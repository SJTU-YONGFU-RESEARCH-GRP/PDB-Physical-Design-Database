module ahb_lite_master (hbusreq,
    hclk,
    hgrant,
    hready,
    hreset,
    hwrite,
    start_trans,
    trans_done,
    trans_write,
    haddr,
    hburst,
    hrdata,
    hresp,
    hsize,
    htrans,
    hwdata,
    read_data,
    trans_addr,
    trans_burst,
    trans_resp,
    trans_size,
    write_data);
 output hbusreq;
 input hclk;
 input hgrant;
 input hready;
 input hreset;
 output hwrite;
 input start_trans;
 output trans_done;
 input trans_write;
 output [31:0] haddr;
 output [2:0] hburst;
 input [31:0] hrdata;
 input [1:0] hresp;
 output [2:0] hsize;
 output [1:0] htrans;
 output [31:0] hwdata;
 output [31:0] read_data;
 input [31:0] trans_addr;
 input [2:0] trans_burst;
 output [1:0] trans_resp;
 input [2:0] trans_size;
 input [31:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire \burst_count[0] ;
 wire \burst_count[1] ;
 wire \burst_count[2] ;
 wire \burst_count[3] ;
 wire \burst_count[4] ;
 wire \burst_count[5] ;
 wire \burst_count[6] ;
 wire \burst_count[7] ;
 wire \burst_total[0] ;
 wire \burst_total[2] ;
 wire \burst_total[3] ;
 wire \burst_total[4] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;

 CLKBUF_X2 _0723_ (.A(\burst_total[3] ),
    .Z(_0130_));
 BUF_X1 _0724_ (.A(\burst_total[0] ),
    .Z(_0131_));
 NOR3_X2 _0725_ (.A1(_0130_),
    .A2(\burst_total[2] ),
    .A3(_0131_),
    .ZN(_0681_));
 XNOR2_X1 _0726_ (.A(_0130_),
    .B(_0691_),
    .ZN(_0686_));
 BUF_X2 _0727_ (.A(net146),
    .Z(_0132_));
 CLKBUF_X2 _0728_ (.A(net145),
    .Z(_0133_));
 INV_X1 _0729_ (.A(_0133_),
    .ZN(_0134_));
 NOR2_X1 _0730_ (.A1(_0132_),
    .A2(_0134_),
    .ZN(_0135_));
 NAND2_X1 _0731_ (.A1(_0007_),
    .A2(_0135_),
    .ZN(_0667_));
 INV_X1 _0732_ (.A(_0667_),
    .ZN(_0700_));
 AND3_X1 _0733_ (.A1(_0132_),
    .A2(_0134_),
    .A3(_0007_),
    .ZN(_0703_));
 AND3_X1 _0734_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0007_),
    .ZN(_0706_));
 INV_X1 _0735_ (.A(net147),
    .ZN(_0136_));
 NOR3_X1 _0736_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0136_),
    .ZN(_0709_));
 NOR3_X1 _0737_ (.A1(_0132_),
    .A2(_0134_),
    .A3(_0136_),
    .ZN(_0712_));
 INV_X1 _0738_ (.A(_0132_),
    .ZN(_0137_));
 NOR3_X1 _0739_ (.A1(_0137_),
    .A2(_0133_),
    .A3(_0136_),
    .ZN(_0715_));
 NOR3_X2 _0740_ (.A1(_0137_),
    .A2(_0134_),
    .A3(_0136_),
    .ZN(_0718_));
 BUF_X2 _0741_ (.A(\state[0] ),
    .Z(_0138_));
 BUF_X2 _0742_ (.A(_0138_),
    .Z(_0139_));
 BUF_X2 _0743_ (.A(\state[1] ),
    .Z(_0140_));
 CLKBUF_X3 _0744_ (.A(_0140_),
    .Z(_0141_));
 BUF_X2 _0745_ (.A(\state[2] ),
    .Z(_0142_));
 INV_X1 _0746_ (.A(_0142_),
    .ZN(_0143_));
 NAND3_X1 _0747_ (.A1(_0139_),
    .A2(_0141_),
    .A3(_0143_),
    .ZN(_0144_));
 CLKBUF_X3 _0748_ (.A(_0000_),
    .Z(_0145_));
 INV_X2 _0749_ (.A(_0145_),
    .ZN(_0146_));
 INV_X2 _0750_ (.A(_0140_),
    .ZN(_0147_));
 AOI21_X1 _0751_ (.A(_0145_),
    .B1(_0142_),
    .B2(_0147_),
    .ZN(_0148_));
 OAI221_X1 _0752_ (.A(_0144_),
    .B1(_0146_),
    .B2(_0141_),
    .C1(_0139_),
    .C2(_0148_),
    .ZN(_0149_));
 INV_X1 _0753_ (.A(_0149_),
    .ZN(_0150_));
 NOR3_X1 _0754_ (.A1(_0139_),
    .A2(net35),
    .A3(_0142_),
    .ZN(_0151_));
 INV_X2 _0755_ (.A(_0138_),
    .ZN(_0152_));
 INV_X1 _0756_ (.A(net35),
    .ZN(_0153_));
 NOR2_X1 _0757_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0154_));
 OAI21_X1 _0758_ (.A(_0141_),
    .B1(_0151_),
    .B2(_0154_),
    .ZN(_0155_));
 INV_X1 _0759_ (.A(net2),
    .ZN(_0156_));
 OAI21_X1 _0760_ (.A(_0138_),
    .B1(_0140_),
    .B2(_0156_),
    .ZN(_0157_));
 CLKBUF_X2 _0761_ (.A(start_trans),
    .Z(_0158_));
 AOI21_X1 _0762_ (.A(_0158_),
    .B1(_0143_),
    .B2(_0141_),
    .ZN(_0159_));
 OAI21_X1 _0763_ (.A(_0157_),
    .B1(_0159_),
    .B2(_0139_),
    .ZN(_0160_));
 NAND3_X1 _0764_ (.A1(_0145_),
    .A2(_0155_),
    .A3(_0160_),
    .ZN(_0161_));
 INV_X1 _0765_ (.A(_0682_),
    .ZN(_0162_));
 NAND3_X1 _0766_ (.A1(_0676_),
    .A2(_0679_),
    .A3(_0685_),
    .ZN(_0163_));
 AOI211_X2 _0767_ (.A(_0687_),
    .B(_0693_),
    .C1(_0695_),
    .C2(_0694_),
    .ZN(_0164_));
 BUF_X1 _0768_ (.A(\burst_count[0] ),
    .Z(_0165_));
 OAI211_X2 _0769_ (.A(_0696_),
    .B(_0694_),
    .C1(_0131_),
    .C2(_0165_),
    .ZN(_0166_));
 INV_X1 _0770_ (.A(_0687_),
    .ZN(_0167_));
 INV_X1 _0771_ (.A(_0688_),
    .ZN(_0168_));
 AOI221_X2 _0772_ (.A(_0163_),
    .B1(_0164_),
    .B2(_0166_),
    .C1(_0167_),
    .C2(_0168_),
    .ZN(_0169_));
 NOR2_X1 _0773_ (.A1(_0672_),
    .A2(_0675_),
    .ZN(_0170_));
 AOI21_X1 _0774_ (.A(_0678_),
    .B1(_0679_),
    .B2(_0684_),
    .ZN(_0171_));
 INV_X1 _0775_ (.A(_0676_),
    .ZN(_0172_));
 OAI21_X1 _0776_ (.A(_0170_),
    .B1(_0171_),
    .B2(_0172_),
    .ZN(_0173_));
 OAI221_X2 _0777_ (.A(_0162_),
    .B1(_0169_),
    .B2(_0173_),
    .C1(_0672_),
    .C2(_0673_),
    .ZN(_0174_));
 NAND3_X1 _0778_ (.A1(_0138_),
    .A2(_0140_),
    .A3(net35),
    .ZN(_0175_));
 OR2_X1 _0779_ (.A1(_0146_),
    .A2(_0175_),
    .ZN(_0176_));
 NOR2_X2 _0780_ (.A1(_0174_),
    .A2(_0176_),
    .ZN(_0177_));
 INV_X1 _0781_ (.A(_0177_),
    .ZN(_0178_));
 AOI21_X1 _0782_ (.A(_0150_),
    .B1(_0161_),
    .B2(_0178_),
    .ZN(_0552_));
 NOR3_X1 _0783_ (.A1(_0139_),
    .A2(_0141_),
    .A3(_0142_),
    .ZN(_0179_));
 NOR3_X1 _0784_ (.A1(_0147_),
    .A2(net35),
    .A3(_0142_),
    .ZN(_0180_));
 OAI21_X1 _0785_ (.A(_0145_),
    .B1(_0157_),
    .B2(_0180_),
    .ZN(_0181_));
 AOI21_X1 _0786_ (.A(_0181_),
    .B1(_0142_),
    .B2(_0158_),
    .ZN(_0182_));
 INV_X1 _0787_ (.A(_0182_),
    .ZN(_0183_));
 AOI221_X1 _0788_ (.A(_0179_),
    .B1(_0183_),
    .B2(_0141_),
    .C1(_0139_),
    .C2(_0181_),
    .ZN(_0553_));
 NOR2_X1 _0789_ (.A1(_0139_),
    .A2(_0158_),
    .ZN(_0184_));
 NAND3_X1 _0790_ (.A1(_0139_),
    .A2(_0145_),
    .A3(_0156_),
    .ZN(_0185_));
 OAI21_X1 _0791_ (.A(_0185_),
    .B1(_0158_),
    .B2(_0145_),
    .ZN(_0186_));
 AOI21_X1 _0792_ (.A(_0184_),
    .B1(_0186_),
    .B2(_0147_),
    .ZN(_0187_));
 MUX2_X1 _0793_ (.A(_0175_),
    .B(_0187_),
    .S(_0142_),
    .Z(_0188_));
 NOR2_X1 _0794_ (.A1(_0146_),
    .A2(_0188_),
    .ZN(_0554_));
 INV_X1 _0795_ (.A(_0698_),
    .ZN(_0668_));
 INV_X1 _0796_ (.A(_0130_),
    .ZN(_0189_));
 INV_X1 _0797_ (.A(\burst_total[4] ),
    .ZN(_0190_));
 NAND3_X1 _0798_ (.A1(_0189_),
    .A2(_0190_),
    .A3(_0691_),
    .ZN(_0671_));
 NOR2_X1 _0799_ (.A1(_0130_),
    .A2(\burst_total[2] ),
    .ZN(_0191_));
 NAND2_X1 _0800_ (.A1(_0131_),
    .A2(_0190_),
    .ZN(_0192_));
 NAND3_X1 _0801_ (.A1(_0680_),
    .A2(_0191_),
    .A3(_0192_),
    .ZN(_0674_));
 NAND2_X1 _0802_ (.A1(_0190_),
    .A2(_0681_),
    .ZN(_0677_));
 NOR3_X2 _0803_ (.A1(_0132_),
    .A2(_0133_),
    .A3(net147),
    .ZN(_0697_));
 NAND3_X4 _0804_ (.A1(_0152_),
    .A2(_0140_),
    .A3(_0145_),
    .ZN(_0193_));
 NOR2_X2 _0805_ (.A1(_0153_),
    .A2(_0193_),
    .ZN(_0194_));
 NAND2_X2 _0806_ (.A1(_0174_),
    .A2(_0194_),
    .ZN(_0195_));
 BUF_X2 _0807_ (.A(_0195_),
    .Z(_0196_));
 NOR2_X2 _0808_ (.A1(_0141_),
    .A2(_0146_),
    .ZN(_0197_));
 NAND3_X2 _0809_ (.A1(_0152_),
    .A2(_0158_),
    .A3(_0197_),
    .ZN(_0198_));
 CLKBUF_X3 _0810_ (.A(_0198_),
    .Z(_0199_));
 NAND3_X1 _0811_ (.A1(_0165_),
    .A2(_0196_),
    .A3(_0199_),
    .ZN(_0200_));
 OAI21_X1 _0812_ (.A(_0200_),
    .B1(_0196_),
    .B2(_0165_),
    .ZN(_0009_));
 NAND3_X1 _0813_ (.A1(\burst_count[1] ),
    .A2(_0196_),
    .A3(_0199_),
    .ZN(_0201_));
 INV_X1 _0814_ (.A(_0722_),
    .ZN(_0202_));
 OAI21_X1 _0815_ (.A(_0201_),
    .B1(_0196_),
    .B2(_0202_),
    .ZN(_0010_));
 BUF_X4 _0816_ (.A(_0193_),
    .Z(_0203_));
 XOR2_X1 _0817_ (.A(_0721_),
    .B(_0005_),
    .Z(_0204_));
 NOR2_X1 _0818_ (.A1(_0203_),
    .A2(_0204_),
    .ZN(_0205_));
 AND2_X1 _0819_ (.A1(_0195_),
    .A2(_0198_),
    .ZN(_0206_));
 MUX2_X1 _0820_ (.A(_0205_),
    .B(\burst_count[2] ),
    .S(_0206_),
    .Z(_0011_));
 INV_X1 _0821_ (.A(\burst_count[3] ),
    .ZN(_0207_));
 NAND3_X1 _0822_ (.A1(_0165_),
    .A2(\burst_count[2] ),
    .A3(\burst_count[1] ),
    .ZN(_0208_));
 NOR3_X4 _0823_ (.A1(_0138_),
    .A2(_0147_),
    .A3(_0146_),
    .ZN(_0209_));
 CLKBUF_X3 _0824_ (.A(_0209_),
    .Z(_0210_));
 AOI22_X1 _0825_ (.A1(_0195_),
    .A2(_0198_),
    .B1(_0208_),
    .B2(_0210_),
    .ZN(_0211_));
 OR3_X1 _0826_ (.A1(\burst_count[3] ),
    .A2(_0203_),
    .A3(_0208_),
    .ZN(_0212_));
 OAI22_X1 _0827_ (.A1(_0207_),
    .A2(_0211_),
    .B1(_0212_),
    .B2(_0206_),
    .ZN(_0012_));
 NAND3_X1 _0828_ (.A1(\burst_count[4] ),
    .A2(_0196_),
    .A3(_0199_),
    .ZN(_0213_));
 NAND3_X1 _0829_ (.A1(_0721_),
    .A2(\burst_count[2] ),
    .A3(\burst_count[3] ),
    .ZN(_0214_));
 XNOR2_X1 _0830_ (.A(_0004_),
    .B(_0214_),
    .ZN(_0215_));
 OAI21_X1 _0831_ (.A(_0213_),
    .B1(_0215_),
    .B2(_0196_),
    .ZN(_0013_));
 NAND3_X1 _0832_ (.A1(\burst_count[5] ),
    .A2(_0196_),
    .A3(_0199_),
    .ZN(_0216_));
 INV_X1 _0833_ (.A(\burst_count[4] ),
    .ZN(_0217_));
 NOR3_X1 _0834_ (.A1(_0207_),
    .A2(_0217_),
    .A3(_0208_),
    .ZN(_0218_));
 XOR2_X1 _0835_ (.A(_0003_),
    .B(_0218_),
    .Z(_0219_));
 OAI21_X1 _0836_ (.A(_0216_),
    .B1(_0219_),
    .B2(_0196_),
    .ZN(_0014_));
 NAND3_X1 _0837_ (.A1(\burst_count[6] ),
    .A2(_0195_),
    .A3(_0199_),
    .ZN(_0220_));
 INV_X1 _0838_ (.A(\burst_count[5] ),
    .ZN(_0221_));
 NOR3_X1 _0839_ (.A1(_0217_),
    .A2(_0221_),
    .A3(_0214_),
    .ZN(_0222_));
 XOR2_X1 _0840_ (.A(_0002_),
    .B(_0222_),
    .Z(_0223_));
 OAI21_X1 _0841_ (.A(_0220_),
    .B1(_0223_),
    .B2(_0196_),
    .ZN(_0015_));
 NAND3_X1 _0842_ (.A1(\burst_count[7] ),
    .A2(_0195_),
    .A3(_0199_),
    .ZN(_0224_));
 NAND3_X1 _0843_ (.A1(\burst_count[5] ),
    .A2(\burst_count[6] ),
    .A3(_0218_),
    .ZN(_0225_));
 XNOR2_X1 _0844_ (.A(_0001_),
    .B(_0225_),
    .ZN(_0226_));
 OAI21_X1 _0845_ (.A(_0224_),
    .B1(_0226_),
    .B2(_0196_),
    .ZN(_0016_));
 BUF_X1 _0846_ (.A(trans_burst[1]),
    .Z(_0227_));
 NOR3_X1 _0847_ (.A1(net72),
    .A2(net71),
    .A3(_0227_),
    .ZN(_0228_));
 MUX2_X1 _0848_ (.A(_0228_),
    .B(_0131_),
    .S(_0198_),
    .Z(_0017_));
 NAND2_X1 _0849_ (.A1(\burst_total[2] ),
    .A2(_0199_),
    .ZN(_0229_));
 INV_X1 _0850_ (.A(net72),
    .ZN(_0230_));
 OAI21_X1 _0851_ (.A(_0230_),
    .B1(net71),
    .B2(_0227_),
    .ZN(_0231_));
 OAI21_X1 _0852_ (.A(_0229_),
    .B1(_0231_),
    .B2(_0199_),
    .ZN(_0018_));
 NOR2_X1 _0853_ (.A1(_0230_),
    .A2(_0227_),
    .ZN(_0232_));
 MUX2_X1 _0854_ (.A(_0232_),
    .B(_0130_),
    .S(_0198_),
    .Z(_0019_));
 NAND2_X1 _0855_ (.A1(\burst_total[4] ),
    .A2(_0199_),
    .ZN(_0233_));
 NAND2_X1 _0856_ (.A1(net72),
    .A2(_0227_),
    .ZN(_0234_));
 OAI21_X1 _0857_ (.A(_0233_),
    .B1(_0234_),
    .B2(_0199_),
    .ZN(_0020_));
 BUF_X2 _0858_ (.A(net141),
    .Z(_0235_));
 NOR3_X1 _0859_ (.A1(_0152_),
    .A2(_0140_),
    .A3(_0146_),
    .ZN(_0236_));
 AND2_X1 _0860_ (.A1(net2),
    .A2(_0236_),
    .ZN(_0237_));
 CLKBUF_X3 _0861_ (.A(_0237_),
    .Z(_0238_));
 MUX2_X1 _0862_ (.A(_0235_),
    .B(net71),
    .S(_0238_),
    .Z(_0021_));
 BUF_X2 _0863_ (.A(net142),
    .Z(_0239_));
 MUX2_X1 _0864_ (.A(_0239_),
    .B(_0227_),
    .S(_0238_),
    .Z(_0022_));
 BUF_X2 _0865_ (.A(net143),
    .Z(_0240_));
 MUX2_X1 _0866_ (.A(_0240_),
    .B(net72),
    .S(_0238_),
    .Z(_0023_));
 NOR2_X1 _0867_ (.A1(net144),
    .A2(_0197_),
    .ZN(_0241_));
 NOR2_X1 _0868_ (.A1(_0239_),
    .A2(_0235_),
    .ZN(_0242_));
 NAND2_X1 _0869_ (.A1(_0006_),
    .A2(_0242_),
    .ZN(_0243_));
 NAND2_X1 _0870_ (.A1(_0174_),
    .A2(_0243_),
    .ZN(_0244_));
 AOI221_X1 _0871_ (.A(_0241_),
    .B1(_0244_),
    .B2(_0194_),
    .C1(_0197_),
    .C2(_0184_),
    .ZN(_0024_));
 MUX2_X1 _0872_ (.A(_0133_),
    .B(net73),
    .S(_0238_),
    .Z(_0025_));
 MUX2_X1 _0873_ (.A(_0132_),
    .B(net74),
    .S(_0238_),
    .Z(_0026_));
 MUX2_X1 _0874_ (.A(net147),
    .B(net75),
    .S(_0238_),
    .Z(_0027_));
 NAND4_X1 _0875_ (.A1(_0239_),
    .A2(_0235_),
    .A3(_0240_),
    .A4(_0006_),
    .ZN(_0245_));
 OR3_X1 _0876_ (.A1(_0239_),
    .A2(_0235_),
    .A3(_0240_),
    .ZN(_0246_));
 AND4_X1 _0877_ (.A1(_0174_),
    .A2(_0210_),
    .A3(_0245_),
    .A4(_0246_),
    .ZN(_0247_));
 NOR2_X1 _0878_ (.A1(_0141_),
    .A2(_0156_),
    .ZN(_0248_));
 AOI21_X1 _0879_ (.A(_0139_),
    .B1(_0141_),
    .B2(_0153_),
    .ZN(_0249_));
 OAI21_X1 _0880_ (.A(_0145_),
    .B1(_0248_),
    .B2(_0249_),
    .ZN(_0250_));
 MUX2_X1 _0881_ (.A(_0247_),
    .B(net148),
    .S(_0250_),
    .Z(_0028_));
 OR2_X1 _0882_ (.A1(_0236_),
    .A2(_0247_),
    .ZN(_0251_));
 MUX2_X1 _0883_ (.A(_0251_),
    .B(net149),
    .S(_0250_),
    .Z(_0029_));
 NAND2_X2 _0884_ (.A1(net182),
    .A2(_0194_),
    .ZN(_0252_));
 CLKBUF_X3 _0885_ (.A(_0252_),
    .Z(_0253_));
 MUX2_X1 _0886_ (.A(net77),
    .B(net150),
    .S(_0253_),
    .Z(_0030_));
 MUX2_X1 _0887_ (.A(net78),
    .B(net151),
    .S(_0253_),
    .Z(_0031_));
 MUX2_X1 _0888_ (.A(net79),
    .B(net152),
    .S(_0253_),
    .Z(_0032_));
 MUX2_X1 _0889_ (.A(net80),
    .B(net153),
    .S(_0253_),
    .Z(_0033_));
 MUX2_X1 _0890_ (.A(net81),
    .B(net154),
    .S(_0253_),
    .Z(_0034_));
 MUX2_X1 _0891_ (.A(net82),
    .B(net155),
    .S(_0253_),
    .Z(_0035_));
 MUX2_X1 _0892_ (.A(net83),
    .B(net156),
    .S(_0253_),
    .Z(_0036_));
 MUX2_X1 _0893_ (.A(net84),
    .B(net157),
    .S(_0253_),
    .Z(_0037_));
 MUX2_X1 _0894_ (.A(net85),
    .B(net158),
    .S(_0253_),
    .Z(_0038_));
 MUX2_X1 _0895_ (.A(net86),
    .B(net159),
    .S(_0253_),
    .Z(_0039_));
 CLKBUF_X3 _0896_ (.A(_0252_),
    .Z(_0254_));
 MUX2_X1 _0897_ (.A(net87),
    .B(net160),
    .S(_0254_),
    .Z(_0040_));
 MUX2_X1 _0898_ (.A(net88),
    .B(net161),
    .S(_0254_),
    .Z(_0041_));
 MUX2_X1 _0899_ (.A(net89),
    .B(net162),
    .S(_0254_),
    .Z(_0042_));
 MUX2_X1 _0900_ (.A(net90),
    .B(net163),
    .S(_0254_),
    .Z(_0043_));
 MUX2_X1 _0901_ (.A(net91),
    .B(net164),
    .S(_0254_),
    .Z(_0044_));
 MUX2_X1 _0902_ (.A(net92),
    .B(net165),
    .S(_0254_),
    .Z(_0045_));
 MUX2_X1 _0903_ (.A(net93),
    .B(net166),
    .S(_0254_),
    .Z(_0046_));
 MUX2_X1 _0904_ (.A(net94),
    .B(net167),
    .S(_0254_),
    .Z(_0047_));
 MUX2_X1 _0905_ (.A(net95),
    .B(net168),
    .S(_0254_),
    .Z(_0048_));
 MUX2_X1 _0906_ (.A(net96),
    .B(net169),
    .S(_0254_),
    .Z(_0049_));
 CLKBUF_X3 _0907_ (.A(_0252_),
    .Z(_0255_));
 MUX2_X1 _0908_ (.A(net97),
    .B(net170),
    .S(_0255_),
    .Z(_0050_));
 MUX2_X1 _0909_ (.A(net98),
    .B(net171),
    .S(_0255_),
    .Z(_0051_));
 MUX2_X1 _0910_ (.A(net99),
    .B(net172),
    .S(_0255_),
    .Z(_0052_));
 MUX2_X1 _0911_ (.A(net100),
    .B(net173),
    .S(_0255_),
    .Z(_0053_));
 MUX2_X1 _0912_ (.A(net101),
    .B(net174),
    .S(_0255_),
    .Z(_0054_));
 MUX2_X1 _0913_ (.A(net102),
    .B(net175),
    .S(_0255_),
    .Z(_0055_));
 MUX2_X1 _0914_ (.A(net103),
    .B(net176),
    .S(_0255_),
    .Z(_0056_));
 MUX2_X1 _0915_ (.A(net104),
    .B(net177),
    .S(_0255_),
    .Z(_0057_));
 MUX2_X1 _0916_ (.A(net105),
    .B(net178),
    .S(_0255_),
    .Z(_0058_));
 MUX2_X1 _0917_ (.A(net106),
    .B(net179),
    .S(_0255_),
    .Z(_0059_));
 MUX2_X1 _0918_ (.A(net107),
    .B(net180),
    .S(_0252_),
    .Z(_0060_));
 MUX2_X1 _0919_ (.A(net108),
    .B(net181),
    .S(_0252_),
    .Z(_0061_));
 MUX2_X1 _0920_ (.A(net182),
    .B(net76),
    .S(_0238_),
    .Z(_0062_));
 NAND2_X1 _0921_ (.A1(_0240_),
    .A2(_0006_),
    .ZN(_0256_));
 OAI21_X1 _0922_ (.A(_0246_),
    .B1(_0256_),
    .B2(_0242_),
    .ZN(_0257_));
 NOR3_X2 _0923_ (.A1(_0153_),
    .A2(_0193_),
    .A3(_0257_),
    .ZN(_0258_));
 AOI21_X4 _0924_ (.A(_0238_),
    .B1(_0258_),
    .B2(_0174_),
    .ZN(_0259_));
 CLKBUF_X3 _0925_ (.A(_0259_),
    .Z(_0260_));
 NAND2_X1 _0926_ (.A1(net109),
    .A2(_0260_),
    .ZN(_0261_));
 AND3_X1 _0927_ (.A1(_0239_),
    .A2(_0240_),
    .A3(_0006_),
    .ZN(_0262_));
 NOR2_X2 _0928_ (.A1(_0239_),
    .A2(_0240_),
    .ZN(_0263_));
 OR3_X1 _0929_ (.A1(_0235_),
    .A2(_0262_),
    .A3(_0263_),
    .ZN(_0264_));
 BUF_X8 _0930_ (.A(_0264_),
    .Z(_0265_));
 AND3_X1 _0931_ (.A1(_0699_),
    .A2(_0210_),
    .A3(_0265_),
    .ZN(_0266_));
 BUF_X4 _0932_ (.A(_0203_),
    .Z(_0267_));
 AOI21_X1 _0933_ (.A(_0266_),
    .B1(_0267_),
    .B2(net39),
    .ZN(_0268_));
 BUF_X4 _0934_ (.A(_0259_),
    .Z(_0269_));
 BUF_X4 _0935_ (.A(_0269_),
    .Z(_0270_));
 OAI21_X1 _0936_ (.A(_0261_),
    .B1(_0268_),
    .B2(_0270_),
    .ZN(_0063_));
 BUF_X4 _0937_ (.A(_0259_),
    .Z(_0271_));
 BUF_X4 _0938_ (.A(_0271_),
    .Z(_0272_));
 CLKBUF_X2 _0939_ (.A(net110),
    .Z(_0273_));
 NOR2_X1 _0940_ (.A1(_0716_),
    .A2(_0719_),
    .ZN(_0274_));
 AOI21_X1 _0941_ (.A(_0713_),
    .B1(_0710_),
    .B2(_0714_),
    .ZN(_0275_));
 NAND2_X1 _0942_ (.A1(_0274_),
    .A2(_0275_),
    .ZN(_0276_));
 BUF_X1 _0943_ (.A(_0704_),
    .Z(_0277_));
 BUF_X1 _0944_ (.A(_0707_),
    .Z(_0278_));
 NOR2_X1 _0945_ (.A1(_0277_),
    .A2(_0278_),
    .ZN(_0279_));
 BUF_X1 _0946_ (.A(_0705_),
    .Z(_0280_));
 INV_X1 _0947_ (.A(_0280_),
    .ZN(_0281_));
 BUF_X1 _0948_ (.A(_0669_),
    .Z(_0282_));
 OAI21_X2 _0949_ (.A(_0279_),
    .B1(_0281_),
    .B2(_0282_),
    .ZN(_0283_));
 BUF_X1 _0950_ (.A(_0711_),
    .Z(_0284_));
 AND2_X1 _0951_ (.A1(_0284_),
    .A2(_0714_),
    .ZN(_0285_));
 CLKBUF_X2 _0952_ (.A(_0708_),
    .Z(_0286_));
 OR2_X1 _0953_ (.A1(_0286_),
    .A2(_0278_),
    .ZN(_0287_));
 AND2_X1 _0954_ (.A1(_0285_),
    .A2(_0287_),
    .ZN(_0288_));
 AOI21_X4 _0955_ (.A(_0276_),
    .B1(_0283_),
    .B2(_0288_),
    .ZN(_0289_));
 BUF_X2 _0956_ (.A(net140),
    .Z(_0290_));
 CLKBUF_X2 _0957_ (.A(net139),
    .Z(_0291_));
 INV_X1 _0958_ (.A(_0719_),
    .ZN(_0292_));
 BUF_X1 _0959_ (.A(_0717_),
    .Z(_0293_));
 OAI21_X1 _0960_ (.A(_0720_),
    .B1(_0716_),
    .B2(_0293_),
    .ZN(_0294_));
 NAND2_X2 _0961_ (.A1(_0292_),
    .A2(_0294_),
    .ZN(_0295_));
 NAND3_X1 _0962_ (.A1(_0290_),
    .A2(_0291_),
    .A3(_0295_),
    .ZN(_0296_));
 NAND2_X4 _0963_ (.A1(_0209_),
    .A2(_0265_),
    .ZN(_0297_));
 NOR4_X1 _0964_ (.A1(_0273_),
    .A2(_0289_),
    .A3(_0296_),
    .A4(_0297_),
    .ZN(_0298_));
 AOI21_X1 _0965_ (.A(_0298_),
    .B1(_0267_),
    .B2(net40),
    .ZN(_0299_));
 OR2_X1 _0966_ (.A1(_0289_),
    .A2(_0296_),
    .ZN(_0300_));
 NOR3_X4 _0967_ (.A1(_0235_),
    .A2(_0262_),
    .A3(_0263_),
    .ZN(_0301_));
 NOR2_X4 _0968_ (.A1(_0193_),
    .A2(_0301_),
    .ZN(_0302_));
 BUF_X4 _0969_ (.A(_0302_),
    .Z(_0303_));
 AOI21_X1 _0970_ (.A(_0271_),
    .B1(_0300_),
    .B2(_0303_),
    .ZN(_0304_));
 INV_X1 _0971_ (.A(_0273_),
    .ZN(_0305_));
 OAI22_X1 _0972_ (.A1(_0272_),
    .A2(_0299_),
    .B1(_0304_),
    .B2(_0305_),
    .ZN(_0064_));
 NAND2_X1 _0973_ (.A1(_0290_),
    .A2(_0273_),
    .ZN(_0306_));
 INV_X1 _0974_ (.A(_0008_),
    .ZN(_0307_));
 AOI21_X2 _0975_ (.A(_0701_),
    .B1(_0702_),
    .B2(_0698_),
    .ZN(_0308_));
 NAND3_X1 _0976_ (.A1(_0280_),
    .A2(_0286_),
    .A3(_0284_),
    .ZN(_0309_));
 AOI21_X1 _0977_ (.A(_0278_),
    .B1(_0277_),
    .B2(_0286_),
    .ZN(_0310_));
 INV_X1 _0978_ (.A(_0284_),
    .ZN(_0311_));
 OAI22_X2 _0979_ (.A1(_0308_),
    .A2(_0309_),
    .B1(_0310_),
    .B2(_0311_),
    .ZN(_0312_));
 AOI21_X1 _0980_ (.A(_0710_),
    .B1(_0713_),
    .B2(_0293_),
    .ZN(_0313_));
 NAND2_X1 _0981_ (.A1(_0274_),
    .A2(_0313_),
    .ZN(_0314_));
 INV_X1 _0982_ (.A(_0720_),
    .ZN(_0315_));
 INV_X1 _0983_ (.A(_0716_),
    .ZN(_0316_));
 OAI21_X1 _0984_ (.A(_0293_),
    .B1(_0713_),
    .B2(_0714_),
    .ZN(_0317_));
 AOI21_X1 _0985_ (.A(_0315_),
    .B1(_0316_),
    .B2(_0317_),
    .ZN(_0318_));
 OAI221_X1 _0986_ (.A(_0307_),
    .B1(_0312_),
    .B2(_0314_),
    .C1(_0318_),
    .C2(_0719_),
    .ZN(_0319_));
 BUF_X2 _0987_ (.A(_0319_),
    .Z(_0320_));
 NOR4_X1 _0988_ (.A1(net111),
    .A2(_0297_),
    .A3(_0306_),
    .A4(_0320_),
    .ZN(_0321_));
 AOI21_X1 _0989_ (.A(_0321_),
    .B1(_0267_),
    .B2(net41),
    .ZN(_0322_));
 CLKBUF_X3 _0990_ (.A(_0302_),
    .Z(_0323_));
 BUF_X4 _0991_ (.A(_0320_),
    .Z(_0324_));
 OR2_X1 _0992_ (.A1(_0306_),
    .A2(_0324_),
    .ZN(_0325_));
 AOI21_X1 _0993_ (.A(_0271_),
    .B1(_0323_),
    .B2(_0325_),
    .ZN(_0326_));
 INV_X1 _0994_ (.A(net111),
    .ZN(_0327_));
 OAI22_X1 _0995_ (.A1(_0272_),
    .A2(_0322_),
    .B1(_0326_),
    .B2(_0327_),
    .ZN(_0065_));
 BUF_X2 _0996_ (.A(net112),
    .Z(_0328_));
 CLKBUF_X3 _0997_ (.A(_0297_),
    .Z(_0329_));
 AND3_X2 _0998_ (.A1(_0290_),
    .A2(_0273_),
    .A3(net111),
    .ZN(_0330_));
 AND3_X1 _0999_ (.A1(_0291_),
    .A2(_0295_),
    .A3(_0330_),
    .ZN(_0331_));
 AND2_X1 _1000_ (.A1(_0274_),
    .A2(_0275_),
    .ZN(_0332_));
 OR2_X1 _1001_ (.A1(_0277_),
    .A2(_0278_),
    .ZN(_0333_));
 INV_X1 _1002_ (.A(_0282_),
    .ZN(_0334_));
 AOI21_X1 _1003_ (.A(_0333_),
    .B1(_0280_),
    .B2(_0334_),
    .ZN(_0335_));
 NAND2_X1 _1004_ (.A1(_0285_),
    .A2(_0287_),
    .ZN(_0336_));
 OAI21_X1 _1005_ (.A(_0332_),
    .B1(_0335_),
    .B2(_0336_),
    .ZN(_0337_));
 BUF_X2 _1006_ (.A(_0337_),
    .Z(_0338_));
 AOI21_X1 _1007_ (.A(_0329_),
    .B1(_0331_),
    .B2(_0338_),
    .ZN(_0339_));
 OAI21_X1 _1008_ (.A(_0328_),
    .B1(_0260_),
    .B2(_0339_),
    .ZN(_0340_));
 NAND3_X1 _1009_ (.A1(_0291_),
    .A2(_0295_),
    .A3(_0330_),
    .ZN(_0341_));
 NOR2_X1 _1010_ (.A1(_0289_),
    .A2(_0341_),
    .ZN(_0342_));
 NOR2_X1 _1011_ (.A1(_0328_),
    .A2(_0329_),
    .ZN(_0343_));
 AOI22_X1 _1012_ (.A1(net42),
    .A2(_0267_),
    .B1(_0342_),
    .B2(_0343_),
    .ZN(_0344_));
 OAI21_X1 _1013_ (.A(_0340_),
    .B1(_0344_),
    .B2(_0270_),
    .ZN(_0066_));
 BUF_X2 _1014_ (.A(net113),
    .Z(_0345_));
 CLKBUF_X3 _1015_ (.A(_0259_),
    .Z(_0346_));
 NAND2_X1 _1016_ (.A1(_0345_),
    .A2(_0346_),
    .ZN(_0347_));
 NAND3_X2 _1017_ (.A1(_0290_),
    .A2(_0273_),
    .A3(net111),
    .ZN(_0348_));
 NOR2_X2 _1018_ (.A1(_0320_),
    .A2(_0348_),
    .ZN(_0349_));
 INV_X1 _1019_ (.A(_0328_),
    .ZN(_0350_));
 NOR3_X1 _1020_ (.A1(_0350_),
    .A2(_0345_),
    .A3(_0297_),
    .ZN(_0351_));
 AOI22_X1 _1021_ (.A1(net43),
    .A2(_0203_),
    .B1(_0349_),
    .B2(_0351_),
    .ZN(_0352_));
 NOR3_X1 _1022_ (.A1(_0350_),
    .A2(_0324_),
    .A3(_0348_),
    .ZN(_0353_));
 NAND2_X1 _1023_ (.A1(_0345_),
    .A2(_0323_),
    .ZN(_0354_));
 OAI221_X1 _1024_ (.A(_0347_),
    .B1(_0352_),
    .B2(_0260_),
    .C1(_0353_),
    .C2(_0354_),
    .ZN(_0067_));
 BUF_X4 _1025_ (.A(net114),
    .Z(_0355_));
 AND2_X2 _1026_ (.A1(_0328_),
    .A2(_0345_),
    .ZN(_0356_));
 AND4_X2 _1027_ (.A1(_0291_),
    .A2(_0295_),
    .A3(_0330_),
    .A4(_0356_),
    .ZN(_0357_));
 AOI21_X1 _1028_ (.A(_0329_),
    .B1(_0357_),
    .B2(_0338_),
    .ZN(_0358_));
 OAI21_X1 _1029_ (.A(_0355_),
    .B1(_0260_),
    .B2(_0358_),
    .ZN(_0359_));
 NAND4_X2 _1030_ (.A1(_0291_),
    .A2(_0295_),
    .A3(_0330_),
    .A4(_0356_),
    .ZN(_0360_));
 NOR2_X1 _1031_ (.A1(_0289_),
    .A2(_0360_),
    .ZN(_0361_));
 NOR2_X1 _1032_ (.A1(_0355_),
    .A2(_0329_),
    .ZN(_0362_));
 AOI22_X1 _1033_ (.A1(net44),
    .A2(_0267_),
    .B1(_0361_),
    .B2(_0362_),
    .ZN(_0363_));
 OAI21_X1 _1034_ (.A(_0359_),
    .B1(_0363_),
    .B2(_0270_),
    .ZN(_0068_));
 BUF_X4 _1035_ (.A(net115),
    .Z(_0364_));
 NAND2_X1 _1036_ (.A1(_0364_),
    .A2(_0346_),
    .ZN(_0365_));
 NAND2_X1 _1037_ (.A1(_0355_),
    .A2(_0356_),
    .ZN(_0366_));
 NOR3_X1 _1038_ (.A1(_0364_),
    .A2(_0297_),
    .A3(_0366_),
    .ZN(_0367_));
 AOI22_X1 _1039_ (.A1(net45),
    .A2(_0203_),
    .B1(_0349_),
    .B2(_0367_),
    .ZN(_0368_));
 NOR3_X1 _1040_ (.A1(_0324_),
    .A2(_0348_),
    .A3(_0366_),
    .ZN(_0369_));
 NAND2_X1 _1041_ (.A1(_0364_),
    .A2(_0323_),
    .ZN(_0370_));
 OAI221_X1 _1042_ (.A(_0365_),
    .B1(_0368_),
    .B2(_0346_),
    .C1(_0369_),
    .C2(_0370_),
    .ZN(_0069_));
 BUF_X4 _1043_ (.A(net116),
    .Z(_0371_));
 INV_X1 _1044_ (.A(_0371_),
    .ZN(_0372_));
 AND3_X1 _1045_ (.A1(_0355_),
    .A2(_0364_),
    .A3(_0356_),
    .ZN(_0373_));
 AND3_X1 _1046_ (.A1(_0372_),
    .A2(_0302_),
    .A3(_0373_),
    .ZN(_0374_));
 AOI22_X1 _1047_ (.A1(net46),
    .A2(_0267_),
    .B1(_0342_),
    .B2(_0374_),
    .ZN(_0375_));
 NAND3_X1 _1048_ (.A1(_0338_),
    .A2(_0331_),
    .A3(_0373_),
    .ZN(_0376_));
 AOI21_X1 _1049_ (.A(_0271_),
    .B1(_0323_),
    .B2(_0376_),
    .ZN(_0377_));
 OAI22_X1 _1050_ (.A1(_0272_),
    .A2(_0375_),
    .B1(_0377_),
    .B2(_0372_),
    .ZN(_0070_));
 BUF_X4 _1051_ (.A(net117),
    .Z(_0378_));
 NAND2_X1 _1052_ (.A1(_0378_),
    .A2(_0346_),
    .ZN(_0379_));
 NAND2_X1 _1053_ (.A1(_0378_),
    .A2(_0303_),
    .ZN(_0380_));
 NAND2_X2 _1054_ (.A1(_0330_),
    .A2(_0356_),
    .ZN(_0381_));
 NAND3_X1 _1055_ (.A1(_0355_),
    .A2(_0364_),
    .A3(_0371_),
    .ZN(_0382_));
 NOR3_X1 _1056_ (.A1(_0324_),
    .A2(_0381_),
    .A3(_0382_),
    .ZN(_0383_));
 CLKBUF_X3 _1057_ (.A(_0193_),
    .Z(_0384_));
 NOR2_X1 _1058_ (.A1(_0378_),
    .A2(_0382_),
    .ZN(_0385_));
 NOR3_X1 _1059_ (.A1(_0297_),
    .A2(_0320_),
    .A3(_0381_),
    .ZN(_0386_));
 AOI22_X1 _1060_ (.A1(net47),
    .A2(_0384_),
    .B1(_0385_),
    .B2(_0386_),
    .ZN(_0387_));
 OAI221_X1 _1061_ (.A(_0379_),
    .B1(_0380_),
    .B2(_0383_),
    .C1(_0260_),
    .C2(_0387_),
    .ZN(_0071_));
 INV_X1 _1062_ (.A(net118),
    .ZN(_0388_));
 INV_X1 _1063_ (.A(_0378_),
    .ZN(_0389_));
 NOR2_X1 _1064_ (.A1(_0389_),
    .A2(_0382_),
    .ZN(_0390_));
 AND3_X1 _1065_ (.A1(_0388_),
    .A2(_0302_),
    .A3(_0390_),
    .ZN(_0391_));
 AOI22_X1 _1066_ (.A1(net48),
    .A2(_0267_),
    .B1(_0361_),
    .B2(_0391_),
    .ZN(_0392_));
 NAND3_X1 _1067_ (.A1(_0338_),
    .A2(_0357_),
    .A3(_0390_),
    .ZN(_0393_));
 AOI21_X1 _1068_ (.A(_0271_),
    .B1(_0323_),
    .B2(_0393_),
    .ZN(_0394_));
 OAI22_X1 _1069_ (.A1(_0272_),
    .A2(_0392_),
    .B1(_0394_),
    .B2(_0388_),
    .ZN(_0072_));
 BUF_X4 _1070_ (.A(net119),
    .Z(_0395_));
 NAND2_X1 _1071_ (.A1(_0395_),
    .A2(_0346_),
    .ZN(_0396_));
 NAND2_X1 _1072_ (.A1(_0395_),
    .A2(_0303_),
    .ZN(_0397_));
 NAND4_X1 _1073_ (.A1(_0371_),
    .A2(_0378_),
    .A3(net118),
    .A4(_0373_),
    .ZN(_0398_));
 NOR3_X1 _1074_ (.A1(_0320_),
    .A2(_0348_),
    .A3(_0398_),
    .ZN(_0399_));
 NOR2_X1 _1075_ (.A1(_0395_),
    .A2(_0297_),
    .ZN(_0400_));
 AOI22_X1 _1076_ (.A1(net49),
    .A2(_0384_),
    .B1(_0400_),
    .B2(_0399_),
    .ZN(_0401_));
 OAI221_X1 _1077_ (.A(_0396_),
    .B1(_0397_),
    .B2(_0399_),
    .C1(_0260_),
    .C2(_0401_),
    .ZN(_0073_));
 NAND2_X1 _1078_ (.A1(net120),
    .A2(_0260_),
    .ZN(_0402_));
 AND3_X1 _1079_ (.A1(_0670_),
    .A2(_0210_),
    .A3(_0265_),
    .ZN(_0403_));
 AOI21_X1 _1080_ (.A(_0403_),
    .B1(_0267_),
    .B2(net50),
    .ZN(_0404_));
 OAI21_X1 _1081_ (.A(_0402_),
    .B1(_0404_),
    .B2(_0270_),
    .ZN(_0074_));
 NAND4_X4 _1082_ (.A1(_0355_),
    .A2(_0364_),
    .A3(_0371_),
    .A4(_0395_),
    .ZN(_0405_));
 NAND4_X4 _1083_ (.A1(_0328_),
    .A2(_0345_),
    .A3(_0378_),
    .A4(net118),
    .ZN(_0406_));
 NOR2_X1 _1084_ (.A1(_0405_),
    .A2(_0406_),
    .ZN(_0407_));
 AND3_X1 _1085_ (.A1(_0338_),
    .A2(_0331_),
    .A3(_0407_),
    .ZN(_0408_));
 NOR2_X1 _1086_ (.A1(net121),
    .A2(_0329_),
    .ZN(_0409_));
 AOI22_X1 _1087_ (.A1(net51),
    .A2(_0384_),
    .B1(_0408_),
    .B2(_0409_),
    .ZN(_0410_));
 NAND3_X1 _1088_ (.A1(_0338_),
    .A2(_0331_),
    .A3(_0407_),
    .ZN(_0411_));
 AOI21_X1 _1089_ (.A(_0269_),
    .B1(_0323_),
    .B2(_0411_),
    .ZN(_0412_));
 INV_X1 _1090_ (.A(net121),
    .ZN(_0413_));
 OAI22_X1 _1091_ (.A1(_0272_),
    .A2(_0410_),
    .B1(_0412_),
    .B2(_0413_),
    .ZN(_0075_));
 NOR2_X1 _1092_ (.A1(net122),
    .A2(_0329_),
    .ZN(_0414_));
 OR4_X1 _1093_ (.A1(_0389_),
    .A2(_0388_),
    .A3(_0413_),
    .A4(_0405_),
    .ZN(_0415_));
 NOR3_X1 _1094_ (.A1(_0324_),
    .A2(_0381_),
    .A3(_0415_),
    .ZN(_0416_));
 AOI22_X1 _1095_ (.A1(net52),
    .A2(_0384_),
    .B1(_0414_),
    .B2(_0416_),
    .ZN(_0417_));
 OR3_X1 _1096_ (.A1(_0320_),
    .A2(_0381_),
    .A3(_0415_),
    .ZN(_0418_));
 AOI21_X1 _1097_ (.A(_0269_),
    .B1(_0323_),
    .B2(_0418_),
    .ZN(_0419_));
 INV_X1 _1098_ (.A(net122),
    .ZN(_0420_));
 OAI22_X1 _1099_ (.A1(_0272_),
    .A2(_0417_),
    .B1(_0419_),
    .B2(_0420_),
    .ZN(_0076_));
 NAND4_X2 _1100_ (.A1(_0378_),
    .A2(net118),
    .A3(net121),
    .A4(net122),
    .ZN(_0421_));
 NOR2_X1 _1101_ (.A1(_0405_),
    .A2(_0421_),
    .ZN(_0422_));
 AND3_X1 _1102_ (.A1(_0338_),
    .A2(_0357_),
    .A3(_0422_),
    .ZN(_0423_));
 NOR2_X1 _1103_ (.A1(net123),
    .A2(_0329_),
    .ZN(_0424_));
 AOI22_X1 _1104_ (.A1(net53),
    .A2(_0384_),
    .B1(_0423_),
    .B2(_0424_),
    .ZN(_0425_));
 NAND3_X1 _1105_ (.A1(_0338_),
    .A2(_0357_),
    .A3(_0422_),
    .ZN(_0426_));
 AOI21_X1 _1106_ (.A(_0269_),
    .B1(_0323_),
    .B2(_0426_),
    .ZN(_0427_));
 INV_X1 _1107_ (.A(net123),
    .ZN(_0428_));
 OAI22_X1 _1108_ (.A1(_0272_),
    .A2(_0425_),
    .B1(_0427_),
    .B2(_0428_),
    .ZN(_0077_));
 BUF_X2 _1109_ (.A(net124),
    .Z(_0429_));
 NAND2_X1 _1110_ (.A1(_0429_),
    .A2(_0346_),
    .ZN(_0430_));
 INV_X1 _1111_ (.A(_0429_),
    .ZN(_0431_));
 NAND3_X2 _1112_ (.A1(net121),
    .A2(net122),
    .A3(net123),
    .ZN(_0432_));
 NOR3_X1 _1113_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_0432_),
    .ZN(_0433_));
 AND3_X1 _1114_ (.A1(_0431_),
    .A2(_0302_),
    .A3(_0433_),
    .ZN(_0434_));
 AOI22_X1 _1115_ (.A1(net54),
    .A2(_0203_),
    .B1(_0349_),
    .B2(_0434_),
    .ZN(_0435_));
 AND2_X1 _1116_ (.A1(_0349_),
    .A2(_0433_),
    .ZN(_0436_));
 NAND2_X1 _1117_ (.A1(_0429_),
    .A2(_0323_),
    .ZN(_0437_));
 OAI221_X1 _1118_ (.A(_0430_),
    .B1(_0435_),
    .B2(_0346_),
    .C1(_0436_),
    .C2(_0437_),
    .ZN(_0078_));
 BUF_X4 _1119_ (.A(net125),
    .Z(_0438_));
 NAND2_X1 _1120_ (.A1(_0438_),
    .A2(_0346_),
    .ZN(_0439_));
 OR3_X1 _1121_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_0432_),
    .ZN(_0440_));
 NOR4_X1 _1122_ (.A1(_0431_),
    .A2(_0438_),
    .A3(_0297_),
    .A4(_0440_),
    .ZN(_0441_));
 AOI22_X1 _1123_ (.A1(net55),
    .A2(_0203_),
    .B1(_0342_),
    .B2(_0441_),
    .ZN(_0442_));
 NOR3_X1 _1124_ (.A1(_0431_),
    .A2(_0411_),
    .A3(_0432_),
    .ZN(_0443_));
 NAND2_X1 _1125_ (.A1(_0438_),
    .A2(_0323_),
    .ZN(_0444_));
 OAI221_X1 _1126_ (.A(_0439_),
    .B1(_0442_),
    .B2(_0346_),
    .C1(_0443_),
    .C2(_0444_),
    .ZN(_0079_));
 BUF_X4 _1127_ (.A(net126),
    .Z(_0445_));
 NAND2_X1 _1128_ (.A1(_0445_),
    .A2(_0346_),
    .ZN(_0446_));
 NAND2_X1 _1129_ (.A1(_0445_),
    .A2(_0303_),
    .ZN(_0447_));
 NAND3_X1 _1130_ (.A1(net123),
    .A2(_0429_),
    .A3(_0438_),
    .ZN(_0448_));
 NOR3_X2 _1131_ (.A1(_0405_),
    .A2(_0421_),
    .A3(_0448_),
    .ZN(_0449_));
 INV_X1 _1132_ (.A(_0449_),
    .ZN(_0450_));
 NOR3_X1 _1133_ (.A1(_0324_),
    .A2(_0381_),
    .A3(_0450_),
    .ZN(_0451_));
 NOR2_X1 _1134_ (.A1(_0445_),
    .A2(_0450_),
    .ZN(_0452_));
 AOI22_X1 _1135_ (.A1(net56),
    .A2(_0203_),
    .B1(_0386_),
    .B2(_0452_),
    .ZN(_0453_));
 OAI221_X1 _1136_ (.A(_0446_),
    .B1(_0447_),
    .B2(_0451_),
    .C1(_0260_),
    .C2(_0453_),
    .ZN(_0080_));
 AND4_X1 _1137_ (.A1(_0445_),
    .A2(_0337_),
    .A3(_0357_),
    .A4(_0449_),
    .ZN(_0454_));
 NOR2_X1 _1138_ (.A1(net127),
    .A2(_0329_),
    .ZN(_0455_));
 AOI22_X1 _1139_ (.A1(net57),
    .A2(_0384_),
    .B1(_0454_),
    .B2(_0455_),
    .ZN(_0456_));
 NAND4_X1 _1140_ (.A1(_0445_),
    .A2(_0338_),
    .A3(_0357_),
    .A4(_0449_),
    .ZN(_0457_));
 AOI21_X1 _1141_ (.A(_0269_),
    .B1(_0303_),
    .B2(_0457_),
    .ZN(_0458_));
 INV_X1 _1142_ (.A(net127),
    .ZN(_0459_));
 OAI22_X1 _1143_ (.A1(_0272_),
    .A2(_0456_),
    .B1(_0458_),
    .B2(_0459_),
    .ZN(_0081_));
 CLKBUF_X2 _1144_ (.A(net128),
    .Z(_0460_));
 NAND2_X1 _1145_ (.A1(_0460_),
    .A2(_0271_),
    .ZN(_0461_));
 NAND2_X1 _1146_ (.A1(_0460_),
    .A2(_0303_),
    .ZN(_0462_));
 NAND4_X2 _1147_ (.A1(_0429_),
    .A2(_0438_),
    .A3(_0445_),
    .A4(net127),
    .ZN(_0463_));
 NOR4_X4 _1148_ (.A1(_0405_),
    .A2(_0406_),
    .A3(_0432_),
    .A4(_0463_),
    .ZN(_0464_));
 AND2_X1 _1149_ (.A1(_0349_),
    .A2(_0464_),
    .ZN(_0465_));
 NAND3_X1 _1150_ (.A1(_0210_),
    .A2(_0265_),
    .A3(_0464_),
    .ZN(_0466_));
 NOR2_X1 _1151_ (.A1(_0460_),
    .A2(_0466_),
    .ZN(_0467_));
 AOI22_X1 _1152_ (.A1(net58),
    .A2(_0203_),
    .B1(_0349_),
    .B2(_0467_),
    .ZN(_0468_));
 OAI221_X1 _1153_ (.A(_0461_),
    .B1(_0462_),
    .B2(_0465_),
    .C1(_0260_),
    .C2(_0468_),
    .ZN(_0082_));
 NOR2_X1 _1154_ (.A1(net129),
    .A2(_0329_),
    .ZN(_0469_));
 NAND2_X1 _1155_ (.A1(_0460_),
    .A2(_0464_),
    .ZN(_0470_));
 NOR3_X1 _1156_ (.A1(_0289_),
    .A2(_0341_),
    .A3(_0470_),
    .ZN(_0471_));
 AOI22_X1 _1157_ (.A1(net59),
    .A2(_0384_),
    .B1(_0469_),
    .B2(_0471_),
    .ZN(_0472_));
 OR3_X1 _1158_ (.A1(_0289_),
    .A2(_0341_),
    .A3(_0470_),
    .ZN(_0473_));
 AOI21_X1 _1159_ (.A(_0269_),
    .B1(_0303_),
    .B2(_0473_),
    .ZN(_0474_));
 INV_X1 _1160_ (.A(net129),
    .ZN(_0475_));
 OAI22_X1 _1161_ (.A1(_0270_),
    .A2(_0472_),
    .B1(_0474_),
    .B2(_0475_),
    .ZN(_0083_));
 OR4_X1 _1162_ (.A1(_0428_),
    .A2(_0405_),
    .A3(_0421_),
    .A4(_0463_),
    .ZN(_0476_));
 NAND2_X1 _1163_ (.A1(_0460_),
    .A2(net129),
    .ZN(_0477_));
 OR3_X1 _1164_ (.A1(_0381_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0478_));
 NOR4_X1 _1165_ (.A1(net130),
    .A2(_0297_),
    .A3(_0324_),
    .A4(_0478_),
    .ZN(_0479_));
 AOI21_X1 _1166_ (.A(_0479_),
    .B1(_0267_),
    .B2(net60),
    .ZN(_0480_));
 OR2_X1 _1167_ (.A1(_0324_),
    .A2(_0478_),
    .ZN(_0481_));
 AOI21_X1 _1168_ (.A(_0269_),
    .B1(_0303_),
    .B2(_0481_),
    .ZN(_0482_));
 INV_X1 _1169_ (.A(net130),
    .ZN(_0483_));
 OAI22_X1 _1170_ (.A1(_0270_),
    .A2(_0480_),
    .B1(_0482_),
    .B2(_0483_),
    .ZN(_0084_));
 XOR2_X1 _1171_ (.A(_0282_),
    .B(_0280_),
    .Z(_0484_));
 NOR2_X1 _1172_ (.A1(_0193_),
    .A2(_0484_),
    .ZN(_0485_));
 AOI221_X2 _1173_ (.A(_0259_),
    .B1(_0265_),
    .B2(_0485_),
    .C1(_0193_),
    .C2(net61),
    .ZN(_0486_));
 INV_X1 _1174_ (.A(net131),
    .ZN(_0487_));
 AOI21_X1 _1175_ (.A(_0486_),
    .B1(_0272_),
    .B2(_0487_),
    .ZN(_0085_));
 NOR2_X1 _1176_ (.A1(net132),
    .A2(_0329_),
    .ZN(_0488_));
 OR3_X1 _1177_ (.A1(_0483_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0489_));
 NOR3_X1 _1178_ (.A1(_0289_),
    .A2(_0360_),
    .A3(_0489_),
    .ZN(_0490_));
 AOI22_X1 _1179_ (.A1(net62),
    .A2(_0384_),
    .B1(_0488_),
    .B2(_0490_),
    .ZN(_0491_));
 OR3_X1 _1180_ (.A1(_0289_),
    .A2(_0360_),
    .A3(_0489_),
    .ZN(_0492_));
 AOI21_X1 _1181_ (.A(_0269_),
    .B1(_0303_),
    .B2(_0492_),
    .ZN(_0493_));
 INV_X1 _1182_ (.A(net132),
    .ZN(_0494_));
 OAI22_X1 _1183_ (.A1(_0270_),
    .A2(_0491_),
    .B1(_0493_),
    .B2(_0494_),
    .ZN(_0086_));
 NAND2_X1 _1184_ (.A1(net133),
    .A2(_0271_),
    .ZN(_0495_));
 NAND2_X1 _1185_ (.A1(net133),
    .A2(_0302_),
    .ZN(_0496_));
 NOR2_X1 _1186_ (.A1(_0483_),
    .A2(_0477_),
    .ZN(_0497_));
 AND4_X1 _1187_ (.A1(net132),
    .A2(_0349_),
    .A3(_0464_),
    .A4(_0497_),
    .ZN(_0498_));
 INV_X1 _1188_ (.A(net133),
    .ZN(_0499_));
 NAND3_X1 _1189_ (.A1(net132),
    .A2(_0499_),
    .A3(_0497_),
    .ZN(_0500_));
 NOR2_X1 _1190_ (.A1(_0466_),
    .A2(_0500_),
    .ZN(_0501_));
 AOI22_X1 _1191_ (.A1(net63),
    .A2(_0203_),
    .B1(_0349_),
    .B2(_0501_),
    .ZN(_0502_));
 OAI221_X1 _1192_ (.A(_0495_),
    .B1(_0496_),
    .B2(_0498_),
    .C1(_0260_),
    .C2(_0502_),
    .ZN(_0087_));
 INV_X1 _1193_ (.A(_0277_),
    .ZN(_0503_));
 OAI21_X1 _1194_ (.A(_0503_),
    .B1(_0308_),
    .B2(_0281_),
    .ZN(_0504_));
 NOR2_X1 _1195_ (.A1(_0286_),
    .A2(_0504_),
    .ZN(_0505_));
 OAI21_X1 _1196_ (.A(_0286_),
    .B1(_0277_),
    .B2(_0280_),
    .ZN(_0506_));
 NOR2_X1 _1197_ (.A1(_0701_),
    .A2(_0277_),
    .ZN(_0507_));
 NAND2_X1 _1198_ (.A1(_0698_),
    .A2(_0702_),
    .ZN(_0508_));
 AOI21_X1 _1199_ (.A(_0506_),
    .B1(_0507_),
    .B2(_0508_),
    .ZN(_0509_));
 NOR3_X1 _1200_ (.A1(_0301_),
    .A2(_0505_),
    .A3(_0509_),
    .ZN(_0510_));
 MUX2_X1 _1201_ (.A(net64),
    .B(_0510_),
    .S(_0210_),
    .Z(_0511_));
 MUX2_X1 _1202_ (.A(_0511_),
    .B(net134),
    .S(_0271_),
    .Z(_0088_));
 NOR2_X1 _1203_ (.A1(_0284_),
    .A2(_0301_),
    .ZN(_0512_));
 NOR2_X1 _1204_ (.A1(_0311_),
    .A2(_0301_),
    .ZN(_0513_));
 OAI21_X1 _1205_ (.A(_0503_),
    .B1(_0281_),
    .B2(_0282_),
    .ZN(_0514_));
 AOI21_X1 _1206_ (.A(_0278_),
    .B1(_0514_),
    .B2(_0286_),
    .ZN(_0515_));
 MUX2_X1 _1207_ (.A(_0512_),
    .B(_0513_),
    .S(_0515_),
    .Z(_0516_));
 MUX2_X1 _1208_ (.A(net65),
    .B(_0516_),
    .S(_0210_),
    .Z(_0517_));
 MUX2_X1 _1209_ (.A(_0517_),
    .B(net135),
    .S(_0271_),
    .Z(_0089_));
 INV_X1 _1210_ (.A(net136),
    .ZN(_0518_));
 NOR2_X1 _1211_ (.A1(_0710_),
    .A2(_0312_),
    .ZN(_0519_));
 XNOR2_X1 _1212_ (.A(_0714_),
    .B(_0519_),
    .ZN(_0520_));
 NAND3_X1 _1213_ (.A1(_0210_),
    .A2(_0265_),
    .A3(_0520_),
    .ZN(_0521_));
 AOI21_X1 _1214_ (.A(_0269_),
    .B1(_0384_),
    .B2(net66),
    .ZN(_0522_));
 AOI22_X1 _1215_ (.A1(_0518_),
    .A2(_0270_),
    .B1(_0521_),
    .B2(_0522_),
    .ZN(_0090_));
 AND2_X1 _1216_ (.A1(_0293_),
    .A2(_0265_),
    .ZN(_0523_));
 NOR2_X1 _1217_ (.A1(_0293_),
    .A2(_0301_),
    .ZN(_0524_));
 OAI21_X1 _1218_ (.A(_0275_),
    .B1(_0335_),
    .B2(_0336_),
    .ZN(_0525_));
 MUX2_X1 _1219_ (.A(_0523_),
    .B(_0524_),
    .S(_0525_),
    .Z(_0526_));
 MUX2_X1 _1220_ (.A(net67),
    .B(_0526_),
    .S(_0210_),
    .Z(_0527_));
 MUX2_X1 _1221_ (.A(_0527_),
    .B(net137),
    .S(_0271_),
    .Z(_0091_));
 NOR3_X1 _1222_ (.A1(_0284_),
    .A2(_0710_),
    .A3(_0713_),
    .ZN(_0528_));
 OAI21_X1 _1223_ (.A(_0316_),
    .B1(_0317_),
    .B2(_0528_),
    .ZN(_0529_));
 INV_X1 _1224_ (.A(_0278_),
    .ZN(_0530_));
 NAND3_X1 _1225_ (.A1(_0530_),
    .A2(_0316_),
    .A3(_0313_),
    .ZN(_0531_));
 OAI21_X1 _1226_ (.A(_0529_),
    .B1(_0531_),
    .B2(_0509_),
    .ZN(_0532_));
 XNOR2_X1 _1227_ (.A(_0720_),
    .B(_0532_),
    .ZN(_0533_));
 AOI221_X1 _1228_ (.A(_0259_),
    .B1(_0302_),
    .B2(_0533_),
    .C1(_0193_),
    .C2(net68),
    .ZN(_0534_));
 INV_X1 _1229_ (.A(net138),
    .ZN(_0535_));
 AOI21_X1 _1230_ (.A(_0534_),
    .B1(_0272_),
    .B2(_0535_),
    .ZN(_0092_));
 INV_X1 _1231_ (.A(_0291_),
    .ZN(_0536_));
 NAND3_X1 _1232_ (.A1(_0307_),
    .A2(_0338_),
    .A3(_0295_),
    .ZN(_0537_));
 INV_X1 _1233_ (.A(_0295_),
    .ZN(_0538_));
 OAI21_X1 _1234_ (.A(_0008_),
    .B1(_0289_),
    .B2(_0538_),
    .ZN(_0539_));
 NAND4_X1 _1235_ (.A1(_0210_),
    .A2(_0265_),
    .A3(_0537_),
    .A4(_0539_),
    .ZN(_0540_));
 AOI21_X1 _1236_ (.A(_0259_),
    .B1(_0384_),
    .B2(net69),
    .ZN(_0541_));
 AOI22_X1 _1237_ (.A1(_0536_),
    .A2(_0270_),
    .B1(_0540_),
    .B2(_0541_),
    .ZN(_0093_));
 NOR3_X1 _1238_ (.A1(_0290_),
    .A2(_0297_),
    .A3(_0324_),
    .ZN(_0542_));
 AOI21_X1 _1239_ (.A(_0542_),
    .B1(_0267_),
    .B2(net70),
    .ZN(_0543_));
 AOI21_X1 _1240_ (.A(_0269_),
    .B1(_0303_),
    .B2(_0324_),
    .ZN(_0544_));
 INV_X1 _1241_ (.A(_0290_),
    .ZN(_0545_));
 OAI22_X1 _1242_ (.A1(_0270_),
    .A2(_0543_),
    .B1(_0544_),
    .B2(_0545_),
    .ZN(_0094_));
 NOR2_X2 _1243_ (.A1(net182),
    .A2(_0176_),
    .ZN(_0546_));
 CLKBUF_X3 _1244_ (.A(_0546_),
    .Z(_0547_));
 MUX2_X1 _1245_ (.A(net183),
    .B(net3),
    .S(_0547_),
    .Z(_0095_));
 MUX2_X1 _1246_ (.A(net184),
    .B(net4),
    .S(_0547_),
    .Z(_0096_));
 MUX2_X1 _1247_ (.A(net185),
    .B(net5),
    .S(_0547_),
    .Z(_0097_));
 MUX2_X1 _1248_ (.A(net186),
    .B(net6),
    .S(_0547_),
    .Z(_0098_));
 MUX2_X1 _1249_ (.A(net187),
    .B(net7),
    .S(_0547_),
    .Z(_0099_));
 MUX2_X1 _1250_ (.A(net188),
    .B(net8),
    .S(_0547_),
    .Z(_0100_));
 MUX2_X1 _1251_ (.A(net189),
    .B(net9),
    .S(_0547_),
    .Z(_0101_));
 MUX2_X1 _1252_ (.A(net190),
    .B(net10),
    .S(_0547_),
    .Z(_0102_));
 MUX2_X1 _1253_ (.A(net191),
    .B(net11),
    .S(_0547_),
    .Z(_0103_));
 MUX2_X1 _1254_ (.A(net192),
    .B(net12),
    .S(_0547_),
    .Z(_0104_));
 CLKBUF_X3 _1255_ (.A(_0546_),
    .Z(_0548_));
 MUX2_X1 _1256_ (.A(net193),
    .B(net13),
    .S(_0548_),
    .Z(_0105_));
 MUX2_X1 _1257_ (.A(net194),
    .B(net14),
    .S(_0548_),
    .Z(_0106_));
 MUX2_X1 _1258_ (.A(net195),
    .B(net15),
    .S(_0548_),
    .Z(_0107_));
 MUX2_X1 _1259_ (.A(net196),
    .B(net16),
    .S(_0548_),
    .Z(_0108_));
 MUX2_X1 _1260_ (.A(net197),
    .B(net17),
    .S(_0548_),
    .Z(_0109_));
 MUX2_X1 _1261_ (.A(net198),
    .B(net18),
    .S(_0548_),
    .Z(_0110_));
 MUX2_X1 _1262_ (.A(net199),
    .B(net19),
    .S(_0548_),
    .Z(_0111_));
 MUX2_X1 _1263_ (.A(net200),
    .B(net20),
    .S(_0548_),
    .Z(_0112_));
 MUX2_X1 _1264_ (.A(net201),
    .B(net21),
    .S(_0548_),
    .Z(_0113_));
 MUX2_X1 _1265_ (.A(net202),
    .B(net22),
    .S(_0548_),
    .Z(_0114_));
 CLKBUF_X3 _1266_ (.A(_0546_),
    .Z(_0549_));
 MUX2_X1 _1267_ (.A(net203),
    .B(net23),
    .S(_0549_),
    .Z(_0115_));
 MUX2_X1 _1268_ (.A(net204),
    .B(net24),
    .S(_0549_),
    .Z(_0116_));
 MUX2_X1 _1269_ (.A(net205),
    .B(net25),
    .S(_0549_),
    .Z(_0117_));
 MUX2_X1 _1270_ (.A(net206),
    .B(net26),
    .S(_0549_),
    .Z(_0118_));
 MUX2_X1 _1271_ (.A(net207),
    .B(net27),
    .S(_0549_),
    .Z(_0119_));
 MUX2_X1 _1272_ (.A(net208),
    .B(net28),
    .S(_0549_),
    .Z(_0120_));
 MUX2_X1 _1273_ (.A(net209),
    .B(net29),
    .S(_0549_),
    .Z(_0121_));
 MUX2_X1 _1274_ (.A(net210),
    .B(net30),
    .S(_0549_),
    .Z(_0122_));
 MUX2_X1 _1275_ (.A(net211),
    .B(net31),
    .S(_0549_),
    .Z(_0123_));
 MUX2_X1 _1276_ (.A(net212),
    .B(net32),
    .S(_0549_),
    .Z(_0124_));
 MUX2_X1 _1277_ (.A(net213),
    .B(net33),
    .S(_0546_),
    .Z(_0125_));
 MUX2_X1 _1278_ (.A(net214),
    .B(net34),
    .S(_0546_),
    .Z(_0126_));
 XOR2_X1 _1279_ (.A(_0139_),
    .B(_0142_),
    .Z(_0550_));
 OAI22_X1 _1280_ (.A1(net215),
    .A2(_0177_),
    .B1(_0550_),
    .B2(_0141_),
    .ZN(_0551_));
 INV_X1 _1281_ (.A(_0551_),
    .ZN(_0127_));
 MUX2_X1 _1282_ (.A(net216),
    .B(net37),
    .S(_0177_),
    .Z(_0128_));
 MUX2_X1 _1283_ (.A(net217),
    .B(net38),
    .S(_0177_),
    .Z(_0129_));
 FA_X1 _1284_ (.A(_0666_),
    .B(_0667_),
    .CI(_0668_),
    .CO(_0669_),
    .S(_0670_));
 HA_X1 _1285_ (.A(\burst_count[7] ),
    .B(_0671_),
    .CO(_0672_),
    .S(_0673_));
 HA_X1 _1286_ (.A(\burst_count[6] ),
    .B(_0674_),
    .CO(_0675_),
    .S(_0676_));
 HA_X1 _1287_ (.A(\burst_count[5] ),
    .B(_0677_),
    .CO(_0678_),
    .S(_0679_));
 HA_X1 _1288_ (.A(_0680_),
    .B(_0681_),
    .CO(_0682_),
    .S(_0683_));
 HA_X1 _1289_ (.A(\burst_count[4] ),
    .B(_0683_),
    .CO(_0684_),
    .S(_0685_));
 HA_X1 _1290_ (.A(\burst_count[3] ),
    .B(_0686_),
    .CO(_0687_),
    .S(_0688_));
 HA_X1 _1291_ (.A(_0689_),
    .B(_0690_),
    .CO(_0691_),
    .S(_0692_));
 HA_X1 _1292_ (.A(\burst_count[2] ),
    .B(_0692_),
    .CO(_0693_),
    .S(_0694_));
 HA_X1 _1293_ (.A(\burst_count[1] ),
    .B(\burst_total[0] ),
    .CO(_0695_),
    .S(_0696_));
 HA_X1 _1294_ (.A(net109),
    .B(_0697_),
    .CO(_0698_),
    .S(_0699_));
 HA_X1 _1295_ (.A(net120),
    .B(_0700_),
    .CO(_0701_),
    .S(_0702_));
 HA_X1 _1296_ (.A(net131),
    .B(_0703_),
    .CO(_0704_),
    .S(_0705_));
 HA_X1 _1297_ (.A(net134),
    .B(_0706_),
    .CO(_0707_),
    .S(_0708_));
 HA_X1 _1298_ (.A(net135),
    .B(_0709_),
    .CO(_0710_),
    .S(_0711_));
 HA_X1 _1299_ (.A(net136),
    .B(_0712_),
    .CO(_0713_),
    .S(_0714_));
 HA_X1 _1300_ (.A(net137),
    .B(_0715_),
    .CO(_0716_),
    .S(_0717_));
 HA_X1 _1301_ (.A(net138),
    .B(_0718_),
    .CO(_0719_),
    .S(_0720_));
 HA_X1 _1302_ (.A(\burst_count[0] ),
    .B(\burst_count[1] ),
    .CO(_0721_),
    .S(_0722_));
 DFFR_X1 \burst_count[0]$_DFFE_PN0P_  (.D(_0009_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[0] ),
    .QN(_0662_));
 DFFR_X2 \burst_count[1]$_DFFE_PN0P_  (.D(_0010_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[1] ),
    .QN(_0661_));
 DFFR_X1 \burst_count[2]$_DFFE_PN0P_  (.D(_0011_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[2] ),
    .QN(_0005_));
 DFFR_X1 \burst_count[3]$_DFFE_PN0P_  (.D(_0012_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[3] ),
    .QN(_0660_));
 DFFR_X1 \burst_count[4]$_DFFE_PN0P_  (.D(_0013_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[4] ),
    .QN(_0004_));
 DFFR_X2 \burst_count[5]$_DFFE_PN0P_  (.D(_0014_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[5] ),
    .QN(_0003_));
 DFFR_X1 \burst_count[6]$_DFFE_PN0P_  (.D(_0015_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[6] ),
    .QN(_0002_));
 DFFR_X1 \burst_count[7]$_DFFE_PN0P_  (.D(_0016_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_count[7] ),
    .QN(_0001_));
 DFFR_X1 \burst_total[0]$_DFFE_PN0P_  (.D(_0017_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_total[0] ),
    .QN(_0689_));
 DFFR_X1 \burst_total[2]$_DFFE_PN0P_  (.D(_0018_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_total[2] ),
    .QN(_0690_));
 DFFR_X1 \burst_total[3]$_DFFE_PN0P_  (.D(_0019_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_total[3] ),
    .QN(_0659_));
 DFFR_X1 \burst_total[4]$_DFFE_PN0P_  (.D(_0020_),
    .RN(net36),
    .CK(net1),
    .Q(\burst_total[4] ),
    .QN(_0680_));
 DFFR_X1 \hburst[0]$_DFFE_PN0P_  (.D(_0021_),
    .RN(net36),
    .CK(net1),
    .Q(net141),
    .QN(_0658_));
 DFFR_X1 \hburst[1]$_DFFE_PN0P_  (.D(_0022_),
    .RN(net36),
    .CK(net1),
    .Q(net142),
    .QN(_0657_));
 DFFR_X1 \hburst[2]$_DFFE_PN0P_  (.D(_0023_),
    .RN(net36),
    .CK(net1),
    .Q(net143),
    .QN(_0006_));
 DFFR_X1 \hbusreq$_DFFE_PN0P_  (.D(_0024_),
    .RN(net36),
    .CK(net1),
    .Q(net144),
    .QN(_0656_));
 DFFR_X1 \hsize[0]$_DFFE_PN0P_  (.D(_0025_),
    .RN(net36),
    .CK(net1),
    .Q(net145),
    .QN(_0655_));
 DFFR_X1 \hsize[1]$_DFFE_PN0P_  (.D(_0026_),
    .RN(net36),
    .CK(net1),
    .Q(net146),
    .QN(_0654_));
 DFFR_X1 \hsize[2]$_DFFE_PN0P_  (.D(_0027_),
    .RN(net36),
    .CK(net1),
    .Q(net147),
    .QN(_0007_));
 DFFR_X1 \htrans[0]$_DFFE_PN0P_  (.D(_0028_),
    .RN(net36),
    .CK(net1),
    .Q(net148),
    .QN(_0653_));
 DFFR_X1 \htrans[1]$_DFFE_PN0P_  (.D(_0029_),
    .RN(net36),
    .CK(net1),
    .Q(net149),
    .QN(_0652_));
 DFFR_X1 \hwdata[0]$_DFFE_PN0P_  (.D(_0030_),
    .RN(net36),
    .CK(net1),
    .Q(net150),
    .QN(_0651_));
 DFFR_X1 \hwdata[10]$_DFFE_PN0P_  (.D(_0031_),
    .RN(net36),
    .CK(net1),
    .Q(net151),
    .QN(_0650_));
 DFFR_X1 \hwdata[11]$_DFFE_PN0P_  (.D(_0032_),
    .RN(net36),
    .CK(net1),
    .Q(net152),
    .QN(_0649_));
 DFFR_X1 \hwdata[12]$_DFFE_PN0P_  (.D(_0033_),
    .RN(net36),
    .CK(net1),
    .Q(net153),
    .QN(_0648_));
 DFFR_X1 \hwdata[13]$_DFFE_PN0P_  (.D(_0034_),
    .RN(net36),
    .CK(net1),
    .Q(net154),
    .QN(_0647_));
 DFFR_X1 \hwdata[14]$_DFFE_PN0P_  (.D(_0035_),
    .RN(net36),
    .CK(net1),
    .Q(net155),
    .QN(_0646_));
 DFFR_X1 \hwdata[15]$_DFFE_PN0P_  (.D(_0036_),
    .RN(net36),
    .CK(net1),
    .Q(net156),
    .QN(_0645_));
 DFFR_X1 \hwdata[16]$_DFFE_PN0P_  (.D(_0037_),
    .RN(net36),
    .CK(net1),
    .Q(net157),
    .QN(_0644_));
 DFFR_X1 \hwdata[17]$_DFFE_PN0P_  (.D(_0038_),
    .RN(net36),
    .CK(net1),
    .Q(net158),
    .QN(_0643_));
 DFFR_X1 \hwdata[18]$_DFFE_PN0P_  (.D(_0039_),
    .RN(net36),
    .CK(net1),
    .Q(net159),
    .QN(_0642_));
 DFFR_X1 \hwdata[19]$_DFFE_PN0P_  (.D(_0040_),
    .RN(net36),
    .CK(net1),
    .Q(net160),
    .QN(_0641_));
 DFFR_X1 \hwdata[1]$_DFFE_PN0P_  (.D(_0041_),
    .RN(net36),
    .CK(net1),
    .Q(net161),
    .QN(_0640_));
 DFFR_X1 \hwdata[20]$_DFFE_PN0P_  (.D(_0042_),
    .RN(net36),
    .CK(net1),
    .Q(net162),
    .QN(_0639_));
 DFFR_X1 \hwdata[21]$_DFFE_PN0P_  (.D(_0043_),
    .RN(net36),
    .CK(net1),
    .Q(net163),
    .QN(_0638_));
 DFFR_X1 \hwdata[22]$_DFFE_PN0P_  (.D(_0044_),
    .RN(net36),
    .CK(net1),
    .Q(net164),
    .QN(_0637_));
 DFFR_X1 \hwdata[23]$_DFFE_PN0P_  (.D(_0045_),
    .RN(net36),
    .CK(net1),
    .Q(net165),
    .QN(_0636_));
 DFFR_X1 \hwdata[24]$_DFFE_PN0P_  (.D(_0046_),
    .RN(net36),
    .CK(net1),
    .Q(net166),
    .QN(_0635_));
 DFFR_X1 \hwdata[25]$_DFFE_PN0P_  (.D(_0047_),
    .RN(net36),
    .CK(net1),
    .Q(net167),
    .QN(_0634_));
 DFFR_X1 \hwdata[26]$_DFFE_PN0P_  (.D(_0048_),
    .RN(net36),
    .CK(net1),
    .Q(net168),
    .QN(_0633_));
 DFFR_X1 \hwdata[27]$_DFFE_PN0P_  (.D(_0049_),
    .RN(net36),
    .CK(net1),
    .Q(net169),
    .QN(_0632_));
 DFFR_X1 \hwdata[28]$_DFFE_PN0P_  (.D(_0050_),
    .RN(net36),
    .CK(net1),
    .Q(net170),
    .QN(_0631_));
 DFFR_X1 \hwdata[29]$_DFFE_PN0P_  (.D(_0051_),
    .RN(net36),
    .CK(net1),
    .Q(net171),
    .QN(_0630_));
 DFFR_X1 \hwdata[2]$_DFFE_PN0P_  (.D(_0052_),
    .RN(net36),
    .CK(net1),
    .Q(net172),
    .QN(_0629_));
 DFFR_X1 \hwdata[30]$_DFFE_PN0P_  (.D(_0053_),
    .RN(net36),
    .CK(net1),
    .Q(net173),
    .QN(_0628_));
 DFFR_X1 \hwdata[31]$_DFFE_PN0P_  (.D(_0054_),
    .RN(net36),
    .CK(net1),
    .Q(net174),
    .QN(_0627_));
 DFFR_X1 \hwdata[3]$_DFFE_PN0P_  (.D(_0055_),
    .RN(net36),
    .CK(net1),
    .Q(net175),
    .QN(_0626_));
 DFFR_X1 \hwdata[4]$_DFFE_PN0P_  (.D(_0056_),
    .RN(net36),
    .CK(net1),
    .Q(net176),
    .QN(_0625_));
 DFFR_X1 \hwdata[5]$_DFFE_PN0P_  (.D(_0057_),
    .RN(net36),
    .CK(net1),
    .Q(net177),
    .QN(_0624_));
 DFFR_X1 \hwdata[6]$_DFFE_PN0P_  (.D(_0058_),
    .RN(net36),
    .CK(net1),
    .Q(net178),
    .QN(_0623_));
 DFFR_X1 \hwdata[7]$_DFFE_PN0P_  (.D(_0059_),
    .RN(net36),
    .CK(net1),
    .Q(net179),
    .QN(_0622_));
 DFFR_X1 \hwdata[8]$_DFFE_PN0P_  (.D(_0060_),
    .RN(net36),
    .CK(net1),
    .Q(net180),
    .QN(_0621_));
 DFFR_X1 \hwdata[9]$_DFFE_PN0P_  (.D(_0061_),
    .RN(net36),
    .CK(net1),
    .Q(net181),
    .QN(_0620_));
 DFFR_X2 \hwrite$_DFFE_PN0P_  (.D(_0062_),
    .RN(net36),
    .CK(net1),
    .Q(net182),
    .QN(_0619_));
 DFFR_X1 \next_addr[0]$_DFFE_PN0P_  (.D(_0063_),
    .RN(net36),
    .CK(net1),
    .Q(net109),
    .QN(_0618_));
 DFFR_X1 \next_addr[10]$_DFFE_PN0P_  (.D(_0064_),
    .RN(net36),
    .CK(net1),
    .Q(net110),
    .QN(_0617_));
 DFFR_X2 \next_addr[11]$_DFFE_PN0P_  (.D(_0065_),
    .RN(net36),
    .CK(net1),
    .Q(net111),
    .QN(_0616_));
 DFFR_X1 \next_addr[12]$_DFFE_PN0P_  (.D(_0066_),
    .RN(net36),
    .CK(net1),
    .Q(net112),
    .QN(_0615_));
 DFFR_X1 \next_addr[13]$_DFFE_PN0P_  (.D(_0067_),
    .RN(net36),
    .CK(net1),
    .Q(net113),
    .QN(_0614_));
 DFFR_X1 \next_addr[14]$_DFFE_PN0P_  (.D(_0068_),
    .RN(net36),
    .CK(net1),
    .Q(net114),
    .QN(_0613_));
 DFFR_X1 \next_addr[15]$_DFFE_PN0P_  (.D(_0069_),
    .RN(net36),
    .CK(net1),
    .Q(net115),
    .QN(_0612_));
 DFFR_X1 \next_addr[16]$_DFFE_PN0P_  (.D(_0070_),
    .RN(net36),
    .CK(net1),
    .Q(net116),
    .QN(_0611_));
 DFFR_X1 \next_addr[17]$_DFFE_PN0P_  (.D(_0071_),
    .RN(net36),
    .CK(net1),
    .Q(net117),
    .QN(_0610_));
 DFFR_X2 \next_addr[18]$_DFFE_PN0P_  (.D(_0072_),
    .RN(net36),
    .CK(net1),
    .Q(net118),
    .QN(_0609_));
 DFFR_X1 \next_addr[19]$_DFFE_PN0P_  (.D(_0073_),
    .RN(net36),
    .CK(net1),
    .Q(net119),
    .QN(_0608_));
 DFFR_X1 \next_addr[1]$_DFFE_PN0P_  (.D(_0074_),
    .RN(net36),
    .CK(net1),
    .Q(net120),
    .QN(_0666_));
 DFFR_X2 \next_addr[20]$_DFFE_PN0P_  (.D(_0075_),
    .RN(net36),
    .CK(net1),
    .Q(net121),
    .QN(_0607_));
 DFFR_X2 \next_addr[21]$_DFFE_PN0P_  (.D(_0076_),
    .RN(net36),
    .CK(net1),
    .Q(net122),
    .QN(_0606_));
 DFFR_X2 \next_addr[22]$_DFFE_PN0P_  (.D(_0077_),
    .RN(net36),
    .CK(net1),
    .Q(net123),
    .QN(_0605_));
 DFFR_X1 \next_addr[23]$_DFFE_PN0P_  (.D(_0078_),
    .RN(net36),
    .CK(net1),
    .Q(net124),
    .QN(_0604_));
 DFFR_X1 \next_addr[24]$_DFFE_PN0P_  (.D(_0079_),
    .RN(net36),
    .CK(net1),
    .Q(net125),
    .QN(_0603_));
 DFFR_X1 \next_addr[25]$_DFFE_PN0P_  (.D(_0080_),
    .RN(net36),
    .CK(net1),
    .Q(net126),
    .QN(_0602_));
 DFFR_X2 \next_addr[26]$_DFFE_PN0P_  (.D(_0081_),
    .RN(net36),
    .CK(net1),
    .Q(net127),
    .QN(_0601_));
 DFFR_X1 \next_addr[27]$_DFFE_PN0P_  (.D(_0082_),
    .RN(net36),
    .CK(net1),
    .Q(net128),
    .QN(_0600_));
 DFFR_X1 \next_addr[28]$_DFFE_PN0P_  (.D(_0083_),
    .RN(net36),
    .CK(net1),
    .Q(net129),
    .QN(_0599_));
 DFFR_X1 \next_addr[29]$_DFFE_PN0P_  (.D(_0084_),
    .RN(net36),
    .CK(net1),
    .Q(net130),
    .QN(_0598_));
 DFFR_X1 \next_addr[2]$_DFFE_PN0P_  (.D(_0085_),
    .RN(net36),
    .CK(net1),
    .Q(net131),
    .QN(_0597_));
 DFFR_X1 \next_addr[30]$_DFFE_PN0P_  (.D(_0086_),
    .RN(net36),
    .CK(net1),
    .Q(net132),
    .QN(_0596_));
 DFFR_X1 \next_addr[31]$_DFFE_PN0P_  (.D(_0087_),
    .RN(net36),
    .CK(net1),
    .Q(net133),
    .QN(_0595_));
 DFFR_X1 \next_addr[3]$_DFFE_PN0P_  (.D(_0088_),
    .RN(net36),
    .CK(net1),
    .Q(net134),
    .QN(_0594_));
 DFFR_X1 \next_addr[4]$_DFFE_PN0P_  (.D(_0089_),
    .RN(net36),
    .CK(net1),
    .Q(net135),
    .QN(_0593_));
 DFFR_X1 \next_addr[5]$_DFFE_PN0P_  (.D(_0090_),
    .RN(net36),
    .CK(net1),
    .Q(net136),
    .QN(_0592_));
 DFFR_X1 \next_addr[6]$_DFFE_PN0P_  (.D(_0091_),
    .RN(net36),
    .CK(net1),
    .Q(net137),
    .QN(_0591_));
 DFFR_X1 \next_addr[7]$_DFFE_PN0P_  (.D(_0092_),
    .RN(net36),
    .CK(net1),
    .Q(net138),
    .QN(_0590_));
 DFFR_X1 \next_addr[8]$_DFFE_PN0P_  (.D(_0093_),
    .RN(net36),
    .CK(net1),
    .Q(net139),
    .QN(_0008_));
 DFFR_X1 \next_addr[9]$_DFFE_PN0P_  (.D(_0094_),
    .RN(net36),
    .CK(net1),
    .Q(net140),
    .QN(_0589_));
 DFFR_X1 \read_data[0]$_DFFE_PN0P_  (.D(_0095_),
    .RN(net36),
    .CK(net1),
    .Q(net183),
    .QN(_0588_));
 DFFR_X1 \read_data[10]$_DFFE_PN0P_  (.D(_0096_),
    .RN(net36),
    .CK(net1),
    .Q(net184),
    .QN(_0587_));
 DFFR_X1 \read_data[11]$_DFFE_PN0P_  (.D(_0097_),
    .RN(net36),
    .CK(net1),
    .Q(net185),
    .QN(_0586_));
 DFFR_X1 \read_data[12]$_DFFE_PN0P_  (.D(_0098_),
    .RN(net36),
    .CK(net1),
    .Q(net186),
    .QN(_0585_));
 DFFR_X1 \read_data[13]$_DFFE_PN0P_  (.D(_0099_),
    .RN(net36),
    .CK(net1),
    .Q(net187),
    .QN(_0584_));
 DFFR_X1 \read_data[14]$_DFFE_PN0P_  (.D(_0100_),
    .RN(net36),
    .CK(net1),
    .Q(net188),
    .QN(_0583_));
 DFFR_X1 \read_data[15]$_DFFE_PN0P_  (.D(_0101_),
    .RN(net36),
    .CK(net1),
    .Q(net189),
    .QN(_0582_));
 DFFR_X1 \read_data[16]$_DFFE_PN0P_  (.D(_0102_),
    .RN(net36),
    .CK(net1),
    .Q(net190),
    .QN(_0581_));
 DFFR_X1 \read_data[17]$_DFFE_PN0P_  (.D(_0103_),
    .RN(net36),
    .CK(net1),
    .Q(net191),
    .QN(_0580_));
 DFFR_X1 \read_data[18]$_DFFE_PN0P_  (.D(_0104_),
    .RN(net36),
    .CK(net1),
    .Q(net192),
    .QN(_0579_));
 DFFR_X1 \read_data[19]$_DFFE_PN0P_  (.D(_0105_),
    .RN(net36),
    .CK(net1),
    .Q(net193),
    .QN(_0578_));
 DFFR_X1 \read_data[1]$_DFFE_PN0P_  (.D(_0106_),
    .RN(net36),
    .CK(net1),
    .Q(net194),
    .QN(_0577_));
 DFFR_X1 \read_data[20]$_DFFE_PN0P_  (.D(_0107_),
    .RN(net36),
    .CK(net1),
    .Q(net195),
    .QN(_0576_));
 DFFR_X1 \read_data[21]$_DFFE_PN0P_  (.D(_0108_),
    .RN(net36),
    .CK(net1),
    .Q(net196),
    .QN(_0575_));
 DFFR_X1 \read_data[22]$_DFFE_PN0P_  (.D(_0109_),
    .RN(net36),
    .CK(net1),
    .Q(net197),
    .QN(_0574_));
 DFFR_X1 \read_data[23]$_DFFE_PN0P_  (.D(_0110_),
    .RN(net36),
    .CK(net1),
    .Q(net198),
    .QN(_0573_));
 DFFR_X1 \read_data[24]$_DFFE_PN0P_  (.D(_0111_),
    .RN(net36),
    .CK(net1),
    .Q(net199),
    .QN(_0572_));
 DFFR_X1 \read_data[25]$_DFFE_PN0P_  (.D(_0112_),
    .RN(net36),
    .CK(net1),
    .Q(net200),
    .QN(_0571_));
 DFFR_X1 \read_data[26]$_DFFE_PN0P_  (.D(_0113_),
    .RN(net36),
    .CK(net1),
    .Q(net201),
    .QN(_0570_));
 DFFR_X1 \read_data[27]$_DFFE_PN0P_  (.D(_0114_),
    .RN(net36),
    .CK(net1),
    .Q(net202),
    .QN(_0569_));
 DFFR_X1 \read_data[28]$_DFFE_PN0P_  (.D(_0115_),
    .RN(net36),
    .CK(net1),
    .Q(net203),
    .QN(_0568_));
 DFFR_X1 \read_data[29]$_DFFE_PN0P_  (.D(_0116_),
    .RN(net36),
    .CK(net1),
    .Q(net204),
    .QN(_0567_));
 DFFR_X1 \read_data[2]$_DFFE_PN0P_  (.D(_0117_),
    .RN(net36),
    .CK(net1),
    .Q(net205),
    .QN(_0566_));
 DFFR_X1 \read_data[30]$_DFFE_PN0P_  (.D(_0118_),
    .RN(net36),
    .CK(net1),
    .Q(net206),
    .QN(_0565_));
 DFFR_X1 \read_data[31]$_DFFE_PN0P_  (.D(_0119_),
    .RN(net36),
    .CK(net1),
    .Q(net207),
    .QN(_0564_));
 DFFR_X1 \read_data[3]$_DFFE_PN0P_  (.D(_0120_),
    .RN(net36),
    .CK(net1),
    .Q(net208),
    .QN(_0563_));
 DFFR_X1 \read_data[4]$_DFFE_PN0P_  (.D(_0121_),
    .RN(net36),
    .CK(net1),
    .Q(net209),
    .QN(_0562_));
 DFFR_X1 \read_data[5]$_DFFE_PN0P_  (.D(_0122_),
    .RN(net36),
    .CK(net1),
    .Q(net210),
    .QN(_0561_));
 DFFR_X1 \read_data[6]$_DFFE_PN0P_  (.D(_0123_),
    .RN(net36),
    .CK(net1),
    .Q(net211),
    .QN(_0560_));
 DFFR_X1 \read_data[7]$_DFFE_PN0P_  (.D(_0124_),
    .RN(net36),
    .CK(net1),
    .Q(net212),
    .QN(_0559_));
 DFFR_X1 \read_data[8]$_DFFE_PN0P_  (.D(_0125_),
    .RN(net36),
    .CK(net1),
    .Q(net213),
    .QN(_0558_));
 DFFR_X1 \read_data[9]$_DFFE_PN0P_  (.D(_0126_),
    .RN(net36),
    .CK(net1),
    .Q(net214),
    .QN(_0663_));
 DFFR_X1 \state[0]$_DFF_PN0_  (.D(_0552_),
    .RN(net36),
    .CK(net1),
    .Q(\state[0] ),
    .QN(_0664_));
 DFFR_X1 \state[1]$_DFF_PN0_  (.D(_0553_),
    .RN(net36),
    .CK(net1),
    .Q(\state[1] ),
    .QN(_0665_));
 DFFR_X1 \state[2]$_DFF_PN0_  (.D(_0554_),
    .RN(net36),
    .CK(net1),
    .Q(\state[2] ),
    .QN(_0000_));
 DFFR_X1 \trans_done$_DFFE_PN0P_  (.D(_0127_),
    .RN(net36),
    .CK(net1),
    .Q(net215),
    .QN(_0557_));
 DFFR_X1 \trans_resp[0]$_DFFE_PN0P_  (.D(_0128_),
    .RN(net36),
    .CK(net1),
    .Q(net216),
    .QN(_0556_));
 DFFR_X1 \trans_resp[1]$_DFFE_PN0P_  (.D(_0129_),
    .RN(net36),
    .CK(net1),
    .Q(net217),
    .QN(_0555_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_73 ();
 BUF_X16 input1 (.A(hclk),
    .Z(net1));
 BUF_X1 input2 (.A(hgrant),
    .Z(net2));
 BUF_X1 input3 (.A(hrdata[0]),
    .Z(net3));
 BUF_X1 input4 (.A(hrdata[10]),
    .Z(net4));
 BUF_X1 input5 (.A(hrdata[11]),
    .Z(net5));
 BUF_X1 input6 (.A(hrdata[12]),
    .Z(net6));
 BUF_X1 input7 (.A(hrdata[13]),
    .Z(net7));
 BUF_X1 input8 (.A(hrdata[14]),
    .Z(net8));
 BUF_X1 input9 (.A(hrdata[15]),
    .Z(net9));
 BUF_X1 input10 (.A(hrdata[16]),
    .Z(net10));
 BUF_X1 input11 (.A(hrdata[17]),
    .Z(net11));
 BUF_X1 input12 (.A(hrdata[18]),
    .Z(net12));
 BUF_X1 input13 (.A(hrdata[19]),
    .Z(net13));
 BUF_X1 input14 (.A(hrdata[1]),
    .Z(net14));
 BUF_X1 input15 (.A(hrdata[20]),
    .Z(net15));
 BUF_X1 input16 (.A(hrdata[21]),
    .Z(net16));
 BUF_X1 input17 (.A(hrdata[22]),
    .Z(net17));
 BUF_X1 input18 (.A(hrdata[23]),
    .Z(net18));
 BUF_X1 input19 (.A(hrdata[24]),
    .Z(net19));
 BUF_X1 input20 (.A(hrdata[25]),
    .Z(net20));
 BUF_X1 input21 (.A(hrdata[26]),
    .Z(net21));
 BUF_X1 input22 (.A(hrdata[27]),
    .Z(net22));
 BUF_X1 input23 (.A(hrdata[28]),
    .Z(net23));
 BUF_X1 input24 (.A(hrdata[29]),
    .Z(net24));
 BUF_X1 input25 (.A(hrdata[2]),
    .Z(net25));
 BUF_X1 input26 (.A(hrdata[30]),
    .Z(net26));
 BUF_X1 input27 (.A(hrdata[31]),
    .Z(net27));
 BUF_X1 input28 (.A(hrdata[3]),
    .Z(net28));
 BUF_X1 input29 (.A(hrdata[4]),
    .Z(net29));
 BUF_X1 input30 (.A(hrdata[5]),
    .Z(net30));
 BUF_X1 input31 (.A(hrdata[6]),
    .Z(net31));
 BUF_X1 input32 (.A(hrdata[7]),
    .Z(net32));
 BUF_X1 input33 (.A(hrdata[8]),
    .Z(net33));
 BUF_X1 input34 (.A(hrdata[9]),
    .Z(net34));
 BUF_X1 input35 (.A(hready),
    .Z(net35));
 BUF_X32 input36 (.A(hreset),
    .Z(net36));
 BUF_X1 input37 (.A(hresp[0]),
    .Z(net37));
 BUF_X1 input38 (.A(hresp[1]),
    .Z(net38));
 BUF_X1 input39 (.A(trans_addr[0]),
    .Z(net39));
 BUF_X1 input40 (.A(trans_addr[10]),
    .Z(net40));
 BUF_X1 input41 (.A(trans_addr[11]),
    .Z(net41));
 BUF_X1 input42 (.A(trans_addr[12]),
    .Z(net42));
 BUF_X1 input43 (.A(trans_addr[13]),
    .Z(net43));
 BUF_X1 input44 (.A(trans_addr[14]),
    .Z(net44));
 BUF_X1 input45 (.A(trans_addr[15]),
    .Z(net45));
 BUF_X1 input46 (.A(trans_addr[16]),
    .Z(net46));
 BUF_X1 input47 (.A(trans_addr[17]),
    .Z(net47));
 BUF_X1 input48 (.A(trans_addr[18]),
    .Z(net48));
 BUF_X1 input49 (.A(trans_addr[19]),
    .Z(net49));
 BUF_X1 input50 (.A(trans_addr[1]),
    .Z(net50));
 BUF_X1 input51 (.A(trans_addr[20]),
    .Z(net51));
 BUF_X1 input52 (.A(trans_addr[21]),
    .Z(net52));
 BUF_X1 input53 (.A(trans_addr[22]),
    .Z(net53));
 BUF_X1 input54 (.A(trans_addr[23]),
    .Z(net54));
 BUF_X1 input55 (.A(trans_addr[24]),
    .Z(net55));
 BUF_X1 input56 (.A(trans_addr[25]),
    .Z(net56));
 BUF_X1 input57 (.A(trans_addr[26]),
    .Z(net57));
 BUF_X1 input58 (.A(trans_addr[27]),
    .Z(net58));
 BUF_X1 input59 (.A(trans_addr[28]),
    .Z(net59));
 BUF_X1 input60 (.A(trans_addr[29]),
    .Z(net60));
 BUF_X1 input61 (.A(trans_addr[2]),
    .Z(net61));
 BUF_X1 input62 (.A(trans_addr[30]),
    .Z(net62));
 BUF_X1 input63 (.A(trans_addr[31]),
    .Z(net63));
 BUF_X1 input64 (.A(trans_addr[3]),
    .Z(net64));
 BUF_X1 input65 (.A(trans_addr[4]),
    .Z(net65));
 BUF_X1 input66 (.A(trans_addr[5]),
    .Z(net66));
 BUF_X1 input67 (.A(trans_addr[6]),
    .Z(net67));
 BUF_X1 input68 (.A(trans_addr[7]),
    .Z(net68));
 BUF_X1 input69 (.A(trans_addr[8]),
    .Z(net69));
 BUF_X1 input70 (.A(trans_addr[9]),
    .Z(net70));
 BUF_X1 input71 (.A(trans_burst[0]),
    .Z(net71));
 BUF_X1 input72 (.A(trans_burst[2]),
    .Z(net72));
 BUF_X1 input73 (.A(trans_size[0]),
    .Z(net73));
 BUF_X1 input74 (.A(trans_size[1]),
    .Z(net74));
 BUF_X1 input75 (.A(trans_size[2]),
    .Z(net75));
 BUF_X1 input76 (.A(trans_write),
    .Z(net76));
 BUF_X1 input77 (.A(write_data[0]),
    .Z(net77));
 BUF_X1 input78 (.A(write_data[10]),
    .Z(net78));
 BUF_X1 input79 (.A(write_data[11]),
    .Z(net79));
 BUF_X1 input80 (.A(write_data[12]),
    .Z(net80));
 BUF_X1 input81 (.A(write_data[13]),
    .Z(net81));
 BUF_X1 input82 (.A(write_data[14]),
    .Z(net82));
 BUF_X1 input83 (.A(write_data[15]),
    .Z(net83));
 BUF_X1 input84 (.A(write_data[16]),
    .Z(net84));
 BUF_X1 input85 (.A(write_data[17]),
    .Z(net85));
 BUF_X1 input86 (.A(write_data[18]),
    .Z(net86));
 BUF_X1 input87 (.A(write_data[19]),
    .Z(net87));
 BUF_X1 input88 (.A(write_data[1]),
    .Z(net88));
 BUF_X1 input89 (.A(write_data[20]),
    .Z(net89));
 BUF_X1 input90 (.A(write_data[21]),
    .Z(net90));
 BUF_X1 input91 (.A(write_data[22]),
    .Z(net91));
 BUF_X1 input92 (.A(write_data[23]),
    .Z(net92));
 BUF_X1 input93 (.A(write_data[24]),
    .Z(net93));
 BUF_X1 input94 (.A(write_data[25]),
    .Z(net94));
 BUF_X1 input95 (.A(write_data[26]),
    .Z(net95));
 BUF_X1 input96 (.A(write_data[27]),
    .Z(net96));
 BUF_X1 input97 (.A(write_data[28]),
    .Z(net97));
 BUF_X1 input98 (.A(write_data[29]),
    .Z(net98));
 BUF_X1 input99 (.A(write_data[2]),
    .Z(net99));
 BUF_X1 input100 (.A(write_data[30]),
    .Z(net100));
 BUF_X1 input101 (.A(write_data[31]),
    .Z(net101));
 BUF_X1 input102 (.A(write_data[3]),
    .Z(net102));
 BUF_X1 input103 (.A(write_data[4]),
    .Z(net103));
 BUF_X1 input104 (.A(write_data[5]),
    .Z(net104));
 BUF_X1 input105 (.A(write_data[6]),
    .Z(net105));
 BUF_X1 input106 (.A(write_data[7]),
    .Z(net106));
 BUF_X1 input107 (.A(write_data[8]),
    .Z(net107));
 BUF_X1 input108 (.A(write_data[9]),
    .Z(net108));
 BUF_X1 output109 (.A(net109),
    .Z(haddr[0]));
 BUF_X1 output110 (.A(net110),
    .Z(haddr[10]));
 BUF_X1 output111 (.A(net111),
    .Z(haddr[11]));
 BUF_X1 output112 (.A(net112),
    .Z(haddr[12]));
 BUF_X1 output113 (.A(net113),
    .Z(haddr[13]));
 BUF_X1 output114 (.A(net114),
    .Z(haddr[14]));
 BUF_X1 output115 (.A(net115),
    .Z(haddr[15]));
 BUF_X1 output116 (.A(net116),
    .Z(haddr[16]));
 BUF_X1 output117 (.A(net117),
    .Z(haddr[17]));
 BUF_X1 output118 (.A(net118),
    .Z(haddr[18]));
 BUF_X1 output119 (.A(net119),
    .Z(haddr[19]));
 BUF_X1 output120 (.A(net120),
    .Z(haddr[1]));
 BUF_X1 output121 (.A(net121),
    .Z(haddr[20]));
 BUF_X1 output122 (.A(net122),
    .Z(haddr[21]));
 BUF_X1 output123 (.A(net123),
    .Z(haddr[22]));
 BUF_X1 output124 (.A(net124),
    .Z(haddr[23]));
 BUF_X1 output125 (.A(net125),
    .Z(haddr[24]));
 BUF_X1 output126 (.A(net126),
    .Z(haddr[25]));
 BUF_X1 output127 (.A(net127),
    .Z(haddr[26]));
 BUF_X1 output128 (.A(net128),
    .Z(haddr[27]));
 BUF_X1 output129 (.A(net129),
    .Z(haddr[28]));
 BUF_X1 output130 (.A(net130),
    .Z(haddr[29]));
 BUF_X1 output131 (.A(net131),
    .Z(haddr[2]));
 BUF_X1 output132 (.A(net132),
    .Z(haddr[30]));
 BUF_X1 output133 (.A(net133),
    .Z(haddr[31]));
 BUF_X1 output134 (.A(net134),
    .Z(haddr[3]));
 BUF_X1 output135 (.A(net135),
    .Z(haddr[4]));
 BUF_X1 output136 (.A(net136),
    .Z(haddr[5]));
 BUF_X1 output137 (.A(net137),
    .Z(haddr[6]));
 BUF_X1 output138 (.A(net138),
    .Z(haddr[7]));
 BUF_X1 output139 (.A(net139),
    .Z(haddr[8]));
 BUF_X1 output140 (.A(net140),
    .Z(haddr[9]));
 BUF_X1 output141 (.A(net141),
    .Z(hburst[0]));
 BUF_X1 output142 (.A(net142),
    .Z(hburst[1]));
 BUF_X1 output143 (.A(net143),
    .Z(hburst[2]));
 BUF_X1 output144 (.A(net144),
    .Z(hbusreq));
 BUF_X1 output145 (.A(net145),
    .Z(hsize[0]));
 BUF_X1 output146 (.A(net146),
    .Z(hsize[1]));
 BUF_X1 output147 (.A(net147),
    .Z(hsize[2]));
 BUF_X1 output148 (.A(net148),
    .Z(htrans[0]));
 BUF_X1 output149 (.A(net149),
    .Z(htrans[1]));
 BUF_X1 output150 (.A(net150),
    .Z(hwdata[0]));
 BUF_X1 output151 (.A(net151),
    .Z(hwdata[10]));
 BUF_X1 output152 (.A(net152),
    .Z(hwdata[11]));
 BUF_X1 output153 (.A(net153),
    .Z(hwdata[12]));
 BUF_X1 output154 (.A(net154),
    .Z(hwdata[13]));
 BUF_X1 output155 (.A(net155),
    .Z(hwdata[14]));
 BUF_X1 output156 (.A(net156),
    .Z(hwdata[15]));
 BUF_X1 output157 (.A(net157),
    .Z(hwdata[16]));
 BUF_X1 output158 (.A(net158),
    .Z(hwdata[17]));
 BUF_X1 output159 (.A(net159),
    .Z(hwdata[18]));
 BUF_X1 output160 (.A(net160),
    .Z(hwdata[19]));
 BUF_X1 output161 (.A(net161),
    .Z(hwdata[1]));
 BUF_X1 output162 (.A(net162),
    .Z(hwdata[20]));
 BUF_X1 output163 (.A(net163),
    .Z(hwdata[21]));
 BUF_X1 output164 (.A(net164),
    .Z(hwdata[22]));
 BUF_X1 output165 (.A(net165),
    .Z(hwdata[23]));
 BUF_X1 output166 (.A(net166),
    .Z(hwdata[24]));
 BUF_X1 output167 (.A(net167),
    .Z(hwdata[25]));
 BUF_X1 output168 (.A(net168),
    .Z(hwdata[26]));
 BUF_X1 output169 (.A(net169),
    .Z(hwdata[27]));
 BUF_X1 output170 (.A(net170),
    .Z(hwdata[28]));
 BUF_X1 output171 (.A(net171),
    .Z(hwdata[29]));
 BUF_X1 output172 (.A(net172),
    .Z(hwdata[2]));
 BUF_X1 output173 (.A(net173),
    .Z(hwdata[30]));
 BUF_X1 output174 (.A(net174),
    .Z(hwdata[31]));
 BUF_X1 output175 (.A(net175),
    .Z(hwdata[3]));
 BUF_X1 output176 (.A(net176),
    .Z(hwdata[4]));
 BUF_X1 output177 (.A(net177),
    .Z(hwdata[5]));
 BUF_X1 output178 (.A(net178),
    .Z(hwdata[6]));
 BUF_X1 output179 (.A(net179),
    .Z(hwdata[7]));
 BUF_X1 output180 (.A(net180),
    .Z(hwdata[8]));
 BUF_X1 output181 (.A(net181),
    .Z(hwdata[9]));
 BUF_X1 output182 (.A(net182),
    .Z(hwrite));
 BUF_X1 output183 (.A(net183),
    .Z(read_data[0]));
 BUF_X1 output184 (.A(net184),
    .Z(read_data[10]));
 BUF_X1 output185 (.A(net185),
    .Z(read_data[11]));
 BUF_X1 output186 (.A(net186),
    .Z(read_data[12]));
 BUF_X1 output187 (.A(net187),
    .Z(read_data[13]));
 BUF_X1 output188 (.A(net188),
    .Z(read_data[14]));
 BUF_X1 output189 (.A(net189),
    .Z(read_data[15]));
 BUF_X1 output190 (.A(net190),
    .Z(read_data[16]));
 BUF_X1 output191 (.A(net191),
    .Z(read_data[17]));
 BUF_X1 output192 (.A(net192),
    .Z(read_data[18]));
 BUF_X1 output193 (.A(net193),
    .Z(read_data[19]));
 BUF_X1 output194 (.A(net194),
    .Z(read_data[1]));
 BUF_X1 output195 (.A(net195),
    .Z(read_data[20]));
 BUF_X1 output196 (.A(net196),
    .Z(read_data[21]));
 BUF_X1 output197 (.A(net197),
    .Z(read_data[22]));
 BUF_X1 output198 (.A(net198),
    .Z(read_data[23]));
 BUF_X1 output199 (.A(net199),
    .Z(read_data[24]));
 BUF_X1 output200 (.A(net200),
    .Z(read_data[25]));
 BUF_X1 output201 (.A(net201),
    .Z(read_data[26]));
 BUF_X1 output202 (.A(net202),
    .Z(read_data[27]));
 BUF_X1 output203 (.A(net203),
    .Z(read_data[28]));
 BUF_X1 output204 (.A(net204),
    .Z(read_data[29]));
 BUF_X1 output205 (.A(net205),
    .Z(read_data[2]));
 BUF_X1 output206 (.A(net206),
    .Z(read_data[30]));
 BUF_X1 output207 (.A(net207),
    .Z(read_data[31]));
 BUF_X1 output208 (.A(net208),
    .Z(read_data[3]));
 BUF_X1 output209 (.A(net209),
    .Z(read_data[4]));
 BUF_X1 output210 (.A(net210),
    .Z(read_data[5]));
 BUF_X1 output211 (.A(net211),
    .Z(read_data[6]));
 BUF_X1 output212 (.A(net212),
    .Z(read_data[7]));
 BUF_X1 output213 (.A(net213),
    .Z(read_data[8]));
 BUF_X1 output214 (.A(net214),
    .Z(read_data[9]));
 BUF_X1 output215 (.A(net215),
    .Z(trans_done));
 BUF_X1 output216 (.A(net216),
    .Z(trans_resp[0]));
 BUF_X1 output217 (.A(net217),
    .Z(trans_resp[1]));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_17 ();
 FILLCELL_X1 FILLER_0_29 ();
 FILLCELL_X16 FILLER_0_36 ();
 FILLCELL_X8 FILLER_0_52 ();
 FILLCELL_X2 FILLER_0_60 ();
 FILLCELL_X1 FILLER_0_62 ();
 FILLCELL_X8 FILLER_0_96 ();
 FILLCELL_X2 FILLER_0_110 ();
 FILLCELL_X8 FILLER_0_115 ();
 FILLCELL_X1 FILLER_0_123 ();
 FILLCELL_X32 FILLER_0_130 ();
 FILLCELL_X8 FILLER_0_162 ();
 FILLCELL_X4 FILLER_0_209 ();
 FILLCELL_X1 FILLER_0_232 ();
 FILLCELL_X4 FILLER_0_253 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X8 FILLER_1_40 ();
 FILLCELL_X2 FILLER_1_48 ();
 FILLCELL_X2 FILLER_1_70 ();
 FILLCELL_X4 FILLER_1_82 ();
 FILLCELL_X4 FILLER_1_92 ();
 FILLCELL_X32 FILLER_1_116 ();
 FILLCELL_X2 FILLER_1_148 ();
 FILLCELL_X2 FILLER_1_184 ();
 FILLCELL_X2 FILLER_1_246 ();
 FILLCELL_X1 FILLER_1_248 ();
 FILLCELL_X2 FILLER_1_272 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_53 ();
 FILLCELL_X1 FILLER_2_55 ();
 FILLCELL_X8 FILLER_2_58 ();
 FILLCELL_X2 FILLER_2_66 ();
 FILLCELL_X1 FILLER_2_68 ();
 FILLCELL_X1 FILLER_2_76 ();
 FILLCELL_X1 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_118 ();
 FILLCELL_X4 FILLER_2_150 ();
 FILLCELL_X2 FILLER_2_154 ();
 FILLCELL_X1 FILLER_2_219 ();
 FILLCELL_X8 FILLER_2_230 ();
 FILLCELL_X4 FILLER_2_238 ();
 FILLCELL_X1 FILLER_2_242 ();
 FILLCELL_X4 FILLER_2_250 ();
 FILLCELL_X1 FILLER_2_254 ();
 FILLCELL_X1 FILLER_2_258 ();
 FILLCELL_X1 FILLER_2_272 ();
 FILLCELL_X1 FILLER_2_276 ();
 FILLCELL_X2 FILLER_3_7 ();
 FILLCELL_X8 FILLER_3_36 ();
 FILLCELL_X2 FILLER_3_44 ();
 FILLCELL_X16 FILLER_3_71 ();
 FILLCELL_X4 FILLER_3_87 ();
 FILLCELL_X2 FILLER_3_91 ();
 FILLCELL_X2 FILLER_3_104 ();
 FILLCELL_X32 FILLER_3_110 ();
 FILLCELL_X8 FILLER_3_142 ();
 FILLCELL_X4 FILLER_3_150 ();
 FILLCELL_X2 FILLER_3_154 ();
 FILLCELL_X8 FILLER_3_176 ();
 FILLCELL_X4 FILLER_3_184 ();
 FILLCELL_X1 FILLER_3_188 ();
 FILLCELL_X2 FILLER_3_192 ();
 FILLCELL_X1 FILLER_3_194 ();
 FILLCELL_X1 FILLER_3_201 ();
 FILLCELL_X1 FILLER_3_205 ();
 FILLCELL_X1 FILLER_3_212 ();
 FILLCELL_X2 FILLER_3_220 ();
 FILLCELL_X4 FILLER_3_242 ();
 FILLCELL_X1 FILLER_3_276 ();
 FILLCELL_X16 FILLER_4_31 ();
 FILLCELL_X1 FILLER_4_47 ();
 FILLCELL_X4 FILLER_4_54 ();
 FILLCELL_X2 FILLER_4_58 ();
 FILLCELL_X16 FILLER_4_75 ();
 FILLCELL_X2 FILLER_4_91 ();
 FILLCELL_X1 FILLER_4_93 ();
 FILLCELL_X8 FILLER_4_101 ();
 FILLCELL_X1 FILLER_4_109 ();
 FILLCELL_X32 FILLER_4_112 ();
 FILLCELL_X32 FILLER_4_144 ();
 FILLCELL_X16 FILLER_4_176 ();
 FILLCELL_X4 FILLER_4_192 ();
 FILLCELL_X2 FILLER_4_196 ();
 FILLCELL_X1 FILLER_4_198 ();
 FILLCELL_X16 FILLER_4_219 ();
 FILLCELL_X4 FILLER_4_235 ();
 FILLCELL_X1 FILLER_4_239 ();
 FILLCELL_X2 FILLER_4_243 ();
 FILLCELL_X2 FILLER_4_272 ();
 FILLCELL_X2 FILLER_5_7 ();
 FILLCELL_X16 FILLER_5_29 ();
 FILLCELL_X4 FILLER_5_45 ();
 FILLCELL_X2 FILLER_5_49 ();
 FILLCELL_X1 FILLER_5_75 ();
 FILLCELL_X16 FILLER_5_78 ();
 FILLCELL_X8 FILLER_5_94 ();
 FILLCELL_X1 FILLER_5_113 ();
 FILLCELL_X4 FILLER_5_117 ();
 FILLCELL_X1 FILLER_5_121 ();
 FILLCELL_X32 FILLER_5_153 ();
 FILLCELL_X32 FILLER_5_185 ();
 FILLCELL_X2 FILLER_5_217 ();
 FILLCELL_X2 FILLER_5_272 ();
 FILLCELL_X16 FILLER_6_28 ();
 FILLCELL_X2 FILLER_6_44 ();
 FILLCELL_X1 FILLER_6_71 ();
 FILLCELL_X4 FILLER_6_96 ();
 FILLCELL_X1 FILLER_6_100 ();
 FILLCELL_X2 FILLER_6_105 ();
 FILLCELL_X32 FILLER_6_158 ();
 FILLCELL_X8 FILLER_6_190 ();
 FILLCELL_X4 FILLER_6_198 ();
 FILLCELL_X8 FILLER_6_207 ();
 FILLCELL_X4 FILLER_6_215 ();
 FILLCELL_X1 FILLER_6_239 ();
 FILLCELL_X2 FILLER_6_247 ();
 FILLCELL_X1 FILLER_6_249 ();
 FILLCELL_X2 FILLER_6_253 ();
 FILLCELL_X1 FILLER_6_255 ();
 FILLCELL_X2 FILLER_6_269 ();
 FILLCELL_X4 FILLER_7_4 ();
 FILLCELL_X4 FILLER_7_25 ();
 FILLCELL_X2 FILLER_7_29 ();
 FILLCELL_X1 FILLER_7_51 ();
 FILLCELL_X1 FILLER_7_64 ();
 FILLCELL_X1 FILLER_7_71 ();
 FILLCELL_X1 FILLER_7_78 ();
 FILLCELL_X8 FILLER_7_83 ();
 FILLCELL_X2 FILLER_7_91 ();
 FILLCELL_X2 FILLER_7_97 ();
 FILLCELL_X1 FILLER_7_99 ();
 FILLCELL_X2 FILLER_7_133 ();
 FILLCELL_X8 FILLER_7_137 ();
 FILLCELL_X2 FILLER_7_145 ();
 FILLCELL_X1 FILLER_7_147 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X16 FILLER_7_225 ();
 FILLCELL_X2 FILLER_7_241 ();
 FILLCELL_X1 FILLER_7_243 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_29 ();
 FILLCELL_X8 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_41 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X1 FILLER_8_59 ();
 FILLCELL_X16 FILLER_8_87 ();
 FILLCELL_X8 FILLER_8_103 ();
 FILLCELL_X2 FILLER_8_111 ();
 FILLCELL_X4 FILLER_8_116 ();
 FILLCELL_X1 FILLER_8_126 ();
 FILLCELL_X4 FILLER_8_130 ();
 FILLCELL_X8 FILLER_8_138 ();
 FILLCELL_X2 FILLER_8_146 ();
 FILLCELL_X1 FILLER_8_154 ();
 FILLCELL_X32 FILLER_8_165 ();
 FILLCELL_X32 FILLER_8_197 ();
 FILLCELL_X8 FILLER_8_229 ();
 FILLCELL_X1 FILLER_8_237 ();
 FILLCELL_X4 FILLER_8_243 ();
 FILLCELL_X1 FILLER_8_247 ();
 FILLCELL_X2 FILLER_8_275 ();
 FILLCELL_X4 FILLER_9_7 ();
 FILLCELL_X1 FILLER_9_11 ();
 FILLCELL_X8 FILLER_9_32 ();
 FILLCELL_X2 FILLER_9_40 ();
 FILLCELL_X4 FILLER_9_44 ();
 FILLCELL_X1 FILLER_9_48 ();
 FILLCELL_X1 FILLER_9_52 ();
 FILLCELL_X32 FILLER_9_87 ();
 FILLCELL_X8 FILLER_9_139 ();
 FILLCELL_X2 FILLER_9_147 ();
 FILLCELL_X1 FILLER_9_149 ();
 FILLCELL_X32 FILLER_9_181 ();
 FILLCELL_X8 FILLER_9_213 ();
 FILLCELL_X2 FILLER_9_221 ();
 FILLCELL_X1 FILLER_9_223 ();
 FILLCELL_X1 FILLER_10_13 ();
 FILLCELL_X4 FILLER_10_24 ();
 FILLCELL_X2 FILLER_10_28 ();
 FILLCELL_X4 FILLER_10_33 ();
 FILLCELL_X2 FILLER_10_37 ();
 FILLCELL_X1 FILLER_10_39 ();
 FILLCELL_X4 FILLER_10_49 ();
 FILLCELL_X2 FILLER_10_53 ();
 FILLCELL_X4 FILLER_10_59 ();
 FILLCELL_X8 FILLER_10_102 ();
 FILLCELL_X4 FILLER_10_110 ();
 FILLCELL_X2 FILLER_10_114 ();
 FILLCELL_X8 FILLER_10_141 ();
 FILLCELL_X2 FILLER_10_160 ();
 FILLCELL_X2 FILLER_10_164 ();
 FILLCELL_X32 FILLER_10_175 ();
 FILLCELL_X16 FILLER_10_207 ();
 FILLCELL_X8 FILLER_10_223 ();
 FILLCELL_X4 FILLER_10_231 ();
 FILLCELL_X2 FILLER_10_235 ();
 FILLCELL_X4 FILLER_10_244 ();
 FILLCELL_X4 FILLER_10_251 ();
 FILLCELL_X2 FILLER_10_255 ();
 FILLCELL_X1 FILLER_10_257 ();
 FILLCELL_X2 FILLER_10_265 ();
 FILLCELL_X1 FILLER_10_267 ();
 FILLCELL_X2 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_60 ();
 FILLCELL_X2 FILLER_11_69 ();
 FILLCELL_X1 FILLER_11_71 ();
 FILLCELL_X2 FILLER_11_77 ();
 FILLCELL_X1 FILLER_11_79 ();
 FILLCELL_X16 FILLER_11_86 ();
 FILLCELL_X8 FILLER_11_102 ();
 FILLCELL_X4 FILLER_11_110 ();
 FILLCELL_X1 FILLER_11_114 ();
 FILLCELL_X2 FILLER_11_144 ();
 FILLCELL_X32 FILLER_11_154 ();
 FILLCELL_X16 FILLER_11_186 ();
 FILLCELL_X8 FILLER_11_202 ();
 FILLCELL_X4 FILLER_11_210 ();
 FILLCELL_X2 FILLER_11_214 ();
 FILLCELL_X1 FILLER_11_216 ();
 FILLCELL_X1 FILLER_11_250 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_30 ();
 FILLCELL_X8 FILLER_12_46 ();
 FILLCELL_X1 FILLER_12_54 ();
 FILLCELL_X8 FILLER_12_59 ();
 FILLCELL_X2 FILLER_12_67 ();
 FILLCELL_X1 FILLER_12_69 ();
 FILLCELL_X2 FILLER_12_75 ();
 FILLCELL_X1 FILLER_12_77 ();
 FILLCELL_X4 FILLER_12_87 ();
 FILLCELL_X1 FILLER_12_91 ();
 FILLCELL_X4 FILLER_12_125 ();
 FILLCELL_X2 FILLER_12_143 ();
 FILLCELL_X1 FILLER_12_145 ();
 FILLCELL_X1 FILLER_12_154 ();
 FILLCELL_X4 FILLER_12_158 ();
 FILLCELL_X32 FILLER_12_182 ();
 FILLCELL_X16 FILLER_12_214 ();
 FILLCELL_X4 FILLER_12_230 ();
 FILLCELL_X8 FILLER_12_239 ();
 FILLCELL_X2 FILLER_12_247 ();
 FILLCELL_X1 FILLER_12_276 ();
 FILLCELL_X1 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_29 ();
 FILLCELL_X1 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_54 ();
 FILLCELL_X2 FILLER_13_62 ();
 FILLCELL_X2 FILLER_13_69 ();
 FILLCELL_X8 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_105 ();
 FILLCELL_X2 FILLER_13_109 ();
 FILLCELL_X2 FILLER_13_117 ();
 FILLCELL_X8 FILLER_13_123 ();
 FILLCELL_X8 FILLER_13_135 ();
 FILLCELL_X4 FILLER_13_143 ();
 FILLCELL_X2 FILLER_13_147 ();
 FILLCELL_X2 FILLER_13_157 ();
 FILLCELL_X32 FILLER_13_181 ();
 FILLCELL_X32 FILLER_13_213 ();
 FILLCELL_X4 FILLER_13_245 ();
 FILLCELL_X1 FILLER_13_249 ();
 FILLCELL_X4 FILLER_14_13 ();
 FILLCELL_X1 FILLER_14_17 ();
 FILLCELL_X8 FILLER_14_23 ();
 FILLCELL_X4 FILLER_14_31 ();
 FILLCELL_X2 FILLER_14_35 ();
 FILLCELL_X1 FILLER_14_44 ();
 FILLCELL_X4 FILLER_14_67 ();
 FILLCELL_X2 FILLER_14_71 ();
 FILLCELL_X1 FILLER_14_73 ();
 FILLCELL_X16 FILLER_14_93 ();
 FILLCELL_X2 FILLER_14_109 ();
 FILLCELL_X1 FILLER_14_127 ();
 FILLCELL_X4 FILLER_14_134 ();
 FILLCELL_X1 FILLER_14_138 ();
 FILLCELL_X1 FILLER_14_150 ();
 FILLCELL_X32 FILLER_14_163 ();
 FILLCELL_X16 FILLER_14_195 ();
 FILLCELL_X4 FILLER_14_211 ();
 FILLCELL_X1 FILLER_14_215 ();
 FILLCELL_X2 FILLER_14_249 ();
 FILLCELL_X1 FILLER_14_251 ();
 FILLCELL_X1 FILLER_14_258 ();
 FILLCELL_X2 FILLER_14_269 ();
 FILLCELL_X1 FILLER_15_31 ();
 FILLCELL_X16 FILLER_15_38 ();
 FILLCELL_X4 FILLER_15_54 ();
 FILLCELL_X2 FILLER_15_58 ();
 FILLCELL_X1 FILLER_15_60 ();
 FILLCELL_X1 FILLER_15_81 ();
 FILLCELL_X1 FILLER_15_92 ();
 FILLCELL_X2 FILLER_15_98 ();
 FILLCELL_X1 FILLER_15_100 ();
 FILLCELL_X1 FILLER_15_153 ();
 FILLCELL_X32 FILLER_15_185 ();
 FILLCELL_X4 FILLER_15_217 ();
 FILLCELL_X2 FILLER_15_221 ();
 FILLCELL_X1 FILLER_15_256 ();
 FILLCELL_X2 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_30 ();
 FILLCELL_X8 FILLER_16_62 ();
 FILLCELL_X4 FILLER_16_70 ();
 FILLCELL_X2 FILLER_16_74 ();
 FILLCELL_X2 FILLER_16_99 ();
 FILLCELL_X1 FILLER_16_163 ();
 FILLCELL_X32 FILLER_16_173 ();
 FILLCELL_X32 FILLER_16_205 ();
 FILLCELL_X8 FILLER_16_237 ();
 FILLCELL_X1 FILLER_16_245 ();
 FILLCELL_X1 FILLER_16_276 ();
 FILLCELL_X2 FILLER_17_4 ();
 FILLCELL_X4 FILLER_17_32 ();
 FILLCELL_X2 FILLER_17_36 ();
 FILLCELL_X32 FILLER_17_58 ();
 FILLCELL_X4 FILLER_17_90 ();
 FILLCELL_X2 FILLER_17_94 ();
 FILLCELL_X1 FILLER_17_96 ();
 FILLCELL_X4 FILLER_17_110 ();
 FILLCELL_X1 FILLER_17_119 ();
 FILLCELL_X32 FILLER_17_126 ();
 FILLCELL_X32 FILLER_17_158 ();
 FILLCELL_X32 FILLER_17_190 ();
 FILLCELL_X32 FILLER_17_222 ();
 FILLCELL_X4 FILLER_17_254 ();
 FILLCELL_X1 FILLER_17_258 ();
 FILLCELL_X2 FILLER_17_272 ();
 FILLCELL_X2 FILLER_18_4 ();
 FILLCELL_X4 FILLER_18_16 ();
 FILLCELL_X2 FILLER_18_20 ();
 FILLCELL_X1 FILLER_18_22 ();
 FILLCELL_X8 FILLER_18_29 ();
 FILLCELL_X1 FILLER_18_37 ();
 FILLCELL_X4 FILLER_18_45 ();
 FILLCELL_X2 FILLER_18_49 ();
 FILLCELL_X1 FILLER_18_51 ();
 FILLCELL_X8 FILLER_18_56 ();
 FILLCELL_X32 FILLER_18_78 ();
 FILLCELL_X4 FILLER_18_110 ();
 FILLCELL_X2 FILLER_18_114 ();
 FILLCELL_X16 FILLER_18_125 ();
 FILLCELL_X2 FILLER_18_141 ();
 FILLCELL_X32 FILLER_18_150 ();
 FILLCELL_X32 FILLER_18_182 ();
 FILLCELL_X2 FILLER_18_214 ();
 FILLCELL_X1 FILLER_18_216 ();
 FILLCELL_X2 FILLER_18_241 ();
 FILLCELL_X1 FILLER_18_243 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X16 FILLER_19_28 ();
 FILLCELL_X8 FILLER_19_44 ();
 FILLCELL_X2 FILLER_19_52 ();
 FILLCELL_X1 FILLER_19_74 ();
 FILLCELL_X2 FILLER_19_95 ();
 FILLCELL_X2 FILLER_19_107 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X8 FILLER_19_114 ();
 FILLCELL_X4 FILLER_19_122 ();
 FILLCELL_X2 FILLER_19_126 ();
 FILLCELL_X1 FILLER_19_128 ();
 FILLCELL_X32 FILLER_19_136 ();
 FILLCELL_X4 FILLER_19_168 ();
 FILLCELL_X1 FILLER_19_172 ();
 FILLCELL_X8 FILLER_19_193 ();
 FILLCELL_X1 FILLER_19_201 ();
 FILLCELL_X16 FILLER_19_230 ();
 FILLCELL_X2 FILLER_19_246 ();
 FILLCELL_X1 FILLER_19_248 ();
 FILLCELL_X2 FILLER_19_252 ();
 FILLCELL_X1 FILLER_19_254 ();
 FILLCELL_X2 FILLER_19_275 ();
 FILLCELL_X1 FILLER_20_28 ();
 FILLCELL_X16 FILLER_20_39 ();
 FILLCELL_X4 FILLER_20_55 ();
 FILLCELL_X1 FILLER_20_59 ();
 FILLCELL_X16 FILLER_20_74 ();
 FILLCELL_X1 FILLER_20_90 ();
 FILLCELL_X8 FILLER_20_104 ();
 FILLCELL_X2 FILLER_20_112 ();
 FILLCELL_X1 FILLER_20_114 ();
 FILLCELL_X4 FILLER_20_124 ();
 FILLCELL_X2 FILLER_20_128 ();
 FILLCELL_X32 FILLER_20_135 ();
 FILLCELL_X2 FILLER_20_167 ();
 FILLCELL_X8 FILLER_20_193 ();
 FILLCELL_X8 FILLER_20_224 ();
 FILLCELL_X4 FILLER_20_232 ();
 FILLCELL_X2 FILLER_20_236 ();
 FILLCELL_X8 FILLER_20_241 ();
 FILLCELL_X4 FILLER_20_249 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X1 FILLER_20_255 ();
 FILLCELL_X1 FILLER_20_276 ();
 FILLCELL_X2 FILLER_21_7 ();
 FILLCELL_X4 FILLER_21_16 ();
 FILLCELL_X1 FILLER_21_20 ();
 FILLCELL_X4 FILLER_21_24 ();
 FILLCELL_X1 FILLER_21_28 ();
 FILLCELL_X2 FILLER_21_32 ();
 FILLCELL_X1 FILLER_21_34 ();
 FILLCELL_X1 FILLER_21_59 ();
 FILLCELL_X2 FILLER_21_70 ();
 FILLCELL_X16 FILLER_21_82 ();
 FILLCELL_X2 FILLER_21_98 ();
 FILLCELL_X2 FILLER_21_110 ();
 FILLCELL_X8 FILLER_21_122 ();
 FILLCELL_X2 FILLER_21_130 ();
 FILLCELL_X16 FILLER_21_143 ();
 FILLCELL_X8 FILLER_21_159 ();
 FILLCELL_X4 FILLER_21_167 ();
 FILLCELL_X1 FILLER_21_171 ();
 FILLCELL_X1 FILLER_21_190 ();
 FILLCELL_X2 FILLER_21_194 ();
 FILLCELL_X4 FILLER_21_221 ();
 FILLCELL_X2 FILLER_21_248 ();
 FILLCELL_X1 FILLER_21_250 ();
 FILLCELL_X4 FILLER_21_260 ();
 FILLCELL_X2 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_3 ();
 FILLCELL_X1 FILLER_22_30 ();
 FILLCELL_X16 FILLER_22_41 ();
 FILLCELL_X2 FILLER_22_72 ();
 FILLCELL_X2 FILLER_22_77 ();
 FILLCELL_X1 FILLER_22_79 ();
 FILLCELL_X2 FILLER_22_95 ();
 FILLCELL_X1 FILLER_22_97 ();
 FILLCELL_X4 FILLER_22_123 ();
 FILLCELL_X1 FILLER_22_127 ();
 FILLCELL_X1 FILLER_22_148 ();
 FILLCELL_X4 FILLER_22_163 ();
 FILLCELL_X2 FILLER_22_167 ();
 FILLCELL_X1 FILLER_22_169 ();
 FILLCELL_X2 FILLER_22_174 ();
 FILLCELL_X1 FILLER_22_176 ();
 FILLCELL_X1 FILLER_22_187 ();
 FILLCELL_X8 FILLER_22_196 ();
 FILLCELL_X2 FILLER_22_204 ();
 FILLCELL_X1 FILLER_22_206 ();
 FILLCELL_X8 FILLER_22_212 ();
 FILLCELL_X4 FILLER_22_220 ();
 FILLCELL_X2 FILLER_22_224 ();
 FILLCELL_X2 FILLER_22_229 ();
 FILLCELL_X1 FILLER_22_241 ();
 FILLCELL_X1 FILLER_22_249 ();
 FILLCELL_X16 FILLER_22_253 ();
 FILLCELL_X8 FILLER_22_269 ();
 FILLCELL_X2 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_6 ();
 FILLCELL_X1 FILLER_23_8 ();
 FILLCELL_X16 FILLER_23_16 ();
 FILLCELL_X2 FILLER_23_32 ();
 FILLCELL_X1 FILLER_23_34 ();
 FILLCELL_X8 FILLER_23_55 ();
 FILLCELL_X2 FILLER_23_63 ();
 FILLCELL_X1 FILLER_23_90 ();
 FILLCELL_X1 FILLER_23_95 ();
 FILLCELL_X1 FILLER_23_115 ();
 FILLCELL_X1 FILLER_23_123 ();
 FILLCELL_X2 FILLER_23_140 ();
 FILLCELL_X1 FILLER_23_142 ();
 FILLCELL_X8 FILLER_23_155 ();
 FILLCELL_X2 FILLER_23_163 ();
 FILLCELL_X1 FILLER_23_165 ();
 FILLCELL_X16 FILLER_23_188 ();
 FILLCELL_X2 FILLER_23_204 ();
 FILLCELL_X1 FILLER_23_237 ();
 FILLCELL_X1 FILLER_23_242 ();
 FILLCELL_X4 FILLER_23_258 ();
 FILLCELL_X2 FILLER_23_262 ();
 FILLCELL_X1 FILLER_23_273 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_5 ();
 FILLCELL_X16 FILLER_24_30 ();
 FILLCELL_X4 FILLER_24_46 ();
 FILLCELL_X1 FILLER_24_50 ();
 FILLCELL_X1 FILLER_24_72 ();
 FILLCELL_X1 FILLER_24_104 ();
 FILLCELL_X1 FILLER_24_135 ();
 FILLCELL_X2 FILLER_24_141 ();
 FILLCELL_X2 FILLER_24_147 ();
 FILLCELL_X1 FILLER_24_149 ();
 FILLCELL_X16 FILLER_24_155 ();
 FILLCELL_X8 FILLER_24_171 ();
 FILLCELL_X2 FILLER_24_179 ();
 FILLCELL_X8 FILLER_24_190 ();
 FILLCELL_X4 FILLER_24_198 ();
 FILLCELL_X2 FILLER_24_202 ();
 FILLCELL_X2 FILLER_24_218 ();
 FILLCELL_X2 FILLER_24_223 ();
 FILLCELL_X1 FILLER_24_225 ();
 FILLCELL_X1 FILLER_24_230 ();
 FILLCELL_X4 FILLER_24_273 ();
 FILLCELL_X16 FILLER_25_31 ();
 FILLCELL_X2 FILLER_25_47 ();
 FILLCELL_X1 FILLER_25_78 ();
 FILLCELL_X2 FILLER_25_90 ();
 FILLCELL_X4 FILLER_25_99 ();
 FILLCELL_X2 FILLER_25_103 ();
 FILLCELL_X4 FILLER_25_111 ();
 FILLCELL_X2 FILLER_25_115 ();
 FILLCELL_X1 FILLER_25_123 ();
 FILLCELL_X4 FILLER_25_126 ();
 FILLCELL_X1 FILLER_25_130 ();
 FILLCELL_X2 FILLER_25_135 ();
 FILLCELL_X16 FILLER_25_143 ();
 FILLCELL_X4 FILLER_25_159 ();
 FILLCELL_X2 FILLER_25_163 ();
 FILLCELL_X2 FILLER_25_170 ();
 FILLCELL_X2 FILLER_25_176 ();
 FILLCELL_X1 FILLER_25_178 ();
 FILLCELL_X2 FILLER_25_183 ();
 FILLCELL_X1 FILLER_25_185 ();
 FILLCELL_X8 FILLER_25_191 ();
 FILLCELL_X4 FILLER_25_199 ();
 FILLCELL_X1 FILLER_25_203 ();
 FILLCELL_X2 FILLER_25_218 ();
 FILLCELL_X4 FILLER_26_20 ();
 FILLCELL_X1 FILLER_26_24 ();
 FILLCELL_X8 FILLER_26_28 ();
 FILLCELL_X4 FILLER_26_36 ();
 FILLCELL_X2 FILLER_26_40 ();
 FILLCELL_X2 FILLER_26_62 ();
 FILLCELL_X2 FILLER_26_66 ();
 FILLCELL_X4 FILLER_26_72 ();
 FILLCELL_X2 FILLER_26_76 ();
 FILLCELL_X1 FILLER_26_78 ();
 FILLCELL_X16 FILLER_26_101 ();
 FILLCELL_X4 FILLER_26_117 ();
 FILLCELL_X2 FILLER_26_121 ();
 FILLCELL_X4 FILLER_26_129 ();
 FILLCELL_X1 FILLER_26_133 ();
 FILLCELL_X16 FILLER_26_145 ();
 FILLCELL_X2 FILLER_26_161 ();
 FILLCELL_X1 FILLER_26_163 ();
 FILLCELL_X16 FILLER_26_189 ();
 FILLCELL_X2 FILLER_26_205 ();
 FILLCELL_X1 FILLER_26_207 ();
 FILLCELL_X2 FILLER_26_226 ();
 FILLCELL_X2 FILLER_27_4 ();
 FILLCELL_X1 FILLER_27_6 ();
 FILLCELL_X32 FILLER_27_37 ();
 FILLCELL_X8 FILLER_27_69 ();
 FILLCELL_X4 FILLER_27_77 ();
 FILLCELL_X2 FILLER_27_81 ();
 FILLCELL_X1 FILLER_27_83 ();
 FILLCELL_X1 FILLER_27_87 ();
 FILLCELL_X16 FILLER_27_98 ();
 FILLCELL_X2 FILLER_27_114 ();
 FILLCELL_X1 FILLER_27_116 ();
 FILLCELL_X8 FILLER_27_123 ();
 FILLCELL_X4 FILLER_27_131 ();
 FILLCELL_X1 FILLER_27_155 ();
 FILLCELL_X4 FILLER_27_163 ();
 FILLCELL_X2 FILLER_27_167 ();
 FILLCELL_X1 FILLER_27_169 ();
 FILLCELL_X4 FILLER_27_173 ();
 FILLCELL_X2 FILLER_27_182 ();
 FILLCELL_X16 FILLER_27_186 ();
 FILLCELL_X4 FILLER_27_202 ();
 FILLCELL_X1 FILLER_27_206 ();
 FILLCELL_X4 FILLER_27_225 ();
 FILLCELL_X2 FILLER_27_275 ();
 FILLCELL_X1 FILLER_28_13 ();
 FILLCELL_X16 FILLER_28_37 ();
 FILLCELL_X8 FILLER_28_53 ();
 FILLCELL_X4 FILLER_28_61 ();
 FILLCELL_X1 FILLER_28_65 ();
 FILLCELL_X8 FILLER_28_80 ();
 FILLCELL_X8 FILLER_28_102 ();
 FILLCELL_X1 FILLER_28_110 ();
 FILLCELL_X8 FILLER_28_131 ();
 FILLCELL_X2 FILLER_28_139 ();
 FILLCELL_X2 FILLER_28_152 ();
 FILLCELL_X8 FILLER_28_158 ();
 FILLCELL_X2 FILLER_28_166 ();
 FILLCELL_X16 FILLER_28_181 ();
 FILLCELL_X8 FILLER_28_197 ();
 FILLCELL_X4 FILLER_28_205 ();
 FILLCELL_X2 FILLER_28_209 ();
 FILLCELL_X4 FILLER_28_227 ();
 FILLCELL_X2 FILLER_28_231 ();
 FILLCELL_X1 FILLER_28_233 ();
 FILLCELL_X2 FILLER_28_255 ();
 FILLCELL_X1 FILLER_28_257 ();
 FILLCELL_X2 FILLER_28_261 ();
 FILLCELL_X1 FILLER_28_263 ();
 FILLCELL_X1 FILLER_28_267 ();
 FILLCELL_X2 FILLER_29_34 ();
 FILLCELL_X1 FILLER_29_36 ();
 FILLCELL_X16 FILLER_29_40 ();
 FILLCELL_X8 FILLER_29_56 ();
 FILLCELL_X1 FILLER_29_64 ();
 FILLCELL_X16 FILLER_29_111 ();
 FILLCELL_X8 FILLER_29_127 ();
 FILLCELL_X16 FILLER_29_139 ();
 FILLCELL_X4 FILLER_29_155 ();
 FILLCELL_X1 FILLER_29_190 ();
 FILLCELL_X1 FILLER_29_195 ();
 FILLCELL_X1 FILLER_29_201 ();
 FILLCELL_X4 FILLER_29_217 ();
 FILLCELL_X1 FILLER_29_221 ();
 FILLCELL_X2 FILLER_29_227 ();
 FILLCELL_X16 FILLER_30_34 ();
 FILLCELL_X8 FILLER_30_50 ();
 FILLCELL_X4 FILLER_30_58 ();
 FILLCELL_X1 FILLER_30_62 ();
 FILLCELL_X8 FILLER_30_75 ();
 FILLCELL_X4 FILLER_30_83 ();
 FILLCELL_X2 FILLER_30_87 ();
 FILLCELL_X1 FILLER_30_89 ();
 FILLCELL_X4 FILLER_30_100 ();
 FILLCELL_X16 FILLER_30_107 ();
 FILLCELL_X2 FILLER_30_123 ();
 FILLCELL_X16 FILLER_30_151 ();
 FILLCELL_X8 FILLER_30_167 ();
 FILLCELL_X1 FILLER_30_175 ();
 FILLCELL_X1 FILLER_30_184 ();
 FILLCELL_X2 FILLER_30_189 ();
 FILLCELL_X1 FILLER_30_195 ();
 FILLCELL_X2 FILLER_30_201 ();
 FILLCELL_X2 FILLER_30_208 ();
 FILLCELL_X1 FILLER_30_210 ();
 FILLCELL_X1 FILLER_30_221 ();
 FILLCELL_X16 FILLER_30_228 ();
 FILLCELL_X1 FILLER_30_244 ();
 FILLCELL_X16 FILLER_30_253 ();
 FILLCELL_X8 FILLER_30_269 ();
 FILLCELL_X32 FILLER_31_17 ();
 FILLCELL_X32 FILLER_31_49 ();
 FILLCELL_X1 FILLER_31_81 ();
 FILLCELL_X4 FILLER_31_110 ();
 FILLCELL_X2 FILLER_31_114 ();
 FILLCELL_X1 FILLER_31_116 ();
 FILLCELL_X4 FILLER_31_159 ();
 FILLCELL_X2 FILLER_31_163 ();
 FILLCELL_X2 FILLER_31_172 ();
 FILLCELL_X1 FILLER_31_187 ();
 FILLCELL_X1 FILLER_31_193 ();
 FILLCELL_X2 FILLER_31_199 ();
 FILLCELL_X2 FILLER_31_221 ();
 FILLCELL_X1 FILLER_31_236 ();
 FILLCELL_X2 FILLER_31_241 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_3 ();
 FILLCELL_X32 FILLER_32_34 ();
 FILLCELL_X32 FILLER_32_66 ();
 FILLCELL_X2 FILLER_32_98 ();
 FILLCELL_X8 FILLER_32_111 ();
 FILLCELL_X4 FILLER_32_119 ();
 FILLCELL_X2 FILLER_32_123 ();
 FILLCELL_X2 FILLER_32_127 ();
 FILLCELL_X1 FILLER_32_129 ();
 FILLCELL_X1 FILLER_32_139 ();
 FILLCELL_X2 FILLER_32_144 ();
 FILLCELL_X1 FILLER_32_156 ();
 FILLCELL_X1 FILLER_32_160 ();
 FILLCELL_X2 FILLER_32_165 ();
 FILLCELL_X2 FILLER_32_169 ();
 FILLCELL_X1 FILLER_32_185 ();
 FILLCELL_X4 FILLER_32_189 ();
 FILLCELL_X4 FILLER_32_199 ();
 FILLCELL_X1 FILLER_32_211 ();
 FILLCELL_X8 FILLER_32_240 ();
 FILLCELL_X2 FILLER_32_248 ();
 FILLCELL_X16 FILLER_32_260 ();
 FILLCELL_X1 FILLER_32_276 ();
 FILLCELL_X1 FILLER_33_1 ();
 FILLCELL_X4 FILLER_33_22 ();
 FILLCELL_X4 FILLER_33_46 ();
 FILLCELL_X2 FILLER_33_50 ();
 FILLCELL_X16 FILLER_33_72 ();
 FILLCELL_X4 FILLER_33_88 ();
 FILLCELL_X8 FILLER_33_112 ();
 FILLCELL_X4 FILLER_33_120 ();
 FILLCELL_X2 FILLER_33_124 ();
 FILLCELL_X2 FILLER_33_130 ();
 FILLCELL_X1 FILLER_33_137 ();
 FILLCELL_X1 FILLER_33_144 ();
 FILLCELL_X4 FILLER_33_149 ();
 FILLCELL_X2 FILLER_33_153 ();
 FILLCELL_X8 FILLER_33_174 ();
 FILLCELL_X1 FILLER_33_182 ();
 FILLCELL_X1 FILLER_33_202 ();
 FILLCELL_X2 FILLER_33_235 ();
 FILLCELL_X1 FILLER_33_237 ();
 FILLCELL_X16 FILLER_33_258 ();
 FILLCELL_X2 FILLER_33_274 ();
 FILLCELL_X1 FILLER_33_276 ();
 FILLCELL_X4 FILLER_34_17 ();
 FILLCELL_X4 FILLER_34_27 ();
 FILLCELL_X2 FILLER_34_31 ();
 FILLCELL_X4 FILLER_34_40 ();
 FILLCELL_X2 FILLER_34_44 ();
 FILLCELL_X1 FILLER_34_46 ();
 FILLCELL_X1 FILLER_34_54 ();
 FILLCELL_X2 FILLER_34_75 ();
 FILLCELL_X16 FILLER_34_97 ();
 FILLCELL_X8 FILLER_34_133 ();
 FILLCELL_X1 FILLER_34_141 ();
 FILLCELL_X4 FILLER_34_146 ();
 FILLCELL_X2 FILLER_34_150 ();
 FILLCELL_X8 FILLER_34_176 ();
 FILLCELL_X2 FILLER_34_184 ();
 FILLCELL_X1 FILLER_34_186 ();
 FILLCELL_X4 FILLER_34_194 ();
 FILLCELL_X2 FILLER_34_225 ();
 FILLCELL_X16 FILLER_34_252 ();
 FILLCELL_X8 FILLER_34_268 ();
 FILLCELL_X1 FILLER_34_276 ();
 FILLCELL_X1 FILLER_35_69 ();
 FILLCELL_X1 FILLER_35_73 ();
 FILLCELL_X2 FILLER_35_81 ();
 FILLCELL_X16 FILLER_35_103 ();
 FILLCELL_X2 FILLER_35_119 ();
 FILLCELL_X1 FILLER_35_144 ();
 FILLCELL_X8 FILLER_35_216 ();
 FILLCELL_X4 FILLER_35_224 ();
 FILLCELL_X16 FILLER_35_255 ();
 FILLCELL_X4 FILLER_35_271 ();
 FILLCELL_X2 FILLER_35_275 ();
 FILLCELL_X2 FILLER_36_34 ();
 FILLCELL_X1 FILLER_36_39 ();
 FILLCELL_X1 FILLER_36_81 ();
 FILLCELL_X2 FILLER_36_89 ();
 FILLCELL_X2 FILLER_36_94 ();
 FILLCELL_X2 FILLER_36_99 ();
 FILLCELL_X8 FILLER_36_110 ();
 FILLCELL_X4 FILLER_36_118 ();
 FILLCELL_X2 FILLER_36_122 ();
 FILLCELL_X2 FILLER_36_133 ();
 FILLCELL_X1 FILLER_36_135 ();
 FILLCELL_X8 FILLER_36_157 ();
 FILLCELL_X2 FILLER_36_192 ();
 FILLCELL_X1 FILLER_36_194 ();
 FILLCELL_X4 FILLER_36_198 ();
 FILLCELL_X1 FILLER_36_202 ();
 FILLCELL_X4 FILLER_36_209 ();
 FILLCELL_X2 FILLER_36_213 ();
 FILLCELL_X1 FILLER_36_215 ();
 FILLCELL_X1 FILLER_36_222 ();
 FILLCELL_X4 FILLER_36_226 ();
 FILLCELL_X8 FILLER_36_233 ();
 FILLCELL_X1 FILLER_36_241 ();
 FILLCELL_X32 FILLER_36_245 ();
endmodule
