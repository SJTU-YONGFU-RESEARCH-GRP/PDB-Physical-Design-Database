module johnson_counter (clk,
    enable,
    load_en,
    rst_n,
    count,
    load_val);
 input clk;
 input enable;
 input load_en;
 input rst_n;
 output [3:0] count;
 input [3:0] load_val;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net12;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _09_ (.I(net11),
    .ZN(_04_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _10_ (.I0(_04_),
    .I1(net4),
    .S(net3),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11_ (.I0(net8),
    .I1(_05_),
    .S(net2),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12_ (.I0(net8),
    .I1(net5),
    .S(net3),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13_ (.I0(net9),
    .I1(_06_),
    .S(net2),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14_ (.I0(net9),
    .I1(net6),
    .S(net3),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15_ (.I0(net10),
    .I1(_07_),
    .S(net2),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16_ (.I0(net10),
    .I1(net7),
    .S(net3),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17_ (.I0(net11),
    .I1(_08_),
    .S(net2),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \count[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 hold1 (.I(net12),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input2 (.I(load_en),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(load_val[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(load_val[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(load_val[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(load_val[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output7 (.I(net8),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net9),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net10),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net11),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_212 ();
endmodule
