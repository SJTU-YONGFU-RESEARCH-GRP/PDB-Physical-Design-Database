
* cell fwft_fifo
* pin wr_data[3]
* pin NWELL
* pin PWELL
* pin wr_data[4]
* pin wr_data[2]
* pin wr_data[5]
* pin wr_data[1]
* pin wr_data[7]
* pin clk
* pin rd_data[5]
* pin rd_data[7]
* pin rd_data[1]
* pin wr_data[6]
* pin rd_data[6]
* pin rd_data[0]
* pin rd_data[2]
* pin rd_data[3]
* pin rd_data[4]
* pin full
* pin empty
* pin rst_n
* pin rd_en
* pin wr_data[0]
* pin wr_en
* pin data_count[0]
* pin data_count[3]
* pin data_count[2]
* pin almost_empty
* pin almost_full
* pin data_count[1]
* pin data_count[4]
.SUBCKT fwft_fifo 1 2 3 49 58 192 235 290 360 424 425 426 434 474 475 494 495
+ 496 508 515 525 542 582 643 676 677 678 679 680 681 682
* net 1 wr_data[3]
* net 2 NWELL
* net 3 PWELL
* net 49 wr_data[4]
* net 58 wr_data[2]
* net 192 wr_data[5]
* net 235 wr_data[1]
* net 290 wr_data[7]
* net 360 clk
* net 424 rd_data[5]
* net 425 rd_data[7]
* net 426 rd_data[1]
* net 434 wr_data[6]
* net 474 rd_data[6]
* net 475 rd_data[0]
* net 494 rd_data[2]
* net 495 rd_data[3]
* net 496 rd_data[4]
* net 508 full
* net 515 empty
* net 525 rst_n
* net 542 rd_en
* net 582 wr_data[0]
* net 643 wr_en
* net 676 data_count[0]
* net 677 data_count[3]
* net 678 data_count[2]
* net 679 almost_empty
* net 680 almost_full
* net 681 data_count[1]
* net 682 data_count[4]
* cell instance $5 m0 *1 250.04,217
X$5 1 3 2 8 CLKBUF_X2
* cell instance $7 r0 *1 268.28,295.4
X$7 540 592 3 2 594 NOR2_X1
* cell instance $55 r0 *1 247.95,295.4
X$55 513 549 3 2 588 NAND2_X1
* cell instance $59 m0 *1 247.76,298.2
X$59 588 466 580 3 622 2 AOI21_X1
* cell instance $60 m0 *1 248.52,298.2
X$60 503 540 3 2 601 NOR2_X1
* cell instance $62 m0 *1 249.47,298.2
X$62 602 3 2 580 CLKBUF_X3
* cell instance $64 r0 *1 249.66,295.4
X$64 3 467 2 602 BUF_X8
* cell instance $72 m0 *1 255.36,298.2
X$72 576 577 603 3 2 609 MUX2_X1
* cell instance $73 r0 *1 255.74,295.4
X$73 454 603 2 3 589 AND2_X1
* cell instance $75 r0 *1 256.5,295.4
X$75 586 561 589 3 2 590 MUX2_X1
* cell instance $81 m0 *1 256.88,298.2
X$81 3 590 511 603 612 2 DFF_X2
* cell instance $83 m0 *1 262.01,298.2
X$83 591 526 580 3 604 2 AOI21_X1
* cell instance $84 m0 *1 262.77,298.2
X$84 578 605 576 565 3 2 591 NAND4_X1
* cell instance $86 m0 *1 266.76,298.2
X$86 616 526 580 3 608 2 AOI21_X1
* cell instance $88 m0 *1 267.9,298.2
X$88 592 543 2 3 593 AND2_X1
* cell instance $89 m0 *1 268.66,298.2
X$89 593 608 594 3 2 607 MUX2_X1
* cell instance $90 m0 *1 269.99,298.2
X$90 3 742 606 607 507 2 DFF_X1
* cell instance $148 r0 *1 244.72,513.8
X$148 665 3 2 676 BUF_X1
* cell instance $150 r0 *1 245.29,513.8
X$150 666 3 2 678 BUF_X1
* cell instance $151 r0 *1 245.86,513.8
X$151 674 3 2 680 BUF_X1
* cell instance $155 r0 *1 251.75,513.8
X$155 672 3 2 681 BUF_X1
* cell instance $160 r0 *1 266.19,513.8
X$160 466 3 2 682 BUF_X1
* cell instance $836 r0 *1 262.39,242.2
X$836 121 181 3 2 182 OR2_X1
* cell instance $837 r0 *1 263.15,242.2
X$837 195 160 196 179 2 3 181 OAI22_X1
* cell instance $839 r0 *1 264.29,242.2
X$839 177 46 199 3 2 175 MUX2_X1
* cell instance $842 r0 *1 268.85,242.2
X$842 178 46 220 3 2 179 MUX2_X1
* cell instance $862 r0 *1 256.69,242.2
X$862 159 46 174 3 2 173 MUX2_X1
* cell instance $865 m0 *1 256.69,245
X$865 195 161 196 173 2 3 186 OAI22_X1
* cell instance $866 m0 *1 257.64,245
X$866 81 186 3 2 197 OR2_X1
* cell instance $870 m0 *1 261.06,245
X$870 143 3 2 848 INV_X1
* cell instance $871 m0 *1 261.44,245
X$871 195 184 196 175 2 3 205 OAI22_X1
* cell instance $872 m0 *1 262.39,245
X$872 105 3 2 143 CLKBUF_X3
* cell instance $873 m0 *1 263.34,245
X$873 85 205 3 2 201 OR2_X1
* cell instance $2925 m0 *1 244.91,513.8
X$2925 673 3 2 677 BUF_X1
* cell instance $2928 m0 *1 246.05,513.8
X$2928 683 3 2 679 BUF_X1
* cell instance $9437 m0 *1 242.06,306.6
X$9437 3 701 648 640 463 2 DFF_X1
* cell instance $9439 m0 *1 245.29,306.6
X$9439 648 2 536 3 BUF_X4
* cell instance $9441 m0 *1 247.38,306.6
X$9441 642 655 2 3 651 AND2_X1
* cell instance $9443 m0 *1 248.52,306.6
X$9443 3 574 649 672 636 646 2 FA_X1
* cell instance $9444 r0 *1 248.9,303.8
X$9444 645 611 642 2 3 650 HA_X1
* cell instance $9448 r0 *1 254.22,303.8
X$9448 3 560 523 646 578 2 DFF_X2
* cell instance $9452 m0 *1 258.21,306.6
X$9452 3 709 652 644 511 2 DFF_X1
* cell instance $9455 r0 *1 260.49,303.8
X$9455 605 627 3 2 644 XOR2_X1
* cell instance $9456 m0 *1 261.44,306.6
X$9456 652 3 2 605 BUF_X2
* cell instance $9460 m0 *1 262.39,306.6
X$9460 3 731 653 639 511 2 DFF_X1
* cell instance $9462 r0 *1 262.96,303.8
X$9462 623 637 3 2 639 XOR2_X1
* cell instance $9465 r0 *1 265.24,303.8
X$9465 653 3 2 623 BUF_X1
* cell instance $9680 r0 *1 247.19,309.4
X$9680 642 649 3 2 659 XNOR2_X2
* cell instance $9900 m0 *1 244.53,315
X$9900 656 658 2 670 3 XOR2_X2
* cell instance $9903 r0 *1 245.67,312.2
X$9903 669 657 656 2 3 548 MUX2_X2
* cell instance $9904 m0 *1 246.24,315
X$9904 659 3 2 666 INV_X4
* cell instance $9905 m0 *1 247.19,315
X$9905 659 668 641 658 3 2 669 NAND4_X1
* cell instance $9906 r0 *1 247.38,312.2
X$9906 658 641 668 659 2 3 661 AND4_X1
* cell instance $9907 m0 *1 248.14,315
X$9907 667 3 2 668 INV_X1
* cell instance $9908 r0 *1 248.52,312.2
X$9908 661 663 656 2 3 602 MUX2_X2
* cell instance $10335 r0 *1 229.71,289.8
X$10335 3 781 546 568 463 2 DFF_X1
* cell instance $10339 m0 *1 234.08,292.6
X$10339 582 3 2 438 CLKBUF_X2
* cell instance $10346 r0 *1 243.58,289.8
X$10346 549 3 2 535 INV_X4
* cell instance $10349 r0 *1 245.67,289.8
X$10349 547 522 548 2 3 115 OAI21_X4
* cell instance $10351 r0 *1 248.14,289.8
X$10351 3 521 2 548 BUF_X8
* cell instance $10356 r0 *1 254.41,289.8
X$10356 3 787 559 560 523 2 DFF_X1
* cell instance $10357 m0 *1 254.6,292.6
X$10357 566 467 522 3 561 2 AOI21_X2
* cell instance $10359 m0 *1 256.31,292.6
X$10359 586 561 562 3 2 524 MUX2_X1
* cell instance $10364 r0 *1 262.58,289.8
X$10364 3 751 564 539 511 2 DFF_X1
* cell instance $10367 m0 *1 265.43,292.6
X$10367 564 543 2 3 570 AND2_X1
* cell instance $10368 r0 *1 265.81,289.8
X$10368 540 564 3 2 552 NOR2_X1
* cell instance $10369 m0 *1 266.19,292.6
X$10369 565 3 2 566 INV_X1
* cell instance $10372 r0 *1 266.57,289.8
X$10372 567 566 3 2 553 NAND2_X1
* cell instance $10373 r0 *1 267.14,289.8
X$10373 540 553 554 3 558 2 AOI21_X1
* cell instance $10375 m0 *1 267.71,292.6
X$10375 569 565 567 3 581 2 AOI21_X2
* cell instance $10376 r0 *1 267.9,289.8
X$10376 555 3 2 540 INV_X2
* cell instance $10377 r0 *1 268.47,289.8
X$10377 3 558 507 556 567 2 DFF_X2
* cell instance $10381 r0 *1 274.36,289.8
X$10381 542 3 2 565 BUF_X2
* cell instance $20192 r0 *1 244.53,317.8
X$20192 526 670 671 2 3 674 OAI21_X4
* cell instance $20193 m0 *1 244.72,320.6
X$20193 670 3 2 673 INV_X2
* cell instance $21056 m0 *1 230.66,281.4
X$21056 438 52 462 3 2 476 MUX2_X1
* cell instance $21057 m0 *1 231.99,281.4
X$21057 3 724 462 476 463 2 DFF_X1
* cell instance $21068 r0 *1 243.01,278.6
X$21068 3 39 465 466 467 2 AOI21_X4
* cell instance $21069 m0 *1 243.01,281.4
X$21069 3 187 488 466 467 2 AOI21_X4
* cell instance $21073 m0 *1 248.9,281.4
X$21073 3 132 482 469 467 2 AOI21_X4
* cell instance $21080 m0 *1 266.57,281.4
X$21080 445 472 446 3 2 486 NAND3_X1
* cell instance $21081 m0 *1 267.33,281.4
X$21081 444 182 486 487 447 2 3 471 OAI221_X1
* cell instance $21082 m0 *1 268.47,281.4
X$21082 472 454 3 2 487 NAND2_X1
* cell instance $21087 m0 *1 273.22,281.4
X$21087 444 197 492 499 447 2 3 484 OAI221_X1
* cell instance $26549 m0 *1 234.08,222.6
X$26549 3 743 36 20 9 2 DFF_X1
* cell instance $26554 m0 *1 241.3,222.6
X$26554 3 741 10 19 4 2 DFF_X1
* cell instance $26558 m0 *1 247.76,222.6
X$26558 3 740 33 17 4 2 DFF_X1
* cell instance $26564 m0 *1 255.74,222.6
X$26564 5 26 7 3 2 16 MUX2_X1
* cell instance $26565 m0 *1 257.07,222.6
X$26565 3 706 5 16 11 2 DFF_X1
* cell instance $26570 m0 *1 261.63,222.6
X$26570 3 726 12 6 11 2 DFF_X1
* cell instance $26573 m0 *1 265.43,222.6
X$26573 13 15 7 3 2 14 MUX2_X1
* cell instance $30534 m0 *1 244.91,511
X$30534 675 466 666 673 3 2 683 NOR4_X1
* cell instance $35095 r0 *1 230.09,275.8
X$35095 438 125 437 3 2 448 MUX2_X1
* cell instance $35096 r0 *1 231.42,275.8
X$35096 438 115 439 3 2 449 MUX2_X1
* cell instance $35120 m0 *1 233.7,278.6
X$35120 3 722 450 477 389 2 DFF_X1
* cell instance $35121 r0 *1 234.65,275.8
X$35121 450 213 381 3 2 477 MUX2_X1
* cell instance $35122 r0 *1 233.89,275.8
X$35122 438 3 2 381 BUF_X2
* cell instance $35123 r0 *1 235.98,275.8
X$35123 3 815 416 478 389 2 DFF_X1
* cell instance $35126 m0 *1 236.93,278.6
X$35126 416 187 381 3 2 478 MUX2_X1
* cell instance $35129 r0 *1 240.54,275.8
X$35129 105 3 2 389 CLKBUF_X3
* cell instance $35131 r0 *1 241.49,275.8
X$35131 389 3 2 846 INV_X4
* cell instance $35139 m0 *1 242.82,278.6
X$35139 3 213 464 466 467 2 AOI21_X4
* cell instance $35140 r0 *1 245.29,275.8
X$35140 3 15 479 469 467 2 AOI21_X4
* cell instance $35142 r0 *1 247.76,275.8
X$35142 105 3 2 330 CLKBUF_X3
* cell instance $35143 r0 *1 248.71,275.8
X$35143 330 3 2 841 INV_X2
* cell instance $35147 r0 *1 253.27,275.8
X$35147 3 789 417 455 330 2 DFF_X1
* cell instance $35148 r0 *1 256.5,275.8
X$35148 3 774 440 485 314 2 DFF_X1
* cell instance $35149 r0 *1 259.73,275.8
X$35149 440 217 381 3 2 485 MUX2_X1
* cell instance $35150 r0 *1 261.06,275.8
X$35150 3 794 458 441 314 2 DFF_X1
* cell instance $35154 r0 *1 266.76,275.8
X$35154 445 442 446 3 2 443 NAND3_X1
* cell instance $35155 r0 *1 267.52,275.8
X$35155 3 421 314 835 442 2 DFF_X2
* cell instance $35156 r0 *1 271.13,275.8
X$35156 430 454 3 2 431 NAND2_X1
* cell instance $35159 r0 *1 272.65,275.8
X$35159 445 422 446 3 2 456 NAND3_X1
* cell instance $35160 r0 *1 273.41,275.8
X$35160 422 454 3 2 453 NAND2_X1
* cell instance $35162 m0 *1 245.29,278.6
X$35162 3 30 468 469 467 2 AOI21_X4
* cell instance $35168 m0 *1 253.65,278.6
X$35168 3 715 470 483 330 2 DFF_X1
* cell instance $35169 m0 *1 256.88,278.6
X$35169 470 132 381 3 2 483 MUX2_X1
* cell instance $35173 r0 *1 275.5,275.8
X$35173 445 473 446 3 2 481 NAND3_X1
* cell instance $35174 r0 *1 274.36,275.8
X$35174 407 444 481 451 447 2 3 480 OAI221_X1
* cell instance $35175 r0 *1 276.26,275.8
X$35175 473 446 3 2 451 NAND2_X1
* cell instance $35176 r0 *1 276.83,275.8
X$35176 3 480 320 833 473 2 DFF_X2
* cell instance $35261 r0 *1 510.53,275.8
X$35261 442 3 2 474 BUF_X1
* cell instance $35262 r0 *1 511.86,275.8
X$35262 473 3 2 475 BUF_X1
* cell instance $35401 r0 *1 226.67,287
X$35401 3 779 534 527 463 2 DFF_X1
* cell instance $35405 r0 *1 231.61,287
X$35405 534 340 546 3 2 529 MUX2_X1
* cell instance $35412 m0 *1 230.66,289.8
X$35412 438 110 546 3 2 568 MUX2_X1
* cell instance $35415 m0 *1 235.41,289.8
X$35415 557 522 521 2 3 110 OAI21_X4
* cell instance $35418 r0 *1 237.88,287
X$35418 532 522 521 2 3 108 OAI21_X4
* cell instance $35419 r0 *1 240.54,287
X$35419 105 3 2 463 CLKBUF_X3
* cell instance $35420 r0 *1 241.49,287
X$35420 536 535 505 3 2 NOR2_X4
* cell instance $35421 r0 *1 243.2,287
X$35421 3 535 536 506 538 544 2 NOR4_X4
* cell instance $35422 r0 *1 246.62,287
X$35422 545 537 503 2 533 3 NOR3_X2
* cell instance $35423 r0 *1 247.95,287
X$35423 512 3 2 538 INV_X1
* cell instance $35424 r0 *1 248.33,287
X$35424 545 538 503 2 519 3 NOR3_X2
* cell instance $35425 r0 *1 249.66,287
X$35425 105 3 2 523 CLKBUF_X3
* cell instance $35426 r0 *1 250.61,287
X$35426 550 3 2 469 INV_X4
* cell instance $35434 m0 *1 241.49,289.8
X$35434 3 535 536 506 537 557 2 NOR4_X4
* cell instance $35436 m0 *1 245.1,289.8
X$35436 506 489 501 2 3 547 AND3_X1
* cell instance $35438 m0 *1 246.24,289.8
X$35438 549 536 2 3 501 AND2_X2
* cell instance $35440 m0 *1 247.57,289.8
X$35440 536 549 3 2 545 NAND2_X1
* cell instance $35443 m0 *1 250.42,289.8
X$35443 3 522 2 550 BUF_X8
* cell instance $35446 m0 *1 253.46,289.8
X$35446 522 2 526 3 BUF_X4
* cell instance $35455 m0 *1 256.69,289.8
X$35455 559 2 340 3 BUF_X4
* cell instance $35459 m0 *1 264.67,289.8
X$35459 570 217 552 3 2 539 MUX2_X1
* cell instance $35460 r0 *1 265.81,287
X$35460 511 3 2 847 INV_X4
* cell instance $35461 r0 *1 264.86,287
X$35461 105 3 2 511 CLKBUF_X3
* cell instance $35462 r0 *1 266.76,287
X$35462 445 540 3 2 528 NOR2_X1
* cell instance $35464 r0 *1 267.52,287
X$35464 543 3 2 446 BUF_X2
* cell instance $35465 r0 *1 268.28,287
X$35465 445 3 2 541 INV_X1
* cell instance $35470 m0 *1 267.14,289.8
X$35470 466 521 541 2 554 3 OAI21_X1
* cell instance $35472 m0 *1 268.28,289.8
X$35472 555 3 2 543 BUF_X2
* cell instance $35474 m0 *1 269.23,289.8
X$35474 555 556 3 2 569 NAND2_X1
* cell instance $35475 m0 *1 269.8,289.8
X$35475 3 445 556 565 567 2 AOI21_X4
* cell instance $35476 r0 *1 272.27,287
X$35476 525 3 2 555 BUF_X1
* cell instance $35521 r0 *1 514.14,287
X$35521 556 3 2 515 BUF_X1
* cell instance $35525 m0 *1 272.46,289.8
X$35525 555 3 2 454 CLKBUF_X3
* cell instance $35692 m0 *1 228,287
X$35692 438 108 534 3 2 527 MUX2_X1
* cell instance $35696 r0 *1 235.6,284.2
X$35696 518 522 521 2 3 52 OAI21_X4
* cell instance $35698 r0 *1 239.78,284.2
X$35698 531 522 521 2 3 125 OAI21_X4
* cell instance $35700 m0 *1 235.6,287
X$35700 544 522 521 2 3 57 OAI21_X4
* cell instance $35704 m0 *1 240.16,287
X$35704 503 489 505 2 3 532 AND3_X1
* cell instance $35708 m0 *1 241.87,287
X$35708 506 504 501 2 3 531 AND3_X1
* cell instance $35709 r0 *1 242.82,284.2
X$35709 505 504 506 3 2 465 NAND3_X2
* cell instance $35713 m0 *1 242.82,287
X$35713 463 3 2 842 INV_X4
* cell instance $35717 m0 *1 246.24,287
X$35717 513 3 2 537 INV_X1
* cell instance $35720 r0 *1 247.57,284.2
X$35720 501 513 503 3 2 520 NAND3_X2
* cell instance $35722 m0 *1 248.33,287
X$35722 523 3 2 843 INV_X4
* cell instance $35724 r0 *1 249.47,284.2
X$35724 3 217 520 469 467 2 AOI21_X4
* cell instance $35727 r0 *1 253.46,284.2
X$35727 519 522 521 2 3 130 OAI21_X4
* cell instance $35731 r0 *1 258.4,284.2
X$35731 3 778 514 517 511 2 DFF_X1
* cell instance $35737 m0 *1 253.46,287
X$35737 533 522 521 2 3 202 OAI21_X4
* cell instance $35741 m0 *1 255.93,287
X$35741 3 707 530 524 523 2 DFF_X1
* cell instance $35745 r0 *1 265.81,284.2
X$35745 528 466 521 2 3 444 OAI21_X4
* cell instance $35790 m0 *1 266.95,287
X$35790 521 526 516 3 2 NOR2_X4
* cell instance $35793 m0 *1 270.56,287
X$35793 105 3 2 507 CLKBUF_X3
* cell instance $35794 m0 *1 271.51,287
X$35794 507 3 2 844 INV_X4
* cell instance $35851 r0 *1 514.33,284.2
X$35851 516 3 2 508 BUF_X1
* cell instance $35928 r0 *1 217.93,259
X$35928 3 804 310 309 236 2 DFF_X1
* cell instance $35956 r0 *1 225.34,259
X$35956 3 784 295 294 236 2 DFF_X1
* cell instance $35961 r0 *1 235.03,259
X$35961 299 115 300 3 2 313 MUX2_X1
* cell instance $35964 r0 *1 236.74,259
X$35964 3 818 300 313 212 2 DFF_X1
* cell instance $35967 m0 *1 237.5,261.8
X$35967 299 125 334 3 2 352 MUX2_X1
* cell instance $35969 m0 *1 239.59,261.8
X$35969 299 3 2 316 BUF_X2
* cell instance $35972 r0 *1 240.35,259
X$35972 300 155 301 3 2 315 MUX2_X1
* cell instance $35975 r0 *1 246.43,259
X$35975 3 761 325 302 172 2 DFF_X1
* cell instance $35981 r0 *1 265.81,259
X$35981 3 783 304 303 314 2 DFF_X1
* cell instance $35984 r0 *1 269.99,259
X$35984 305 171 307 3 2 323 MUX2_X1
* cell instance $35986 r0 *1 274.36,259
X$35986 306 217 316 3 2 311 MUX2_X1
* cell instance $35987 r0 *1 275.69,259
X$35987 322 203 306 3 2 307 MUX2_X1
* cell instance $36007 m0 *1 242.25,261.8
X$36007 337 171 315 3 2 328 MUX2_X1
* cell instance $36011 m0 *1 245.67,261.8
X$36011 325 30 316 3 2 302 MUX2_X1
* cell instance $36014 m0 *1 248.14,261.8
X$36014 317 15 316 3 2 338 MUX2_X1
* cell instance $36016 m0 *1 250.23,261.8
X$36016 325 27 317 3 2 331 MUX2_X1
* cell instance $36017 m0 *1 251.56,261.8
X$36017 3 702 318 329 330 2 DFF_X1
* cell instance $36018 m0 *1 254.79,261.8
X$36018 318 39 316 3 2 329 MUX2_X1
* cell instance $36024 m0 *1 256.69,261.8
X$36024 339 46 331 3 2 319 MUX2_X1
* cell instance $36025 m0 *1 258.02,261.8
X$36025 87 319 84 296 2 3 327 OAI22_X1
* cell instance $36027 m0 *1 259.35,261.8
X$36027 195 328 196 323 2 3 326 OAI22_X1
* cell instance $36028 m0 *1 260.3,261.8
X$36028 327 326 3 2 347 OR2_X1
* cell instance $36031 m0 *1 267.9,261.8
X$36031 316 130 304 3 2 303 MUX2_X1
* cell instance $36032 m0 *1 269.23,261.8
X$36032 304 158 324 3 2 305 MUX2_X1
* cell instance $36033 m0 *1 270.56,261.8
X$36033 324 132 316 3 2 346 MUX2_X1
* cell instance $36035 m0 *1 274.93,261.8
X$36035 316 202 322 3 2 321 MUX2_X1
* cell instance $36038 m0 *1 277.4,261.8
X$36038 3 705 322 321 320 2 DFF_X1
* cell instance $36219 r0 *1 223.25,264.6
X$36219 362 110 356 3 2 355 MUX2_X1
* cell instance $36220 r0 *1 221.92,264.6
X$36220 362 108 354 3 2 361 MUX2_X1
* cell instance $36223 r0 *1 225.53,264.6
X$36223 354 96 356 3 2 364 MUX2_X1
* cell instance $36228 r0 *1 232.37,264.6
X$36228 340 2 96 3 BUF_X4
* cell instance $36236 m0 *1 223.06,267.4
X$36236 3 737 356 355 236 2 DFF_X1
* cell instance $36241 m0 *1 234.46,267.4
X$36241 362 3 2 344 BUF_X2
* cell instance $36251 r0 *1 248.52,264.6
X$36251 360 3 2 105 CLKBUF_X3
* cell instance $36261 r0 *1 260.49,264.6
X$36261 333 2 203 3 BUF_X4
* cell instance $36267 m0 *1 269.61,267.4
X$36267 3 696 363 358 320 2 DFF_X1
* cell instance $36269 r0 *1 269.8,264.6
X$36269 363 132 344 3 2 358 MUX2_X1
* cell instance $36317 m0 *1 273.98,267.4
X$36317 344 202 370 3 2 373 MUX2_X1
* cell instance $36318 m0 *1 275.31,267.4
X$36318 371 217 344 3 2 359 MUX2_X1
* cell instance $36319 m0 *1 276.64,267.4
X$36319 3 692 371 359 320 2 DFF_X1
* cell instance $36461 m0 *1 221.54,270.2
X$36461 3 727 376 408 389 2 DFF_X1
* cell instance $36462 m0 *1 224.77,270.2
X$36462 376 23 400 3 2 377 MUX2_X1
* cell instance $36463 m0 *1 226.1,270.2
X$36463 377 62 364 3 2 391 MUX2_X1
* cell instance $36467 m0 *1 229.9,270.2
X$36467 362 125 378 3 2 410 MUX2_X1
* cell instance $36472 r0 *1 233.32,267.4
X$36472 340 2 23 3 BUF_X4
* cell instance $36473 r0 *1 237.69,267.4
X$36473 333 2 158 3 BUF_X4
* cell instance $36476 r0 *1 240.73,267.4
X$36476 366 2 62 3 BUF_X4
* cell instance $36479 m0 *1 233.32,270.2
X$36479 378 333 379 3 2 394 MUX2_X1
* cell instance $36482 m0 *1 235.22,270.2
X$36482 394 171 393 3 2 390 MUX2_X1
* cell instance $36487 m0 *1 241.68,270.2
X$36487 395 30 381 3 2 402 MUX2_X1
* cell instance $36489 m0 *1 243.77,270.2
X$36489 395 23 403 3 2 397 MUX2_X1
* cell instance $36491 r0 *1 245.67,267.4
X$36491 3 799 382 380 330 2 DFF_X1
* cell instance $36496 m0 *1 245.86,270.2
X$36496 382 39 381 3 2 380 MUX2_X1
* cell instance $36498 m0 *1 247.95,270.2
X$36498 382 23 383 3 2 396 MUX2_X1
* cell instance $36500 m0 *1 250.04,270.2
X$36500 396 62 397 3 2 384 MUX2_X1
* cell instance $36503 m0 *1 252.51,270.2
X$36503 398 39 344 3 2 365 MUX2_X1
* cell instance $36504 r0 *1 253.27,267.4
X$36504 3 797 398 365 330 2 DFF_X1
* cell instance $36508 m0 *1 255.36,270.2
X$36508 399 26 344 3 2 412 MUX2_X1
* cell instance $36510 r0 *1 256.88,267.4
X$36510 366 2 46 3 BUF_X4
* cell instance $36511 r0 *1 258.21,267.4
X$36511 375 96 3 196 2 NAND2_X4
* cell instance $36512 r0 *1 259.92,267.4
X$36512 203 375 3 2 367 OR2_X1
* cell instance $36513 r0 *1 260.68,267.4
X$36513 96 385 3 2 374 OR2_X1
* cell instance $36514 r0 *1 261.44,267.4
X$36514 374 3 2 195 BUF_X2
* cell instance $36518 m0 *1 256.88,270.2
X$36518 398 340 399 3 2 392 MUX2_X1
* cell instance $36520 m0 *1 258.59,270.2
X$36520 375 3 2 385 INV_X1
* cell instance $36521 m0 *1 258.97,270.2
X$36521 385 203 3 84 2 NAND2_X4
* cell instance $36522 m0 *1 260.68,270.2
X$36522 367 3 2 87 CLKBUF_X3
* cell instance $36523 m0 *1 261.63,270.2
X$36523 392 46 357 3 2 386 MUX2_X1
* cell instance $36525 m0 *1 263.34,270.2
X$36525 195 390 196 388 2 3 406 OAI22_X1
* cell instance $36528 m0 *1 265.43,270.2
X$36528 3 698 368 387 314 2 DFF_X1
* cell instance $36530 r0 *1 266.38,267.4
X$36530 344 130 368 3 2 387 MUX2_X1
* cell instance $36531 r0 *1 269.23,267.4
X$36531 368 158 363 3 2 369 MUX2_X1
* cell instance $36532 r0 *1 270.56,267.4
X$36532 369 171 372 3 2 388 MUX2_X1
* cell instance $36536 r0 *1 273.22,267.4
X$36536 3 806 370 373 320 2 DFF_X1
* cell instance $36538 r0 *1 276.45,267.4
X$36538 370 203 371 3 2 372 MUX2_X1
* cell instance $36751 r0 *1 221.16,270.2
X$36751 362 52 376 3 2 408 MUX2_X1
* cell instance $36753 r0 *1 224.77,270.2
X$36753 362 57 400 3 2 409 MUX2_X1
* cell instance $36757 m0 *1 223.63,273
X$36757 3 689 400 409 389 2 DFF_X1
* cell instance $36759 r0 *1 228.19,270.2
X$36759 3 814 378 410 389 2 DFF_X1
* cell instance $36761 r0 *1 231.42,270.2
X$36761 3 812 379 411 389 2 DFF_X1
* cell instance $36762 r0 *1 234.65,270.2
X$36762 379 213 344 3 2 411 MUX2_X1
* cell instance $36768 m0 *1 237.12,273
X$36768 435 171 401 3 2 404 MUX2_X1
* cell instance $36770 r0 *1 239.59,270.2
X$36770 366 2 171 3 BUF_X4
* cell instance $36772 r0 *1 240.92,270.2
X$36772 3 795 395 402 330 2 DFF_X1
* cell instance $36774 r0 *1 244.91,270.2
X$36774 3 819 383 414 330 2 DFF_X1
* cell instance $36775 r0 *1 248.14,270.2
X$36775 383 26 381 3 2 414 MUX2_X1
* cell instance $36781 m0 *1 241.3,273
X$36781 3 714 403 413 330 2 DFF_X1
* cell instance $36782 m0 *1 244.53,273
X$36782 403 15 381 3 2 413 MUX2_X1
* cell instance $36784 r0 *1 250.8,270.2
X$36784 415 84 384 87 2 3 436 OAI22_X1
* cell instance $36791 r0 *1 254.41,270.2
X$36791 3 796 399 412 330 2 DFF_X1
* cell instance $36794 r0 *1 262.39,270.2
X$36794 87 386 84 391 2 3 405 OAI22_X1
* cell instance $36795 r0 *1 263.34,270.2
X$36795 405 406 3 2 460 OR2_X1
* cell instance $36820 m0 *1 258.59,273
X$36820 418 196 404 195 2 3 419 OAI22_X1
* cell instance $36821 m0 *1 259.54,273
X$36821 436 419 3 2 407 OR2_X1
* cell instance $37013 r0 *1 244.15,306.6
X$37013 654 648 647 2 3 660 HA_X1
* cell instance $37016 r0 *1 246.24,306.6
X$37016 646 574 655 2 3 662 HA_X1
* cell instance $37017 r0 *1 248.14,306.6
X$37017 3 656 662 642 650 651 636 2 AOI221_X4
* cell instance $37021 r0 *1 258.97,306.6
X$37021 3 645 652 517 511 2 DFF_X1
* cell instance $37022 r0 *1 262.2,306.6
X$37022 3 654 653 551 511 2 DFF_X1
* cell instance $37042 m0 *1 244.53,309.4
X$37042 647 3 2 658 BUF_X2
* cell instance $37045 m0 *1 246.43,309.4
X$37045 658 642 2 3 664 AND2_X1
* cell instance $37046 m0 *1 247.19,309.4
X$37046 650 658 660 649 664 575 2 3 AOI221_X2
* cell instance $37211 r0 *1 229.9,261.8
X$37211 3 817 332 348 212 2 DFF_X1
* cell instance $37213 r0 *1 233.32,261.8
X$37213 3 816 350 351 212 2 DFF_X1
* cell instance $37238 m0 *1 220.97,264.6
X$37238 3 728 354 361 236 2 DFF_X1
* cell instance $37242 m0 *1 230.85,264.6
X$37242 362 115 332 3 2 348 MUX2_X1
* cell instance $37244 m0 *1 232.37,264.6
X$37244 332 155 350 3 2 393 MUX2_X1
* cell instance $37246 m0 *1 234.08,264.6
X$37246 350 187 344 3 2 351 MUX2_X1
* cell instance $37249 m0 *1 236.36,264.6
X$37249 333 2 155 3 BUF_X4
* cell instance $37251 r0 *1 236.93,261.8
X$37251 3 808 334 352 212 2 DFF_X1
* cell instance $37252 r0 *1 240.35,261.8
X$37252 336 213 316 3 2 335 MUX2_X1
* cell instance $37253 r0 *1 241.68,261.8
X$37253 334 333 336 3 2 337 MUX2_X1
* cell instance $37260 m0 *1 241.3,264.6
X$37260 3 736 336 335 212 2 DFF_X1
* cell instance $37262 r0 *1 248.14,261.8
X$37262 3 798 317 338 172 2 DFF_X1
* cell instance $37266 r0 *1 253.65,261.8
X$37266 3 768 341 353 330 2 DFF_X1
* cell instance $37267 r0 *1 256.88,261.8
X$37267 341 26 316 3 2 353 MUX2_X1
* cell instance $37268 r0 *1 258.21,261.8
X$37268 3 776 342 349 314 2 DFF_X1
* cell instance $37269 r0 *1 261.44,261.8
X$37269 342 30 344 3 2 349 MUX2_X1
* cell instance $37276 m0 *1 254.98,264.6
X$37276 318 340 341 3 2 339 MUX2_X1
* cell instance $37280 m0 *1 256.31,264.6
X$37280 340 2 27 3 BUF_X4
* cell instance $37283 m0 *1 261.06,264.6
X$37283 342 27 343 3 2 357 MUX2_X1
* cell instance $37287 r0 *1 264.67,261.8
X$37287 343 15 344 3 2 345 MUX2_X1
* cell instance $37290 r0 *1 269.99,261.8
X$37290 3 767 324 346 320 2 DFF_X1
* cell instance $37309 m0 *1 264.86,264.6
X$37309 3 697 343 345 314 2 DFF_X1
* cell instance $37492 m0 *1 243.2,317.8
X$37492 667 641 2 675 3 XOR2_X2
* cell instance $37493 r0 *1 244.91,315
X$37493 641 3 2 665 INV_X2
* cell instance $37495 r0 *1 245.48,315
X$37495 658 665 667 666 3 2 657 OR4_X1
* cell instance $37496 r0 *1 246.62,315
X$37496 666 667 665 658 3 2 663 NOR4_X1
* cell instance $37548 m0 *1 245.67,317.8
X$37548 666 667 3 2 671 NAND2_X1
* cell instance $37551 m0 *1 248.14,317.8
X$37551 672 3 2 667 CLKBUF_X2
* cell instance $37720 r0 *1 242.63,301
X$37720 625 630 629 3 2 640 MUX2_X1
* cell instance $37722 r0 *1 243.96,301
X$37722 626 466 580 3 630 2 AOI21_X1
* cell instance $37726 r0 *1 247.19,301
X$37726 612 573 641 2 3 635 HA_X1
* cell instance $37731 r0 *1 260.49,301
X$37731 633 526 580 3 627 2 AOI21_X1
* cell instance $37736 m0 *1 249.09,303.8
X$37736 635 3 2 636 INV_X1
* cell instance $37742 r0 *1 262.58,301
X$37742 581 578 605 576 3 2 638 NAND4_X1
* cell instance $37790 m0 *1 262.77,303.8
X$37790 638 526 580 3 637 2 AOI21_X1
* cell instance $37926 r0 *1 239.97,292.6
X$37926 572 571 823 2 3 489 HA_X1
* cell instance $37928 r0 *1 243.39,292.6
X$37928 535 467 466 3 583 2 AOI21_X2
* cell instance $37931 r0 *1 249.28,292.6
X$37931 563 575 2 550 3 XOR2_X2
* cell instance $37934 r0 *1 255.55,292.6
X$37934 585 561 584 3 2 560 MUX2_X1
* cell instance $37935 r0 *1 256.88,292.6
X$37935 543 578 2 3 585 AND2_X1
* cell instance $37936 r0 *1 257.64,292.6
X$37936 454 579 2 3 584 AND2_X1
* cell instance $37938 r0 *1 259.92,292.6
X$37938 581 3 2 597 INV_X1
* cell instance $37942 r0 *1 265.05,292.6
X$37942 564 592 3 2 563 XNOR2_X2
* cell instance $37965 m0 *1 237.31,295.4
X$37965 3 596 463 571 574 2 DFF_X2
* cell instance $37968 m0 *1 241.3,295.4
X$37968 573 571 595 2 3 504 HA_X1
* cell instance $37970 m0 *1 243.39,295.4
X$37970 572 574 822 2 3 513 HA_X1
* cell instance $37972 m0 *1 246.05,295.4
X$37972 573 574 821 2 3 512 HA_X1
* cell instance $37976 m0 *1 255.93,295.4
X$37976 543 576 2 3 586 AND2_X1
* cell instance $37977 m0 *1 256.69,295.4
X$37977 576 540 3 2 562 NOR2_X1
* cell instance $37980 m0 *1 258.21,295.4
X$37980 578 577 579 3 2 599 MUX2_X1
* cell instance $37981 m0 *1 259.54,295.4
X$37981 597 526 580 3 577 2 AOI21_X1
* cell instance $37982 m0 *1 260.3,295.4
X$37982 3 599 511 825 578 2 DFF_X2
* cell instance $37985 r0 *1 267.33,292.6
X$37985 580 526 3 2 447 NAND2_X2
* cell instance $38192 r0 *1 237.31,298.2
X$38192 3 617 463 573 572 2 DFF_X2
* cell instance $38195 r0 *1 241.68,298.2
X$38195 620 583 600 3 2 617 MUX2_X1
* cell instance $38199 r0 *1 247,298.2
X$38199 506 540 3 2 610 NOR2_X1
* cell instance $38200 r0 *1 247.57,298.2
X$38200 610 622 601 3 2 631 MUX2_X1
* cell instance $38201 r0 *1 248.9,298.2
X$38201 611 2 503 3 BUF_X4
* cell instance $38202 r0 *1 250.23,298.2
X$38202 611 3 2 506 INV_X4
* cell instance $38211 m0 *1 241.87,301
X$38211 543 536 2 3 625 AND2_X1
* cell instance $38214 m0 *1 244.34,301
X$38214 572 574 503 549 3 2 626 NAND4_X1
* cell instance $38217 m0 *1 245.86,301
X$38217 536 540 3 2 629 NOR2_X1
* cell instance $38218 m0 *1 246.43,301
X$38218 3 631 523 829 611 2 DFF_X2
* cell instance $38222 m0 *1 251.37,301
X$38222 643 3 2 549 BUF_X2
* cell instance $38224 r0 *1 258.21,298.2
X$38224 612 3 2 576 BUF_X1
* cell instance $38225 r0 *1 254.6,298.2
X$38225 3 609 523 831 612 2 DFF_X2
* cell instance $38229 r0 *1 261.06,298.2
X$38229 543 605 2 3 634 AND2_X1
* cell instance $38230 r0 *1 259.16,298.2
X$38230 612 578 579 2 3 613 HA_X1
* cell instance $38231 r0 *1 261.82,298.2
X$38231 605 540 3 2 632 NOR2_X1
* cell instance $38232 r0 *1 262.39,298.2
X$38232 614 526 580 3 624 2 AOI21_X1
* cell instance $38233 r0 *1 263.15,298.2
X$38233 613 565 3 2 614 NAND2_X1
* cell instance $38234 r0 *1 263.72,298.2
X$38234 543 623 2 3 615 AND2_X1
* cell instance $38238 m0 *1 260.87,301
X$38238 581 613 3 2 633 NAND2_X1
* cell instance $38239 m0 *1 261.44,301
X$38239 634 624 632 3 2 517 MUX2_X1
* cell instance $38240 m0 *1 262.77,301
X$38240 615 604 628 3 2 551 MUX2_X1
* cell instance $38241 m0 *1 264.1,301
X$38241 623 540 3 2 628 NOR2_X1
* cell instance $38243 r0 *1 265.05,298.2
X$38243 623 605 613 565 3 2 616 NAND4_X1
* cell instance $38246 r0 *1 266.76,298.2
X$38246 621 526 580 3 619 2 AOI21_X1
* cell instance $38248 r0 *1 269.04,298.2
X$38248 592 619 3 2 618 XOR2_X1
* cell instance $38250 m0 *1 265.05,301
X$38250 581 623 605 613 3 2 621 NAND4_X1
* cell instance $38252 r0 *1 273.79,298.2
X$38252 606 3 2 592 CLKBUF_X2
* cell instance $38253 r0 *1 270.56,298.2
X$38253 3 807 606 618 507 2 DFF_X1
* cell instance $38440 r0 *1 240.73,295.4
X$38440 543 574 2 3 587 AND2_X1
* cell instance $38441 r0 *1 241.49,295.4
X$38441 587 583 598 3 2 596 MUX2_X1
* cell instance $38442 r0 *1 242.82,295.4
X$38442 454 595 2 3 598 AND2_X1
* cell instance $38475 m0 *1 241.3,298.2
X$38475 543 572 2 3 620 AND2_X1
* cell instance $38476 m0 *1 242.06,298.2
X$38476 454 573 2 3 600 AND2_X1
* cell instance $38563 m0 *1 229.52,284.2
X$38563 3 732 497 509 463 2 DFF_X1
* cell instance $38565 r0 *1 231.04,281.4
X$38565 438 57 497 3 2 509 MUX2_X1
* cell instance $38567 r0 *1 233.32,281.4
X$38567 462 340 497 3 2 498 MUX2_X1
* cell instance $38569 r0 *1 235.41,281.4
X$38569 498 366 529 3 2 415 MUX2_X1
* cell instance $38576 m0 *1 240.16,284.2
X$38576 503 504 505 2 3 518 AND3_X1
* cell instance $38581 m0 *1 242.63,284.2
X$38581 501 504 503 3 2 464 NAND3_X2
* cell instance $38583 r0 *1 243.2,281.4
X$38583 501 489 503 3 2 488 NAND3_X2
* cell instance $38586 m0 *1 243.96,284.2
X$38586 505 513 506 3 2 479 NAND3_X2
* cell instance $38587 m0 *1 245.29,284.2
X$38587 505 489 506 3 2 468 NAND3_X2
* cell instance $38588 m0 *1 246.62,284.2
X$38588 505 512 506 3 2 500 NAND3_X2
* cell instance $38590 r0 *1 247.19,281.4
X$38590 501 512 503 3 2 482 NAND3_X2
* cell instance $38600 m0 *1 250.8,284.2
X$38600 3 466 2 469 BUF_X8
* cell instance $38605 m0 *1 257.64,284.2
X$38605 530 3 2 366 CLKBUF_X3
* cell instance $38608 m0 *1 260.87,284.2
X$38608 514 3 2 333 CLKBUF_X3
* cell instance $38609 m0 *1 261.82,284.2
X$38609 3 551 511 826 375 2 DFF_X2
* cell instance $38611 r0 *1 266.57,281.4
X$38611 3 471 507 834 472 2 DFF_X2
* cell instance $38616 m0 *1 268.09,284.2
X$38616 3 510 507 827 491 2 DFF_X2
* cell instance $38617 r0 *1 270.75,281.4
X$38617 444 201 490 502 447 2 3 510 OAI221_X1
* cell instance $38619 r0 *1 271.89,281.4
X$38619 491 454 3 2 502 NAND2_X1
* cell instance $38620 r0 *1 272.46,281.4
X$38620 445 491 446 3 2 490 NAND3_X1
* cell instance $38623 m0 *1 273.22,284.2
X$38623 445 493 446 3 2 492 NAND3_X1
* cell instance $38625 r0 *1 273.6,281.4
X$38625 493 454 3 2 499 NAND2_X1
* cell instance $38626 r0 *1 274.36,281.4
X$38626 3 484 507 830 493 2 DFF_X2
* cell instance $38670 r0 *1 508.82,281.4
X$38670 472 3 2 495 BUF_X1
* cell instance $38672 r0 *1 510.15,281.4
X$38672 491 3 2 496 BUF_X1
* cell instance $38715 r0 *1 511.29,281.4
X$38715 493 3 2 494 BUF_X1
* cell instance $38851 m0 *1 228.38,275.8
X$38851 3 703 437 448 389 2 DFF_X1
* cell instance $38853 m0 *1 232.37,275.8
X$38853 3 704 439 449 389 2 DFF_X1
* cell instance $38854 r0 *1 233.51,273
X$38854 434 3 2 362 BUF_X1
* cell instance $38863 r0 *1 266.19,273
X$38863 105 3 2 314 CLKBUF_X3
* cell instance $38864 r0 *1 267.14,273
X$38864 314 3 2 845 INV_X4
* cell instance $38865 r0 *1 268.09,273
X$38865 444 433 432 431 447 2 3 461 OAI221_X1
* cell instance $38867 r0 *1 269.99,273
X$38867 445 430 446 3 2 432 NAND3_X1
* cell instance $38869 r0 *1 270.94,273
X$38869 3 429 320 832 422 2 DFF_X2
* cell instance $38886 m0 *1 235.6,275.8
X$38886 437 158 450 3 2 435 MUX2_X1
* cell instance $38887 m0 *1 236.93,275.8
X$38887 439 158 416 3 2 401 MUX2_X1
* cell instance $38898 m0 *1 247.19,275.8
X$38898 3 26 500 469 467 2 AOI21_X4
* cell instance $38901 m0 *1 254.22,275.8
X$38901 381 130 417 3 2 455 MUX2_X1
* cell instance $38906 m0 *1 255.93,275.8
X$38906 417 333 470 3 2 457 MUX2_X1
* cell instance $38909 m0 *1 257.83,275.8
X$38909 457 366 459 3 2 418 MUX2_X1
* cell instance $38911 m0 *1 259.35,275.8
X$38911 458 333 440 3 2 459 MUX2_X1
* cell instance $38914 m0 *1 261.25,275.8
X$38914 381 202 458 3 2 441 MUX2_X1
* cell instance $38918 m0 *1 266.19,275.8
X$38918 442 454 3 2 420 NAND2_X1
* cell instance $38919 m0 *1 266.76,275.8
X$38919 444 460 443 420 447 2 3 421 OAI221_X1
* cell instance $38920 m0 *1 267.9,275.8
X$38920 3 461 320 828 430 2 DFF_X2
* cell instance $38921 m0 *1 271.51,275.8
X$38921 444 347 456 453 447 2 3 429 OAI221_X1
* cell instance $38922 m0 *1 272.65,275.8
X$38922 105 3 2 320 CLKBUF_X3
* cell instance $38923 m0 *1 273.6,275.8
X$38923 320 3 2 839 INV_X2
* cell instance $38924 m0 *1 274.17,275.8
X$38924 444 273 428 452 447 2 3 427 OAI221_X1
* cell instance $38925 m0 *1 275.31,275.8
X$38925 423 446 3 2 452 NAND2_X1
* cell instance $38926 m0 *1 275.88,275.8
X$38926 445 423 446 3 2 428 NAND3_X1
* cell instance $38930 m0 *1 279.11,275.8
X$38930 3 427 320 824 423 2 DFF_X2
* cell instance $39014 m0 *1 509.39,275.8
X$39014 430 3 2 424 BUF_X1
* cell instance $39018 m0 *1 512.43,275.8
X$39018 423 3 2 426 BUF_X1
* cell instance $39021 m0 *1 514.9,275.8
X$39021 422 3 2 425 BUF_X1
* cell instance $39160 m0 *1 214.32,245
X$39160 3 718 193 204 236 2 DFF_X1
* cell instance $39161 r0 *1 216.41,242.2
X$39161 3 762 166 180 50 2 DFF_X1
* cell instance $39162 r0 *1 215.08,242.2
X$39162 153 108 166 3 2 180 MUX2_X1
* cell instance $39165 r0 *1 221.92,242.2
X$39165 153 52 167 3 2 183 MUX2_X1
* cell instance $39168 r0 *1 224.2,242.2
X$39168 153 57 168 3 2 185 MUX2_X1
* cell instance $39169 r0 *1 225.53,242.2
X$39169 3 793 168 185 50 2 DFF_X1
* cell instance $39173 r0 *1 232.75,242.2
X$39173 139 155 169 3 2 189 MUX2_X1
* cell instance $39176 r0 *1 235.79,242.2
X$39176 189 171 190 3 2 161 MUX2_X1
* cell instance $39177 r0 *1 237.12,242.2
X$39177 3 773 156 191 9 2 DFF_X1
* cell instance $39178 r0 *1 240.35,242.2
X$39178 156 213 7 3 2 191 MUX2_X1
* cell instance $39181 m0 *1 217.55,245
X$39181 153 110 193 3 2 204 MUX2_X1
* cell instance $39182 m0 *1 218.88,245
X$39182 166 96 193 3 2 206 MUX2_X1
* cell instance $39186 m0 *1 221.54,245
X$39186 3 713 167 183 236 2 DFF_X1
* cell instance $39187 m0 *1 224.77,245
X$39187 167 96 168 3 2 194 MUX2_X1
* cell instance $39188 m0 *1 226.1,245
X$39188 194 62 206 3 2 188 MUX2_X1
* cell instance $39192 m0 *1 229.9,245
X$39192 3 690 169 207 236 2 DFF_X1
* cell instance $39193 m0 *1 233.13,245
X$39193 169 213 22 3 2 207 MUX2_X1
* cell instance $39198 m0 *1 241.3,245
X$39198 170 187 7 3 2 208 MUX2_X1
* cell instance $39201 r0 *1 242.82,242.2
X$39201 164 171 163 3 2 184 MUX2_X1
* cell instance $39207 m0 *1 247,245
X$39207 3 688 230 209 172 2 DFF_X1
* cell instance $39210 m0 *1 250.8,245
X$39210 87 138 84 188 2 3 233 OAI22_X1
* cell instance $39212 m0 *1 254.79,245
X$39212 172 3 2 838 INV_X2
* cell instance $39213 m0 *1 255.36,245
X$39213 105 3 2 172 CLKBUF_X3
* cell instance $39325 m0 *1 221.35,228.2
X$39325 3 744 59 72 50 2 DFF_X1
* cell instance $39327 r0 *1 227.43,225.4
X$39327 51 57 56 3 2 34 MUX2_X1
* cell instance $39329 r0 *1 228.76,225.4
X$39329 3 750 53 35 50 2 DFF_X1
* cell instance $39338 m0 *1 228.19,228.2
X$39338 51 52 53 3 2 35 MUX2_X1
* cell instance $39340 m0 *1 229.9,228.2
X$39340 53 23 56 3 2 89 MUX2_X1
* cell instance $39343 m0 *1 240.35,228.2
X$39343 51 3 2 7 BUF_X2
* cell instance $39352 m0 *1 255.36,228.2
X$39352 54 39 38 3 2 71 MUX2_X1
* cell instance $39353 m0 *1 256.69,228.2
X$39353 3 747 54 71 11 2 DFF_X1
* cell instance $39355 r0 *1 259.73,225.4
X$39355 54 27 41 3 2 70 MUX2_X1
* cell instance $39357 r0 *1 262.77,225.4
X$39357 42 30 38 3 2 69 MUX2_X1
* cell instance $39360 m0 *1 260.68,228.2
X$39360 70 46 55 3 2 68 MUX2_X1
* cell instance $39363 m0 *1 263.15,228.2
X$39363 3 735 42 69 11 2 DFF_X1
* cell instance $39365 r0 *1 264.48,225.4
X$39365 42 27 43 3 2 55 MUX2_X1
* cell instance $39490 r0 *1 217.93,233.8
X$39490 60 108 113 3 2 111 MUX2_X1
* cell instance $39493 r0 *1 220.21,233.8
X$39493 60 110 114 3 2 112 MUX2_X1
* cell instance $39496 r0 *1 222.49,233.8
X$39496 113 96 114 3 2 64 MUX2_X1
* cell instance $39498 r0 *1 224.58,233.8
X$39498 51 108 98 3 2 122 MUX2_X1
* cell instance $39499 r0 *1 225.91,233.8
X$39499 3 753 98 122 50 2 DFF_X1
* cell instance $39505 r0 *1 256.5,233.8
X$39505 3 780 118 116 11 2 DFF_X1
* cell instance $39506 r0 *1 259.73,233.8
X$39506 118 27 119 3 2 123 MUX2_X1
* cell instance $39507 r0 *1 261.06,233.8
X$39507 123 46 120 3 2 176 MUX2_X1
* cell instance $39601 m0 *1 219.83,236.6
X$39601 3 745 114 112 50 2 DFF_X1
* cell instance $39605 m0 *1 232.37,236.6
X$39605 60 115 124 3 2 135 MUX2_X1
* cell instance $39608 m0 *1 237.12,236.6
X$39608 51 125 127 3 2 126 MUX2_X1
* cell instance $39612 m0 *1 239.78,236.6
X$39612 51 115 129 3 2 128 MUX2_X1
* cell instance $39781 r0 *1 234.46,222.6
X$39781 3 791 37 31 9 2 DFF_X1
* cell instance $39784 r0 *1 238.64,222.6
X$39784 3 771 21 18 9 2 DFF_X1
* cell instance $39785 r0 *1 241.87,222.6
X$39785 21 30 22 3 2 18 MUX2_X1
* cell instance $39786 r0 *1 243.2,222.6
X$39786 10 15 22 3 2 19 MUX2_X1
* cell instance $39789 r0 *1 246.24,222.6
X$39789 3 749 48 24 4 2 DFF_X1
* cell instance $39790 r0 *1 249.47,222.6
X$39790 33 26 22 3 2 17 MUX2_X1
* cell instance $39820 m0 *1 227.62,225.4
X$39820 3 716 56 34 50 2 DFF_X1
* cell instance $39823 m0 *1 234.08,225.4
X$39823 8 52 36 3 2 20 MUX2_X1
* cell instance $39824 m0 *1 235.41,225.4
X$39824 8 57 37 3 2 31 MUX2_X1
* cell instance $39826 m0 *1 236.93,225.4
X$39826 36 23 37 3 2 66 MUX2_X1
* cell instance $39834 m0 *1 243.2,225.4
X$39834 21 23 10 3 2 47 MUX2_X1
* cell instance $39837 m0 *1 246.24,225.4
X$39837 48 39 22 3 2 24 MUX2_X1
* cell instance $39839 m0 *1 248.33,225.4
X$39839 8 3 2 38 BUF_X2
* cell instance $39840 m0 *1 249.09,225.4
X$39840 48 27 33 3 2 25 MUX2_X1
* cell instance $39844 r0 *1 253.46,222.6
X$39844 28 39 7 3 2 40 MUX2_X1
* cell instance $39847 r0 *1 257.26,222.6
X$39847 28 27 5 3 2 32 MUX2_X1
* cell instance $39848 r0 *1 258.59,222.6
X$39848 3 772 41 29 11 2 DFF_X1
* cell instance $39849 r0 *1 261.82,222.6
X$39849 12 30 7 3 2 6 MUX2_X1
* cell instance $39850 r0 *1 263.15,222.6
X$39850 12 27 13 3 2 45 MUX2_X1
* cell instance $39852 r0 *1 265.24,222.6
X$39852 3 763 13 14 11 2 DFF_X1
* cell instance $39870 m0 *1 254.22,225.4
X$39870 3 738 28 40 11 2 DFF_X1
* cell instance $39874 m0 *1 257.45,225.4
X$39874 41 26 38 3 2 29 MUX2_X1
* cell instance $39877 m0 *1 259.92,225.4
X$39877 32 46 45 3 2 90 MUX2_X1
* cell instance $39882 m0 *1 268.66,225.4
X$39882 43 15 38 3 2 44 MUX2_X1
* cell instance $39883 m0 *1 269.99,225.4
X$39883 3 733 43 44 11 2 DFF_X1
* cell instance $40037 r0 *1 209.38,245
X$40037 192 3 2 210 BUF_X1
* cell instance $40071 m0 *1 235.41,247.8
X$40071 227 187 117 3 2 226 MUX2_X1
* cell instance $40075 r0 *1 239.97,245
X$40075 3 785 170 208 212 2 DFF_X1
* cell instance $40082 r0 *1 248.71,245
X$40082 231 187 38 3 2 229 MUX2_X1
* cell instance $40083 r0 *1 247.38,245
X$40083 230 213 38 3 2 209 MUX2_X1
* cell instance $40088 m0 *1 247.57,247.8
X$40088 3 687 231 229 172 2 DFF_X1
* cell instance $40092 m0 *1 253.46,247.8
X$40092 216 217 22 3 2 214 MUX2_X1
* cell instance $40094 r0 *1 254.22,245
X$40094 3 754 216 214 172 2 DFF_X1
* cell instance $40097 r0 *1 262.77,245
X$40097 7 202 198 3 2 228 MUX2_X1
* cell instance $40099 m0 *1 254.79,247.8
X$40099 22 202 215 3 2 234 MUX2_X1
* cell instance $40103 m0 *1 256.12,247.8
X$40103 215 203 216 3 2 174 MUX2_X1
* cell instance $40106 m0 *1 262.01,247.8
X$40106 3 719 198 228 143 2 DFF_X1
* cell instance $40108 r0 *1 264.48,245
X$40108 198 203 200 3 2 199 MUX2_X1
* cell instance $40110 r0 *1 270.37,245
X$40110 221 217 38 3 2 223 MUX2_X1
* cell instance $40111 r0 *1 271.7,245
X$40111 3 801 221 223 143 2 DFF_X1
* cell instance $40157 m0 *1 265.24,247.8
X$40157 200 217 7 3 2 218 MUX2_X1
* cell instance $40161 m0 *1 268.66,247.8
X$40161 3 723 219 222 143 2 DFF_X1
* cell instance $40162 m0 *1 271.89,247.8
X$40162 38 202 219 3 2 222 MUX2_X1
* cell instance $40163 m0 *1 273.22,247.8
X$40163 219 203 221 3 2 220 MUX2_X1
* cell instance $40313 m0 *1 214.13,250.6
X$40313 235 3 2 153 CLKBUF_X2
* cell instance $40315 m0 *1 216.41,250.6
X$40315 3 720 237 243 236 2 DFF_X1
* cell instance $40316 r0 *1 217.55,247.8
X$40316 210 110 237 3 2 243 MUX2_X1
* cell instance $40322 r0 *1 224.39,247.8
X$40322 210 57 224 3 2 246 MUX2_X1
* cell instance $40326 m0 *1 219.64,250.6
X$40326 238 96 237 3 2 247 MUX2_X1
* cell instance $40330 m0 *1 223.63,250.6
X$40330 3 699 224 246 236 2 DFF_X1
* cell instance $40331 m0 *1 226.86,250.6
X$40331 245 62 247 3 2 232 MUX2_X1
* cell instance $40333 m0 *1 228.38,250.6
X$40333 105 3 2 236 CLKBUF_X3
* cell instance $40334 m0 *1 229.33,250.6
X$40334 236 3 2 CLKBUF_X1
* cell instance $40335 r0 *1 230.09,247.8
X$40335 210 115 211 3 2 225 MUX2_X1
* cell instance $40337 r0 *1 231.42,247.8
X$40337 3 760 211 225 212 2 DFF_X1
* cell instance $40338 r0 *1 234.65,247.8
X$40338 3 757 227 226 212 2 DFF_X1
* cell instance $40345 m0 *1 234.84,250.6
X$40345 211 155 227 3 2 239 MUX2_X1
* cell instance $40346 m0 *1 236.17,250.6
X$40346 105 3 2 212 CLKBUF_X3
* cell instance $40351 m0 *1 241.3,250.6
X$40351 3 693 240 248 212 2 DFF_X1
* cell instance $40353 r0 *1 242.82,247.8
X$40353 153 3 2 79 BUF_X2
* cell instance $40358 r0 *1 255.17,247.8
X$40358 3 756 215 234 172 2 DFF_X1
* cell instance $40361 r0 *1 265.24,247.8
X$40361 3 802 200 218 143 2 DFF_X1
* cell instance $40387 m0 *1 262.01,250.6
X$40387 87 176 84 232 2 3 241 OAI22_X1
* cell instance $40569 m0 *1 213.37,231
X$40569 58 3 2 60 CLKBUF_X2
* cell instance $40571 r0 *1 215.27,228.2
X$40571 49 3 2 51 CLKBUF_X2
* cell instance $40575 r0 *1 222.68,228.2
X$40575 60 52 59 3 2 72 MUX2_X1
* cell instance $40576 r0 *1 219.45,228.2
X$40576 3 759 61 73 50 2 DFF_X1
* cell instance $40578 r0 *1 224.2,228.2
X$40578 60 57 61 3 2 73 MUX2_X1
* cell instance $40579 r0 *1 225.53,228.2
X$40579 59 23 61 3 2 63 MUX2_X1
* cell instance $40586 r0 *1 249.85,228.2
X$40586 25 62 47 3 2 95 MUX2_X1
* cell instance $40607 m0 *1 226.29,231
X$40607 63 62 64 3 2 74 MUX2_X1
* cell instance $40611 m0 *1 234.27,231
X$40611 3 695 99 65 9 2 DFF_X1
* cell instance $40618 m0 *1 241.87,231
X$40618 3 685 67 75 4 2 DFF_X1
* cell instance $40619 m0 *1 245.1,231
X$40619 67 30 79 3 2 75 MUX2_X1
* cell instance $40624 m0 *1 251.94,231
X$40624 3 717 82 92 4 2 DFF_X1
* cell instance $40781 r0 *1 230.85,231
X$40781 89 62 88 3 2 86 MUX2_X1
* cell instance $40783 r0 *1 232.94,231
X$40783 60 3 2 22 BUF_X2
* cell instance $40805 m0 *1 218.5,233.8
X$40805 3 725 113 111 50 2 DFF_X1
* cell instance $40808 m0 *1 224.01,233.8
X$40808 51 110 97 3 2 106 MUX2_X1
* cell instance $40809 m0 *1 225.34,233.8
X$40809 3 700 97 106 50 2 DFF_X1
* cell instance $40810 m0 *1 228.57,233.8
X$40810 98 96 97 3 2 88 MUX2_X1
* cell instance $40815 m0 *1 234.27,233.8
X$40815 8 108 99 3 2 65 MUX2_X1
* cell instance $40816 r0 *1 235.03,231
X$40816 3 766 76 109 9 2 DFF_X1
* cell instance $40818 r0 *1 238.26,231
X$40818 66 62 77 3 2 80 MUX2_X1
* cell instance $40820 m0 *1 235.6,233.8
X$40820 8 110 76 3 2 109 MUX2_X1
* cell instance $40822 m0 *1 237.12,233.8
X$40822 99 96 76 3 2 77 MUX2_X1
* cell instance $40824 r0 *1 243.2,231
X$40824 78 15 79 3 2 91 MUX2_X1
* cell instance $40825 r0 *1 239.97,231
X$40825 3 786 78 91 9 2 DFF_X1
* cell instance $40826 r0 *1 244.53,231
X$40826 67 23 78 3 2 94 MUX2_X1
* cell instance $40829 r0 *1 248.14,231
X$40829 93 62 94 3 2 138 MUX2_X1
* cell instance $40830 r0 *1 249.47,231
X$40830 82 27 100 3 2 93 MUX2_X1
* cell instance $40831 r0 *1 250.8,231
X$40831 87 95 84 74 2 3 81 OAI22_X1
* cell instance $40834 r0 *1 252.7,231
X$40834 82 39 79 3 2 92 MUX2_X1
* cell instance $40845 m0 *1 247.19,233.8
X$40845 3 721 100 107 4 2 DFF_X1
* cell instance $40846 m0 *1 250.42,233.8
X$40846 100 26 79 3 2 107 MUX2_X1
* cell instance $40848 m0 *1 253.27,233.8
X$40848 105 3 2 4 CLKBUF_X3
* cell instance $40849 m0 *1 254.22,233.8
X$40849 4 3 2 836 INV_X2
* cell instance $40852 m0 *1 255.93,233.8
X$40852 118 39 117 3 2 116 MUX2_X1
* cell instance $40854 r0 *1 257.64,231
X$40854 3 770 119 83 11 2 DFF_X1
* cell instance $40856 r0 *1 260.87,231
X$40856 87 90 84 86 2 3 85 OAI22_X1
* cell instance $40861 m0 *1 258.59,233.8
X$40861 119 26 117 3 2 83 MUX2_X1
* cell instance $40863 m0 *1 260.3,233.8
X$40863 105 3 2 11 CLKBUF_X3
* cell instance $40864 m0 *1 261.25,233.8
X$40864 11 3 2 CLKBUF_X1
* cell instance $40865 m0 *1 261.82,233.8
X$40865 87 68 84 80 2 3 121 OAI22_X1
* cell instance $40866 m0 *1 262.77,233.8
X$40866 101 30 117 3 2 104 MUX2_X1
* cell instance $40867 r0 *1 263.15,231
X$40867 3 813 101 104 11 2 DFF_X1
* cell instance $40872 m0 *1 264.86,233.8
X$40872 101 27 102 3 2 120 MUX2_X1
* cell instance $40876 m0 *1 267.52,233.8
X$40876 102 15 117 3 2 103 MUX2_X1
* cell instance $40877 r0 *1 268.47,231
X$40877 3 764 102 103 11 2 DFF_X1
* cell instance $41094 r0 *1 230.47,239.4
X$41094 60 125 139 3 2 148 MUX2_X1
* cell instance $41095 r0 *1 227.24,239.4
X$41095 3 752 139 148 50 2 DFF_X1
* cell instance $41097 r0 *1 233.32,239.4
X$41097 154 187 22 3 2 165 MUX2_X1
* cell instance $41102 r0 *1 248.52,239.4
X$41102 140 155 231 3 2 162 MUX2_X1
* cell instance $41106 r0 *1 254.6,239.4
X$41106 142 132 22 3 2 141 MUX2_X1
* cell instance $41107 r0 *1 255.93,239.4
X$41107 136 158 142 3 2 159 MUX2_X1
* cell instance $41112 m0 *1 231.61,242.2
X$41112 3 694 154 165 9 2 DFF_X1
* cell instance $41115 m0 *1 235.41,242.2
X$41115 124 158 154 3 2 190 MUX2_X1
* cell instance $41117 m0 *1 239.78,242.2
X$41117 127 155 156 3 2 164 MUX2_X1
* cell instance $41121 m0 *1 241.87,242.2
X$41121 129 155 170 3 2 163 MUX2_X1
* cell instance $41126 m0 *1 247.57,242.2
X$41126 150 155 230 3 2 157 MUX2_X1
* cell instance $41127 m0 *1 248.9,242.2
X$41127 157 171 162 3 2 160 MUX2_X1
* cell instance $41135 r0 *1 263.72,239.4
X$41135 147 158 131 3 2 177 MUX2_X1
* cell instance $41137 r0 *1 268.28,239.4
X$41137 144 158 133 3 2 178 MUX2_X1
* cell instance $41334 r0 *1 219.83,250.6
X$41334 210 108 238 3 2 244 MUX2_X1
* cell instance $41335 r0 *1 216.6,250.6
X$41335 3 755 238 244 236 2 DFF_X1
* cell instance $41338 r0 *1 222.11,250.6
X$41338 3 782 257 256 236 2 DFF_X1
* cell instance $41339 r0 *1 225.34,250.6
X$41339 257 23 224 3 2 245 MUX2_X1
* cell instance $41343 r0 *1 230.66,250.6
X$41343 210 3 2 117 BUF_X2
* cell instance $41348 m0 *1 223.25,253.4
X$41348 210 52 257 3 2 256 MUX2_X1
* cell instance $41352 m0 *1 229.9,253.4
X$41352 210 125 249 3 2 276 MUX2_X1
* cell instance $41355 m0 *1 233.13,253.4
X$41355 249 155 279 3 2 259 MUX2_X1
* cell instance $41359 m0 *1 235.79,253.4
X$41359 259 171 239 3 2 260 MUX2_X1
* cell instance $41363 m0 *1 239.78,253.4
X$41363 153 125 250 3 2 261 MUX2_X1
* cell instance $41365 r0 *1 240.92,250.6
X$41365 153 115 240 3 2 248 MUX2_X1
* cell instance $41369 m0 *1 241.3,253.4
X$41369 3 684 250 261 212 2 DFF_X1
* cell instance $41370 m0 *1 244.53,253.4
X$41370 251 213 79 3 2 262 MUX2_X1
* cell instance $41371 r0 *1 248.14,250.6
X$41371 240 158 268 3 2 265 MUX2_X1
* cell instance $41372 r0 *1 244.91,250.6
X$41372 3 758 251 262 212 2 DFF_X1
* cell instance $41378 m0 *1 245.86,253.4
X$41378 250 155 251 3 2 263 MUX2_X1
* cell instance $41382 m0 *1 248.52,253.4
X$41382 263 171 265 3 2 286 MUX2_X1
* cell instance $41385 m0 *1 252.13,253.4
X$41385 79 130 269 3 2 267 MUX2_X1
* cell instance $41386 m0 *1 253.46,253.4
X$41386 3 686 269 267 172 2 DFF_X1
* cell instance $41391 m0 *1 256.88,253.4
X$41391 233 285 3 2 273 OR2_X1
* cell instance $41395 m0 *1 258.97,253.4
X$41395 79 202 271 3 2 266 MUX2_X1
* cell instance $41396 m0 *1 260.3,253.4
X$41396 3 711 271 266 143 2 DFF_X1
* cell instance $41397 m0 *1 263.53,253.4
X$41397 195 260 196 277 2 3 264 OAI22_X1
* cell instance $41398 m0 *1 264.48,253.4
X$41398 241 264 3 2 433 OR2_X1
* cell instance $41400 m0 *1 268.28,253.4
X$41400 275 158 242 3 2 252 MUX2_X1
* cell instance $41401 m0 *1 269.61,253.4
X$41401 252 46 274 3 2 277 MUX2_X1
* cell instance $41402 r0 *1 269.8,250.6
X$41402 242 132 117 3 2 258 MUX2_X1
* cell instance $41404 r0 *1 271.13,250.6
X$41404 3 800 242 258 143 2 DFF_X1
* cell instance $41407 r0 *1 276.07,250.6
X$41407 3 805 253 254 143 2 DFF_X1
* cell instance $41427 m0 *1 273.41,253.4
X$41427 255 217 117 3 2 272 MUX2_X1
* cell instance $41428 m0 *1 274.74,253.4
X$41428 253 203 255 3 2 274 MUX2_X1
* cell instance $41429 m0 *1 276.07,253.4
X$41429 117 202 253 3 2 254 MUX2_X1
* cell instance $41605 r0 *1 212.04,256.2
X$41605 290 3 2 299 CLKBUF_X2
* cell instance $41607 r0 *1 216.6,256.2
X$41607 3 811 308 291 236 2 DFF_X1
* cell instance $41614 m0 *1 216.98,259
X$41614 299 108 308 3 2 291 MUX2_X1
* cell instance $41615 m0 *1 218.31,259
X$41615 299 110 310 3 2 309 MUX2_X1
* cell instance $41618 m0 *1 220.21,259
X$41618 308 96 310 3 2 298 MUX2_X1
* cell instance $41621 r0 *1 223.44,256.2
X$41621 3 790 293 292 236 2 DFF_X1
* cell instance $41646 m0 *1 223.25,259
X$41646 299 52 293 3 2 292 MUX2_X1
* cell instance $41649 m0 *1 225.53,259
X$41649 299 57 295 3 2 294 MUX2_X1
* cell instance $41652 m0 *1 227.81,259
X$41652 293 23 295 3 2 312 MUX2_X1
* cell instance $41653 m0 *1 229.14,259
X$41653 312 62 298 3 2 296 MUX2_X1
* cell instance $41658 m0 *1 237.88,259
X$41658 3 708 301 297 212 2 DFF_X1
* cell instance $41660 m0 *1 241.3,259
X$41660 301 187 316 3 2 297 MUX2_X1
* cell instance $41670 m0 *1 273.79,259
X$41670 3 710 306 311 320 2 DFF_X1
* cell instance $41852 r0 *1 228.95,253.4
X$41852 3 765 249 276 212 2 DFF_X1
* cell instance $41855 r0 *1 232.94,253.4
X$41855 279 213 117 3 2 278 MUX2_X1
* cell instance $41864 m0 *1 231.42,256.2
X$41864 3 691 279 278 212 2 DFF_X1
* cell instance $41869 r0 *1 246.24,253.4
X$41869 3 792 268 281 172 2 DFF_X1
* cell instance $41871 r0 *1 249.47,253.4
X$41871 268 187 79 3 2 281 MUX2_X1
* cell instance $41877 r0 *1 256.69,253.4
X$41877 195 286 196 287 2 3 285 OAI22_X1
* cell instance $41878 r0 *1 253.46,253.4
X$41878 3 788 284 282 172 2 DFF_X1
* cell instance $41879 r0 *1 257.64,253.4
X$41879 270 46 288 3 2 287 MUX2_X1
* cell instance $41883 m0 *1 254.6,256.2
X$41883 284 132 79 3 2 282 MUX2_X1
* cell instance $41888 m0 *1 256.12,256.2
X$41888 269 203 284 3 2 270 MUX2_X1
* cell instance $41890 r0 *1 260.3,253.4
X$41890 271 203 283 3 2 288 MUX2_X1
* cell instance $41894 r0 *1 264.86,253.4
X$41894 3 803 275 280 143 2 DFF_X1
* cell instance $41895 r0 *1 268.09,253.4
X$41895 117 130 275 3 2 280 MUX2_X1
* cell instance $41897 r0 *1 272.46,253.4
X$41897 3 810 255 272 143 2 DFF_X1
* cell instance $41942 m0 *1 260.49,256.2
X$41942 283 217 79 3 2 289 MUX2_X1
* cell instance $41943 m0 *1 261.82,256.2
X$41943 3 712 283 289 314 2 DFF_X1
* cell instance $42072 r0 *1 232.18,236.6
X$42072 3 775 124 135 9 2 DFF_X1
* cell instance $42100 m0 *1 228.57,239.4
X$42100 105 3 2 50 CLKBUF_X3
* cell instance $42101 m0 *1 229.52,239.4
X$42101 50 3 2 837 INV_X2
* cell instance $42105 m0 *1 235.41,239.4
X$42105 105 3 2 9 CLKBUF_X3
* cell instance $42106 m0 *1 236.36,239.4
X$42106 9 3 2 840 INV_X2
* cell instance $42107 r0 *1 239.78,236.6
X$42107 3 769 129 128 9 2 DFF_X1
* cell instance $42108 r0 *1 236.55,236.6
X$42108 3 777 127 126 9 2 DFF_X1
* cell instance $42116 r0 *1 243.58,236.6
X$42116 8 125 150 3 2 151 MUX2_X1
* cell instance $42122 m0 *1 243.96,239.4
X$42122 3 748 150 151 4 2 DFF_X1
* cell instance $42123 m0 *1 247.19,239.4
X$42123 3 746 140 152 4 2 DFF_X1
* cell instance $42125 r0 *1 247.57,236.6
X$42125 8 115 140 3 2 152 MUX2_X1
* cell instance $42128 r0 *1 252.51,236.6
X$42128 22 130 136 3 2 137 MUX2_X1
* cell instance $42130 r0 *1 253.84,236.6
X$42130 3 820 136 137 4 2 DFF_X1
* cell instance $42134 r0 *1 262.39,236.6
X$42134 7 130 147 3 2 149 MUX2_X1
* cell instance $42136 r0 *1 264.48,236.6
X$42136 131 132 7 3 2 146 MUX2_X1
* cell instance $42138 r0 *1 266,236.6
X$42138 3 809 133 134 11 2 DFF_X1
* cell instance $42139 r0 *1 269.23,236.6
X$42139 133 132 38 3 2 134 MUX2_X1
* cell instance $42188 m0 *1 254.03,239.4
X$42188 3 739 142 141 172 2 DFF_X1
* cell instance $42196 m0 *1 261.63,239.4
X$42196 3 734 147 149 143 2 DFF_X1
* cell instance $42197 m0 *1 264.86,239.4
X$42197 3 729 131 146 143 2 DFF_X1
* cell instance $42198 m0 *1 268.09,239.4
X$42198 38 130 144 3 2 145 MUX2_X1
* cell instance $42199 m0 *1 269.42,239.4
X$42199 3 730 144 145 143 2 DFF_X1
.ENDS fwft_fifo

* cell CLKBUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT CLKBUF_X1 1 3 4
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.19,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.38,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.19,0.2075 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.095U AS=0.009975P AD=0.01015P PS=0.4U PD=0.335U
* device instance $4 r0 *1 0.38,0.2575 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.195U AS=0.01015P AD=0.020475P PS=0.335U PD=0.6U
.ENDS CLKBUF_X1

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell NOR3_X2
* pin A3
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 10 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 9 2 10 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 5 3 9 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 8 3 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 4 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 5 1 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 6 2 5 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 5 3 6 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR3_X2

* cell NOR4_X4
* pin PWELL,VSS
* pin A1
* pin A2
* pin A3
* pin A4
* pin ZN
* pin NWELL,VDD
.SUBCKT NOR4_X4 1 2 3 4 5 6 10
* net 1 PWELL,VSS
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 A4
* net 6 ZN
* net 10 NWELL,VDD
* device instance $1 r0 *1 1.92,0.995 PMOS_VTL
M$1 8 4 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 2.68,0.995 PMOS_VTL
M$5 10 5 9 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.995 PMOS_VTL
M$9 6 2 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $13 r0 *1 0.93,0.995 PMOS_VTL
M$13 8 3 7 10 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $17 r0 *1 1.92,0.2975 NMOS_VTL
M$17 1 4 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $21 r0 *1 2.68,0.2975 NMOS_VTL
M$21 1 5 6 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $25 r0 *1 0.17,0.2975 NMOS_VTL
M$25 6 2 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $29 r0 *1 0.93,0.2975 NMOS_VTL
M$29 6 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NOR4_X4

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell AND4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND4_X1 1 2 3 4 6 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 6 2 5 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 5 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 5 4 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 5 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 10 1 5 7 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 11 2 10 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 9 3 11 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 7 4 9 7 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 5 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND4_X1

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.077175P PS=2.24U PD=1.54U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.050925P PS=1.595U
+ PD=1.11U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell OR4_X1
* pin A1
* pin A2
* pin A3
* pin A4
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR4_X1 1 2 3 4 5 7 8
* net 1 A1
* net 2 A2
* net 3 A3
* net 4 A4
* net 5 PWELL,VSS
* net 7 NWELL,VDD
* net 8 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 10 1 6 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 2 10 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 11 3 9 7 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 8 6 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 6 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 5 2 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $8 r0 *1 0.55,0.195 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.74,0.195 NMOS_VTL
M$9 5 4 6 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 8 6 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR4_X1

* cell AOI221_X2
* pin B1
* pin B2
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI221_X2 1 2 3 4 5 6 8 9
* net 1 B1
* net 2 B2
* net 3 A
* net 4 C2
* net 5 C1
* net 6 ZN
* net 8 NWELL,VDD
* net 9 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 3 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.09135P PS=2.24U PD=1.55U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 1 7 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.32,0.995 PMOS_VTL
M$7 6 4 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.09135P AD=0.11025P PS=1.55U PD=2.24U
* device instance $8 r0 *1 1.51,0.995 PMOS_VTL
M$8 10 5 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 6 3 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.060175P PS=1.595U
+ PD=1.12U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 14 1 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 9 2 14 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 13 2 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 6 1 13 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.32,0.2975 NMOS_VTL
M$17 12 4 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P PS=0.565U
+ PD=0.555U
* device instance $18 r0 *1 1.51,0.2975 NMOS_VTL
M$18 6 5 12 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.7,0.2975 NMOS_VTL
M$19 11 5 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.89,0.2975 NMOS_VTL
M$20 9 4 11 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X2

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 0.385,0.32 NMOS_VTL
M$15 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $16 r0 *1 0.575,0.32 NMOS_VTL
M$16 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 0.765,0.32 NMOS_VTL
M$17 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $18 r0 *1 0.96,0.32 NMOS_VTL
M$18 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $19 r0 *1 1.15,0.32 NMOS_VTL
M$19 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $20 r0 *1 0.195,0.2975 NMOS_VTL
M$20 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
* device instance $21 r0 *1 1.49,0.195 NMOS_VTL
M$21 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $22 r0 *1 1.68,0.195 NMOS_VTL
M$22 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $23 r0 *1 1.87,0.195 NMOS_VTL
M$23 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $24 r0 *1 2.06,0.195 NMOS_VTL
M$24 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $25 r0 *1 2.26,0.195 NMOS_VTL
M$25 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $26 r0 *1 2.45,0.195 NMOS_VTL
M$26 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.64,0.195 NMOS_VTL
M$27 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $28 r0 *1 2.83,0.2975 NMOS_VTL
M$28 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS FA_X1

* cell AOI221_X4
* pin PWELL,VSS
* pin ZN
* pin C1
* pin C2
* pin A
* pin B1
* pin B2
* pin NWELL,VDD
.SUBCKT AOI221_X4 1 4 7 8 9 10 11 14
* net 1 PWELL,VSS
* net 4 ZN
* net 7 C1
* net 8 C2
* net 9 A
* net 10 B1
* net 11 B2
* net 14 NWELL,VDD
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 14 11 13 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U
+ PD=0.77U
* device instance $2 r0 *1 1.35,0.995 PMOS_VTL
M$2 3 2 14 14 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $4 r0 *1 1.73,0.995 PMOS_VTL
M$4 4 3 14 14 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $8 r0 *1 0.25,0.995 PMOS_VTL
M$8 2 7 12 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $9 r0 *1 0.44,0.995 PMOS_VTL
M$9 12 8 2 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 0.63,0.995 PMOS_VTL
M$10 13 9 12 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.82,0.995 PMOS_VTL
M$11 14 10 13 14 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $12 r0 *1 0.25,0.2975 NMOS_VTL
M$12 5 7 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $13 r0 *1 0.44,0.2975 NMOS_VTL
M$13 1 8 5 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0342375P PS=0.555U
+ PD=0.58U
* device instance $14 r0 *1 0.655,0.2975 NMOS_VTL
M$14 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.0342375P AD=0.02905P PS=0.58U
+ PD=0.555U
* device instance $15 r0 *1 0.845,0.2975 NMOS_VTL
M$15 6 10 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0549875P PS=0.555U
+ PD=0.68U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 1 11 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.0549875P AD=0.02905P PS=0.68U
+ PD=0.555U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $19 r0 *1 1.73,0.2975 NMOS_VTL
M$19 4 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AOI221_X4

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell NOR4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 3 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 7 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 5 4 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR4_X1

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell AOI21_X4
* pin PWELL,VSS
* pin ZN
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
.SUBCKT AOI21_X4 1 2 3 4 5 11
* net 1 PWELL,VSS
* net 2 ZN
* net 3 A
* net 4 B2
* net 5 B1
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 11 3 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 2 4 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 10 5 2 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 2 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 8 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 2 5 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 9 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 6 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.895,0.2975 NMOS_VTL
M$22 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.085,0.2975 NMOS_VTL
M$23 7 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.275,0.2975 NMOS_VTL
M$24 1 4 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X4

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell OAI221_X1
* pin B2
* pin B1
* pin A
* pin C2
* pin C1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI221_X1 1 2 3 4 5 7 8 9
* net 1 B2
* net 2 B1
* net 3 A
* net 4 C2
* net 5 C1
* net 7 NWELL,VDD
* net 8 PWELL,VSS
* net 9 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 12 1 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 9 2 12 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 9 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 11 4 7 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 5 11 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 8 1 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 6 2 8 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 10 3 6 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 9 4 10 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.93,0.2975 NMOS_VTL
M$10 10 5 9 8 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI221_X1

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X4 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.345,0.195 NMOS_VTL
M$9 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $10 r0 *1 1.535,0.195 NMOS_VTL
M$10 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $11 r0 *1 1.725,0.2975 NMOS_VTL
M$11 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $12 r0 *1 0.785,0.195 NMOS_VTL
M$12 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $13 r0 *1 0.975,0.195 NMOS_VTL
M$13 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $14 r0 *1 0.21,0.2975 NMOS_VTL
M$14 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $15 r0 *1 0.4,0.2975 NMOS_VTL
M$15 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.59,0.2975 NMOS_VTL
M$16 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
.ENDS HA_X1

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell CLKBUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.17,0.1875 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $5 r0 *1 0.36,0.1875 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.39U AS=0.0273P AD=0.034125P PS=0.67U PD=0.935U
.ENDS CLKBUF_X2

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2

* cell DFF_X2
* pin PWELL,VSS
* pin D
* pin CK
* pin QN
* pin Q
* pin NWELL,VDD
.SUBCKT DFF_X2 1 6 8 10 11 16
* net 1 PWELL,VSS
* net 6 D
* net 8 CK
* net 10 QN
* net 11 Q
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.855,0.995 PMOS_VTL
M$1 10 9 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 3.235,0.995 PMOS_VTL
M$3 11 2 16 16 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.2,0.9275 PMOS_VTL
M$5 16 7 3 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $6 r0 *1 0.39,1.04 PMOS_VTL
M$6 17 4 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $7 r0 *1 0.58,1.04 PMOS_VTL
M$7 17 7 5 16 PMOS_VTL L=0.05U W=0.09U AS=0.01785P AD=0.0063P PS=0.56U PD=0.23U
* device instance $8 r0 *1 0.77,0.975 PMOS_VTL
M$8 18 3 5 16 PMOS_VTL L=0.05U W=0.42U AS=0.01785P AD=0.0294P PS=0.56U PD=0.56U
* device instance $9 r0 *1 0.96,0.975 PMOS_VTL
M$9 16 6 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $10 r0 *1 1.15,1.0275 PMOS_VTL
M$10 4 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $11 r0 *1 2.135,0.915 PMOS_VTL
M$11 20 3 9 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $12 r0 *1 2.325,0.915 PMOS_VTL
M$12 20 2 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.0252P AD=0.0063P PS=0.77U PD=0.23U
* device instance $13 r0 *1 1.565,1.0275 PMOS_VTL
M$13 16 8 7 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $14 r0 *1 1.755,1.0275 PMOS_VTL
M$14 19 5 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $15 r0 *1 1.945,1.0275 PMOS_VTL
M$15 9 7 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $16 r0 *1 2.515,0.995 PMOS_VTL
M$16 2 9 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0252P AD=0.06615P PS=0.77U PD=1.47U
* device instance $17 r0 *1 2.855,0.2975 NMOS_VTL
M$17 10 9 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U
+ PD=1.11U
* device instance $19 r0 *1 3.235,0.2975 NMOS_VTL
M$19 11 2 1 1 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U
+ PD=1.595U
* device instance $21 r0 *1 0.39,0.31 NMOS_VTL
M$21 12 4 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $22 r0 *1 0.58,0.31 NMOS_VTL
M$22 12 3 5 1 NMOS_VTL L=0.05U W=0.09U AS=0.012775P AD=0.0063P PS=0.415U
+ PD=0.23U
* device instance $23 r0 *1 1.15,0.25 NMOS_VTL
M$23 4 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $24 r0 *1 0.77,0.2825 NMOS_VTL
M$24 13 7 5 1 NMOS_VTL L=0.05U W=0.275U AS=0.012775P AD=0.01925P PS=0.415U
+ PD=0.415U
* device instance $25 r0 *1 0.96,0.2825 NMOS_VTL
M$25 1 6 13 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
* device instance $26 r0 *1 0.2,0.37 NMOS_VTL
M$26 1 7 3 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $27 r0 *1 1.565,0.35 NMOS_VTL
M$27 1 8 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $28 r0 *1 1.755,0.35 NMOS_VTL
M$28 14 5 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $29 r0 *1 1.945,0.35 NMOS_VTL
M$29 9 3 14 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $30 r0 *1 2.135,0.41 NMOS_VTL
M$30 15 7 9 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $31 r0 *1 2.325,0.41 NMOS_VTL
M$31 15 2 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.017675P AD=0.0063P PS=0.555U
+ PD=0.23U
* device instance $32 r0 *1 2.515,0.2975 NMOS_VTL
M$32 2 9 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.017675P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS DFF_X2

* cell DFF_X1
* pin PWELL,VSS
* pin QN
* pin Q
* pin D
* pin CK
* pin NWELL,VDD
.SUBCKT DFF_X1 1 8 9 14 15 16
* net 1 PWELL,VSS
* net 8 QN
* net 9 Q
* net 14 D
* net 15 CK
* net 16 NWELL,VDD
* device instance $1 r0 *1 2.85,0.995 PMOS_VTL
M$1 16 6 8 16 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 3.04,0.995 PMOS_VTL
M$2 9 7 16 16 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.9425 PMOS_VTL
M$3 16 5 2 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.014175P PS=0.84U
+ PD=0.455U
* device instance $4 r0 *1 0.375,1.055 PMOS_VTL
M$4 17 3 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.0063P PS=0.455U
+ PD=0.23U
* device instance $5 r0 *1 0.565,1.055 PMOS_VTL
M$5 17 5 4 16 PMOS_VTL L=0.05U W=0.09U AS=0.018075P AD=0.0063P PS=0.565U
+ PD=0.23U
* device instance $6 r0 *1 0.76,0.975 PMOS_VTL
M$6 18 2 4 16 PMOS_VTL L=0.05U W=0.42U AS=0.018075P AD=0.0294P PS=0.565U
+ PD=0.56U
* device instance $7 r0 *1 0.95,0.975 PMOS_VTL
M$7 16 14 18 16 PMOS_VTL L=0.05U W=0.42U AS=0.0294P AD=0.025725P PS=0.56U
+ PD=0.56U
* device instance $8 r0 *1 1.14,1.0275 PMOS_VTL
M$8 3 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.025725P AD=0.0567P PS=0.56U
+ PD=0.99U
* device instance $9 r0 *1 1.555,1.0275 PMOS_VTL
M$9 16 15 5 16 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $10 r0 *1 1.745,1.0275 PMOS_VTL
M$10 19 4 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $11 r0 *1 1.935,1.0275 PMOS_VTL
M$11 6 5 19 16 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.014175P PS=0.455U
+ PD=0.455U
* device instance $12 r0 *1 2.125,1.14 PMOS_VTL
M$12 20 2 6 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $13 r0 *1 2.32,1.14 PMOS_VTL
M$13 20 7 16 16 PMOS_VTL L=0.05U W=0.09U AS=0.014175P AD=0.006525P PS=0.455U
+ PD=0.235U
* device instance $14 r0 *1 2.51,1.0275 PMOS_VTL
M$14 7 6 16 16 PMOS_VTL L=0.05U W=0.315U AS=0.014175P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $15 r0 *1 2.85,0.2975 NMOS_VTL
M$15 1 6 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $16 r0 *1 3.04,0.2975 NMOS_VTL
M$16 9 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $17 r0 *1 2.125,0.345 NMOS_VTL
M$17 12 5 6 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $18 r0 *1 2.32,0.345 NMOS_VTL
M$18 12 7 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.006525P PS=0.35U
+ PD=0.235U
* device instance $19 r0 *1 1.555,0.36 NMOS_VTL
M$19 1 15 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $20 r0 *1 1.745,0.36 NMOS_VTL
M$20 13 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $21 r0 *1 1.935,0.36 NMOS_VTL
M$21 6 2 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0105P PS=0.35U PD=0.35U
* device instance $22 r0 *1 2.51,0.36 NMOS_VTL
M$22 7 6 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0105P AD=0.02205P PS=0.35U PD=0.63U
* device instance $23 r0 *1 0.185,0.285 NMOS_VTL
M$23 1 5 2 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0105P PS=0.63U PD=0.35U
* device instance $24 r0 *1 0.375,0.345 NMOS_VTL
M$24 10 3 1 1 NMOS_VTL L=0.05U W=0.09U AS=0.0105P AD=0.0063P PS=0.35U PD=0.23U
* device instance $25 r0 *1 0.565,0.345 NMOS_VTL
M$25 10 2 4 1 NMOS_VTL L=0.05U W=0.09U AS=0.013P AD=0.0063P PS=0.42U PD=0.23U
* device instance $26 r0 *1 1.14,0.285 NMOS_VTL
M$26 3 4 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.016975P AD=0.02205P PS=0.415U
+ PD=0.63U
* device instance $27 r0 *1 0.76,0.3175 NMOS_VTL
M$27 11 5 4 1 NMOS_VTL L=0.05U W=0.275U AS=0.013P AD=0.01925P PS=0.42U PD=0.415U
* device instance $28 r0 *1 0.95,0.3175 NMOS_VTL
M$28 1 14 11 1 NMOS_VTL L=0.05U W=0.275U AS=0.01925P AD=0.016975P PS=0.415U
+ PD=0.415U
.ENDS DFF_X1

* cell OAI22_X1
* pin B2
* pin B1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI22_X1 1 2 3 4 6 7 8
* net 1 B2
* net 2 B1
* net 3 A1
* net 4 A2
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 10 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 8 2 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 9 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 6 4 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.185,0.2975 NMOS_VTL
M$5 7 1 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.375,0.2975 NMOS_VTL
M$6 5 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.565,0.2975 NMOS_VTL
M$7 8 3 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.755,0.2975 NMOS_VTL
M$8 5 4 8 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI22_X1

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1
