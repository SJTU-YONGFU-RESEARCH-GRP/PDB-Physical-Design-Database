module cordic (clk,
    done,
    rst_n,
    start,
    x_in,
    x_out,
    y_in,
    y_out,
    z_in,
    z_out);
 input clk;
 output done;
 input rst_n;
 input start;
 input [15:0] x_in;
 output [15:0] x_out;
 input [15:0] y_in;
 output [15:0] y_out;
 input [15:0] z_in;
 output [15:0] z_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire net2;
 wire net1;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire \iteration[0] ;
 wire \iteration[1] ;
 wire \iteration[2] ;
 wire \iteration[3] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \x[0] ;
 wire \x[10] ;
 wire \x[11] ;
 wire \x[12] ;
 wire \x[13] ;
 wire \x[14] ;
 wire \x[15] ;
 wire \x[1] ;
 wire \x[2] ;
 wire \x[3] ;
 wire \x[4] ;
 wire \x[5] ;
 wire \x[6] ;
 wire \x[7] ;
 wire \x[8] ;
 wire \x[9] ;
 wire \y[0] ;
 wire \y[10] ;
 wire \y[11] ;
 wire \y[12] ;
 wire \y[13] ;
 wire \y[14] ;
 wire \y[15] ;
 wire \y[1] ;
 wire \y[2] ;
 wire \y[3] ;
 wire \y[4] ;
 wire \y[5] ;
 wire \y[6] ;
 wire \y[7] ;
 wire \y[8] ;
 wire \y[9] ;
 wire \z[0] ;
 wire \z[10] ;
 wire \z[11] ;
 wire \z[12] ;
 wire \z[13] ;
 wire \z[14] ;
 wire \z[15] ;
 wire \z[1] ;
 wire \z[2] ;
 wire \z[3] ;
 wire \z[4] ;
 wire \z[5] ;
 wire \z[6] ;
 wire \z[7] ;
 wire \z[8] ;
 wire \z[9] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net102;
 wire net103;
 wire net142;
 wire net105;
 wire net141;
 wire net151;
 wire net148;
 wire net150;
 wire net149;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net145;
 wire net146;
 wire net140;
 wire net143;
 wire net144;
 wire net147;

 CLKBUF_X3 _1279_ (.A(rst_n),
    .Z(_0549_));
 CLKBUF_X3 _1280_ (.A(\state[1] ),
    .Z(_0550_));
 NAND2_X1 _1281_ (.A1(_1120_),
    .A2(_0550_),
    .ZN(_0551_));
 BUF_X4 _1282_ (.A(\iteration[1] ),
    .Z(_0552_));
 CLKBUF_X3 _1283_ (.A(_0552_),
    .Z(_0553_));
 CLKBUF_X3 _1284_ (.A(\state[2] ),
    .Z(_0554_));
 NOR2_X4 _1285_ (.A1(_0554_),
    .A2(_0550_),
    .ZN(_0555_));
 NAND2_X1 _1286_ (.A1(_0553_),
    .A2(_0555_),
    .ZN(_0556_));
 NAND2_X2 _1287_ (.A1(_0556_),
    .A2(_0551_),
    .ZN(_0557_));
 NAND2_X4 _1288_ (.A1(_0549_),
    .A2(_0557_),
    .ZN(_1121_));
 INV_X4 _1289_ (.A(_1121_),
    .ZN(_1130_));
 INV_X1 _1290_ (.A(_0549_),
    .ZN(_0558_));
 BUF_X4 _1291_ (.A(_0558_),
    .Z(_0559_));
 BUF_X2 _1292_ (.A(\state[3] ),
    .Z(_0560_));
 CLKBUF_X3 _1293_ (.A(_0560_),
    .Z(_0561_));
 NOR2_X1 _1294_ (.A1(_0559_),
    .A2(_0561_),
    .ZN(_0562_));
 INV_X1 _1295_ (.A(\state[0] ),
    .ZN(_0563_));
 OAI21_X1 _1296_ (.A(_0562_),
    .B1(net4),
    .B2(_0563_),
    .ZN(_0008_));
 BUF_X4 _1297_ (.A(_0559_),
    .Z(_0564_));
 BUF_X4 _1298_ (.A(_0554_),
    .Z(_0565_));
 BUF_X4 _1299_ (.A(_0565_),
    .Z(_0566_));
 BUF_X4 _1300_ (.A(_0550_),
    .Z(_0567_));
 BUF_X4 _1301_ (.A(_0567_),
    .Z(_0568_));
 BUF_X4 _1302_ (.A(_0568_),
    .Z(_0569_));
 BUF_X4 _1303_ (.A(\iteration[2] ),
    .Z(_0570_));
 INV_X4 _1304_ (.A(_0570_),
    .ZN(_0571_));
 CLKBUF_X3 _1305_ (.A(_0571_),
    .Z(_0572_));
 BUF_X4 _1306_ (.A(\iteration[3] ),
    .Z(_0573_));
 BUF_X4 _1307_ (.A(_0573_),
    .Z(_0574_));
 NAND3_X1 _1308_ (.A1(_0572_),
    .A2(_1119_),
    .A3(_0574_),
    .ZN(_0575_));
 AOI21_X1 _1309_ (.A(_0566_),
    .B1(_0569_),
    .B2(_0575_),
    .ZN(_0576_));
 NOR2_X1 _1310_ (.A1(_0564_),
    .A2(_0576_),
    .ZN(_0009_));
 BUF_X8 _1311_ (.A(\iteration[0] ),
    .Z(_0577_));
 BUF_X8 _1312_ (.A(_0577_),
    .Z(_0578_));
 INV_X1 _1313_ (.A(net2),
    .ZN(_0579_));
 NAND2_X1 _1314_ (.A1(_0550_),
    .A2(_0579_),
    .ZN(_0580_));
 INV_X1 _1315_ (.A(_0555_),
    .ZN(_0581_));
 OAI21_X2 _1316_ (.A(_0580_),
    .B1(_0581_),
    .B2(_0012_),
    .ZN(_0582_));
 NAND2_X2 _1317_ (.A1(_0549_),
    .A2(_0582_),
    .ZN(_1122_));
 INV_X2 _1318_ (.A(_1122_),
    .ZN(_1125_));
 BUF_X2 _1319_ (.A(_0010_),
    .Z(_0583_));
 BUF_X4 _1320_ (.A(_0570_),
    .Z(_0584_));
 BUF_X8 _1321_ (.A(net2),
    .Z(_0585_));
 NAND3_X1 _1322_ (.A1(_0553_),
    .A2(_0584_),
    .A3(_0585_),
    .ZN(_0586_));
 XOR2_X1 _1323_ (.A(_0583_),
    .B(_0586_),
    .Z(_0587_));
 NAND2_X1 _1324_ (.A1(_0567_),
    .A2(_0587_),
    .ZN(_0588_));
 NAND2_X1 _1325_ (.A1(_0574_),
    .A2(_0555_),
    .ZN(_0589_));
 NAND2_X1 _1326_ (.A1(_0588_),
    .A2(_0589_),
    .ZN(_0590_));
 NAND2_X2 _1327_ (.A1(_0549_),
    .A2(_0590_),
    .ZN(_0591_));
 CLKBUF_X3 _1328_ (.A(_0011_),
    .Z(_0592_));
 XNOR2_X2 _1329_ (.A(_0592_),
    .B(_1119_),
    .ZN(_0593_));
 AOI22_X4 _1330_ (.A1(_0584_),
    .A2(_0555_),
    .B1(_0550_),
    .B2(_0593_),
    .ZN(_0594_));
 NOR2_X4 _1331_ (.A1(_0594_),
    .A2(_0558_),
    .ZN(_0038_));
 NOR2_X1 _1332_ (.A1(_1121_),
    .A2(_0038_),
    .ZN(_0595_));
 INV_X1 _1333_ (.A(_0038_),
    .ZN(_0596_));
 NOR2_X1 _1334_ (.A1(_1126_),
    .A2(_0596_),
    .ZN(_0597_));
 OAI21_X1 _1335_ (.A(_0591_),
    .B1(_0595_),
    .B2(_0597_),
    .ZN(_0598_));
 OAI21_X1 _1336_ (.A(_0598_),
    .B1(_0591_),
    .B2(_1124_),
    .ZN(_0000_));
 MUX2_X1 _1337_ (.A(_1122_),
    .B(_0038_),
    .S(_1121_),
    .Z(_0599_));
 MUX2_X1 _1338_ (.A(_1131_),
    .B(_0599_),
    .S(_0591_),
    .Z(_0001_));
 INV_X2 _1339_ (.A(_0591_),
    .ZN(_0039_));
 MUX2_X1 _1340_ (.A(_1128_),
    .B(_0582_),
    .S(_0039_),
    .Z(_0002_));
 NAND4_X1 _1341_ (.A1(_1123_),
    .A2(_0588_),
    .A3(_0589_),
    .A4(_0038_),
    .ZN(_0600_));
 NOR2_X1 _1342_ (.A1(_1123_),
    .A2(_1131_),
    .ZN(_0601_));
 INV_X1 _1343_ (.A(_1131_),
    .ZN(_0602_));
 OAI221_X1 _1344_ (.A(_0600_),
    .B1(_0601_),
    .B2(_0591_),
    .C1(net144),
    .C2(_0602_),
    .ZN(_0003_));
 NAND2_X1 _1345_ (.A1(_1128_),
    .A2(_0039_),
    .ZN(_0603_));
 AOI21_X1 _1346_ (.A(_0595_),
    .B1(net144),
    .B2(_1133_),
    .ZN(_0604_));
 OAI21_X1 _1347_ (.A(_0603_),
    .B1(_0604_),
    .B2(_0039_),
    .ZN(_0004_));
 MUX2_X1 _1348_ (.A(_1124_),
    .B(_1131_),
    .S(_0038_),
    .Z(_0605_));
 MUX2_X1 _1349_ (.A(_0605_),
    .B(_1123_),
    .S(_0039_),
    .Z(_0005_));
 INV_X1 _1350_ (.A(_0025_),
    .ZN(_0606_));
 INV_X1 _1351_ (.A(_0995_),
    .ZN(_0607_));
 BUF_X1 _1352_ (.A(_1005_),
    .Z(_0608_));
 BUF_X1 _1353_ (.A(_1000_),
    .Z(_0609_));
 OR4_X1 _1354_ (.A1(_0609_),
    .A2(_1001_),
    .A3(_1002_),
    .A4(_1003_),
    .ZN(_0610_));
 OR2_X1 _1355_ (.A1(_1004_),
    .A2(_0610_),
    .ZN(_0611_));
 NOR4_X2 _1356_ (.A1(_0608_),
    .A2(_1006_),
    .A3(_0994_),
    .A4(_0611_),
    .ZN(_0612_));
 NAND2_X1 _1357_ (.A1(_0607_),
    .A2(_0612_),
    .ZN(_0613_));
 NOR2_X1 _1358_ (.A1(_0996_),
    .A2(_0613_),
    .ZN(_0614_));
 INV_X1 _1359_ (.A(_0999_),
    .ZN(_0615_));
 NAND2_X2 _1360_ (.A1(_1138_),
    .A2(_0615_),
    .ZN(_0616_));
 NOR2_X1 _1361_ (.A1(_0997_),
    .A2(_0616_),
    .ZN(_0617_));
 AOI21_X1 _1362_ (.A(_0606_),
    .B1(_0614_),
    .B2(_0617_),
    .ZN(_1178_));
 INV_X4 _1363_ (.A(_0573_),
    .ZN(_0618_));
 BUF_X4 _1364_ (.A(_0618_),
    .Z(_0619_));
 CLKBUF_X3 _1365_ (.A(\x[15] ),
    .Z(_0620_));
 BUF_X8 _1366_ (.A(net139),
    .Z(_0621_));
 MUX2_X1 _1367_ (.A(\x[14] ),
    .B(_0620_),
    .S(_0621_),
    .Z(_0622_));
 MUX2_X2 _1368_ (.A(\x[12] ),
    .B(\x[13] ),
    .S(_0621_),
    .Z(_0623_));
 INV_X4 _1369_ (.A(_0552_),
    .ZN(_0624_));
 BUF_X8 _1370_ (.A(_0624_),
    .Z(_0625_));
 MUX2_X2 _1371_ (.A(_0622_),
    .B(_0623_),
    .S(_0625_),
    .Z(_0626_));
 INV_X4 _1372_ (.A(_0626_),
    .ZN(_0627_));
 NOR2_X2 _1373_ (.A1(_0572_),
    .A2(_0627_),
    .ZN(_0628_));
 MUX2_X1 _1374_ (.A(\x[10] ),
    .B(\x[11] ),
    .S(_0621_),
    .Z(_0629_));
 MUX2_X1 _1375_ (.A(\x[8] ),
    .B(\x[9] ),
    .S(_0621_),
    .Z(_0630_));
 MUX2_X1 _1376_ (.A(_0629_),
    .B(_0630_),
    .S(_0625_),
    .Z(_0631_));
 AND2_X4 _1377_ (.A1(_0572_),
    .A2(_0631_),
    .ZN(_0632_));
 NOR2_X4 _1378_ (.A1(_0628_),
    .A2(_0632_),
    .ZN(_0633_));
 NOR2_X1 _1379_ (.A1(_0619_),
    .A2(_0633_),
    .ZN(_0634_));
 MUX2_X1 _1380_ (.A(\x[6] ),
    .B(\x[7] ),
    .S(net1),
    .Z(_0635_));
 MUX2_X1 _1381_ (.A(\x[4] ),
    .B(\x[5] ),
    .S(_0585_),
    .Z(_0636_));
 BUF_X4 _1382_ (.A(_0625_),
    .Z(_0637_));
 MUX2_X1 _1383_ (.A(_0635_),
    .B(_0636_),
    .S(_0637_),
    .Z(_0638_));
 MUX2_X1 _1384_ (.A(\x[2] ),
    .B(\x[3] ),
    .S(_0585_),
    .Z(_0639_));
 MUX2_X1 _1385_ (.A(\x[0] ),
    .B(\x[1] ),
    .S(_0585_),
    .Z(_0640_));
 MUX2_X1 _1386_ (.A(_0639_),
    .B(_0640_),
    .S(_0637_),
    .Z(_0641_));
 MUX2_X1 _1387_ (.A(_0638_),
    .B(_0641_),
    .S(_0572_),
    .Z(_0642_));
 AOI21_X2 _1388_ (.A(_0634_),
    .B1(_0642_),
    .B2(_0619_),
    .ZN(_1186_));
 INV_X1 _1389_ (.A(_1186_),
    .ZN(_1182_));
 BUF_X4 _1390_ (.A(_0637_),
    .Z(_0643_));
 MUX2_X1 _1391_ (.A(_0636_),
    .B(_0639_),
    .S(_0643_),
    .Z(_0644_));
 NOR2_X4 _1392_ (.A1(_0570_),
    .A2(_0573_),
    .ZN(_0645_));
 NOR2_X4 _1393_ (.A1(_0571_),
    .A2(\iteration[3] ),
    .ZN(_0646_));
 MUX2_X1 _1394_ (.A(_0630_),
    .B(_0635_),
    .S(_0643_),
    .Z(_0647_));
 AOI22_X2 _1395_ (.A1(_0644_),
    .A2(_0645_),
    .B1(_0646_),
    .B2(_0647_),
    .ZN(_0648_));
 NOR2_X2 _1396_ (.A1(_0643_),
    .A2(_0584_),
    .ZN(_0649_));
 MUX2_X1 _1397_ (.A(_0622_),
    .B(_0629_),
    .S(_0572_),
    .Z(_0650_));
 AOI22_X4 _1398_ (.A1(net137),
    .A2(_0649_),
    .B1(_0650_),
    .B2(_0643_),
    .ZN(_0651_));
 OAI21_X2 _1399_ (.A(_0648_),
    .B1(_0651_),
    .B2(_0619_),
    .ZN(_0652_));
 BUF_X2 _1400_ (.A(\z[15] ),
    .Z(_0653_));
 BUF_X4 _1401_ (.A(_0653_),
    .Z(_0654_));
 BUF_X4 _1402_ (.A(_0654_),
    .Z(_0655_));
 NOR2_X1 _1403_ (.A1(_0655_),
    .A2(_1187_),
    .ZN(_0656_));
 XNOR2_X1 _1404_ (.A(_0652_),
    .B(_0656_),
    .ZN(_1191_));
 NAND2_X2 _1405_ (.A1(_0571_),
    .A2(_0618_),
    .ZN(_0657_));
 MUX2_X1 _1406_ (.A(\x[5] ),
    .B(\x[6] ),
    .S(_0585_),
    .Z(_0658_));
 MUX2_X1 _1407_ (.A(\x[3] ),
    .B(\x[4] ),
    .S(_0585_),
    .Z(_0659_));
 MUX2_X1 _1408_ (.A(_0658_),
    .B(_0659_),
    .S(_0637_),
    .Z(_0660_));
 NAND2_X4 _1409_ (.A1(_0571_),
    .A2(_0573_),
    .ZN(_0661_));
 MUX2_X1 _1410_ (.A(\x[13] ),
    .B(\x[14] ),
    .S(_0621_),
    .Z(_0662_));
 MUX2_X1 _1411_ (.A(\x[11] ),
    .B(\x[12] ),
    .S(net1),
    .Z(_0663_));
 MUX2_X2 _1412_ (.A(_0662_),
    .B(_0663_),
    .S(_0637_),
    .Z(_0664_));
 OAI22_X2 _1413_ (.A1(_0657_),
    .A2(_0660_),
    .B1(_0661_),
    .B2(_0664_),
    .ZN(_0665_));
 CLKBUF_X2 _1414_ (.A(_0026_),
    .Z(_0666_));
 AND4_X1 _1415_ (.A1(_0579_),
    .A2(_0573_),
    .A3(_0620_),
    .A4(_0666_),
    .ZN(_0667_));
 MUX2_X1 _1416_ (.A(\x[9] ),
    .B(\x[10] ),
    .S(net1),
    .Z(_0668_));
 MUX2_X1 _1417_ (.A(\x[7] ),
    .B(\x[8] ),
    .S(_0585_),
    .Z(_0669_));
 MUX2_X1 _1418_ (.A(_0668_),
    .B(_0669_),
    .S(_0637_),
    .Z(_0670_));
 AOI21_X2 _1419_ (.A(_0667_),
    .B1(_0670_),
    .B2(_0619_),
    .ZN(_0671_));
 AOI21_X4 _1420_ (.A(_0665_),
    .B1(_0671_),
    .B2(_0584_),
    .ZN(_0672_));
 CLKBUF_X3 _1421_ (.A(_0654_),
    .Z(_0673_));
 MUX2_X1 _1422_ (.A(_0631_),
    .B(_0641_),
    .S(_0583_),
    .Z(_0674_));
 MUX2_X1 _1423_ (.A(_0626_),
    .B(_0638_),
    .S(_0583_),
    .Z(_0675_));
 MUX2_X1 _1424_ (.A(_0674_),
    .B(_0675_),
    .S(_0584_),
    .Z(_0676_));
 AND2_X1 _1425_ (.A1(_0625_),
    .A2(_0662_),
    .ZN(_0677_));
 AND3_X1 _1426_ (.A1(_0552_),
    .A2(_0579_),
    .A3(_0620_),
    .ZN(_0678_));
 NOR3_X4 _1427_ (.A1(_0618_),
    .A2(_0677_),
    .A3(_0678_),
    .ZN(_0679_));
 NAND2_X1 _1428_ (.A1(_0637_),
    .A2(_0618_),
    .ZN(_0680_));
 NAND2_X1 _1429_ (.A1(_0553_),
    .A2(_0618_),
    .ZN(_0681_));
 OAI22_X2 _1430_ (.A1(_0658_),
    .A2(_0680_),
    .B1(_0681_),
    .B2(_0669_),
    .ZN(_0682_));
 NOR3_X2 _1431_ (.A1(_0572_),
    .A2(_0679_),
    .A3(_0682_),
    .ZN(_0683_));
 NOR2_X1 _1432_ (.A1(_0643_),
    .A2(_0663_),
    .ZN(_0684_));
 NOR2_X1 _1433_ (.A1(_0553_),
    .A2(_0668_),
    .ZN(_0685_));
 NOR2_X1 _1434_ (.A1(_0643_),
    .A2(_0659_),
    .ZN(_0686_));
 MUX2_X1 _1435_ (.A(\x[1] ),
    .B(\x[2] ),
    .S(_0585_),
    .Z(_0687_));
 NOR2_X1 _1436_ (.A1(_0553_),
    .A2(_0687_),
    .ZN(_0688_));
 OAI33_X1 _1437_ (.A1(_0661_),
    .A2(_0684_),
    .A3(_0685_),
    .B1(_0688_),
    .B2(_0686_),
    .B3(_0657_),
    .ZN(_0689_));
 NOR4_X4 _1438_ (.A1(_0652_),
    .A2(net143),
    .A3(_0683_),
    .A4(net138),
    .ZN(_0690_));
 NOR2_X1 _1439_ (.A1(_0673_),
    .A2(_0690_),
    .ZN(_0691_));
 XNOR2_X1 _1440_ (.A(_0672_),
    .B(_0691_),
    .ZN(_1194_));
 INV_X1 _1441_ (.A(_1183_),
    .ZN(_1110_));
 AOI22_X2 _1442_ (.A1(net136),
    .A2(_0645_),
    .B1(_0646_),
    .B2(_0631_),
    .ZN(_0692_));
 OAI21_X2 _1443_ (.A(_0692_),
    .B1(_0661_),
    .B2(_0627_),
    .ZN(_0693_));
 INV_X2 _1444_ (.A(_0653_),
    .ZN(_0694_));
 INV_X1 _1445_ (.A(_1187_),
    .ZN(_0695_));
 OR2_X4 _1446_ (.A1(_0695_),
    .A2(_0652_),
    .ZN(_0696_));
 OAI21_X4 _1447_ (.A(_0694_),
    .B1(_0672_),
    .B2(_0696_),
    .ZN(_0697_));
 XOR2_X2 _1448_ (.A(_0693_),
    .B(_0697_),
    .Z(_1197_));
 NAND2_X4 _1449_ (.A1(_0570_),
    .A2(_0618_),
    .ZN(_0698_));
 OAI33_X1 _1450_ (.A1(_0679_),
    .A2(_0584_),
    .A3(_0682_),
    .B1(_0684_),
    .B2(_0685_),
    .B3(_0698_),
    .ZN(_0699_));
 NOR2_X1 _1451_ (.A1(_0672_),
    .A2(_0693_),
    .ZN(_0700_));
 AOI21_X2 _1452_ (.A(_0673_),
    .B1(_0690_),
    .B2(_0700_),
    .ZN(_0701_));
 XNOR2_X2 _1453_ (.A(_0699_),
    .B(_0701_),
    .ZN(_1200_));
 NAND4_X1 _1454_ (.A1(_0592_),
    .A2(_0574_),
    .A3(_0666_),
    .A4(_0622_),
    .ZN(_0702_));
 MUX2_X1 _1455_ (.A(_0623_),
    .B(_0629_),
    .S(_0643_),
    .Z(_0703_));
 AOI22_X1 _1456_ (.A1(_0647_),
    .A2(_0645_),
    .B1(_0646_),
    .B2(_0703_),
    .ZN(_0704_));
 NAND2_X1 _1457_ (.A1(_0702_),
    .A2(_0704_),
    .ZN(_0705_));
 NOR4_X4 _1458_ (.A1(_0696_),
    .A2(_0693_),
    .A3(_0672_),
    .A4(net140),
    .ZN(_0706_));
 NOR2_X1 _1459_ (.A1(_0706_),
    .A2(_0673_),
    .ZN(_0707_));
 XNOR2_X1 _1460_ (.A(_0705_),
    .B(_0707_),
    .ZN(_1203_));
 NOR2_X2 _1461_ (.A1(_0552_),
    .A2(net2),
    .ZN(_0708_));
 NAND3_X1 _1462_ (.A1(_0592_),
    .A2(_0620_),
    .A3(_0708_),
    .ZN(_0709_));
 AND2_X1 _1463_ (.A1(_0574_),
    .A2(_0709_),
    .ZN(_0710_));
 MUX2_X1 _1464_ (.A(_0664_),
    .B(_0670_),
    .S(_0572_),
    .Z(_0711_));
 NOR2_X2 _1465_ (.A1(_0574_),
    .A2(_0711_),
    .ZN(_0712_));
 NOR2_X2 _1466_ (.A1(_0710_),
    .A2(_0712_),
    .ZN(_0713_));
 BUF_X4 _1467_ (.A(_0694_),
    .Z(_0714_));
 OR4_X4 _1468_ (.A1(_0652_),
    .A2(net138),
    .A3(_0683_),
    .A4(_0676_),
    .ZN(_0715_));
 OR4_X4 _1469_ (.A1(_0672_),
    .A2(_0693_),
    .A3(net140),
    .A4(_0705_),
    .ZN(_0716_));
 OR2_X4 _1470_ (.A1(_0716_),
    .A2(_0715_),
    .ZN(_0717_));
 NAND2_X4 _1471_ (.A1(_0717_),
    .A2(_0714_),
    .ZN(_0718_));
 XOR2_X2 _1472_ (.A(_0713_),
    .B(_0718_),
    .Z(_1206_));
 OAI21_X2 _1473_ (.A(_0619_),
    .B1(_0628_),
    .B2(_0632_),
    .ZN(_0719_));
 NOR3_X2 _1474_ (.A1(_0696_),
    .A2(_0713_),
    .A3(_0716_),
    .ZN(_0720_));
 NOR2_X1 _1475_ (.A1(_0673_),
    .A2(_0720_),
    .ZN(_0721_));
 XOR2_X2 _1476_ (.A(_0721_),
    .B(_0719_),
    .Z(_1209_));
 MUX2_X1 _1477_ (.A(_0663_),
    .B(_0668_),
    .S(_0625_),
    .Z(_0722_));
 OR2_X1 _1478_ (.A1(_0570_),
    .A2(_0722_),
    .ZN(_0723_));
 OR3_X1 _1479_ (.A1(_0572_),
    .A2(_0677_),
    .A3(_0678_),
    .ZN(_0724_));
 NAND2_X1 _1480_ (.A1(_0723_),
    .A2(_0724_),
    .ZN(_0725_));
 NOR3_X4 _1481_ (.A1(_0715_),
    .A2(_0713_),
    .A3(_0716_),
    .ZN(_0726_));
 AOI21_X1 _1482_ (.A(_0654_),
    .B1(_0633_),
    .B2(_0726_),
    .ZN(_0727_));
 NOR3_X1 _1483_ (.A1(_0727_),
    .A2(_0725_),
    .A3(_0574_),
    .ZN(_0728_));
 INV_X1 _1484_ (.A(_0725_),
    .ZN(_0729_));
 NOR2_X1 _1485_ (.A1(_0574_),
    .A2(_0725_),
    .ZN(_0730_));
 OAI22_X1 _1486_ (.A1(_0719_),
    .A2(_0729_),
    .B1(_0726_),
    .B2(_0730_),
    .ZN(_0731_));
 AOI21_X1 _1487_ (.A(_0728_),
    .B1(_0731_),
    .B2(_0714_),
    .ZN(_1212_));
 OR2_X1 _1488_ (.A1(_0574_),
    .A2(_0651_),
    .ZN(_0732_));
 AOI221_X2 _1489_ (.A(_0632_),
    .B1(_0723_),
    .B2(_0724_),
    .C1(_0626_),
    .C2(_0584_),
    .ZN(_0733_));
 OAI22_X4 _1490_ (.A1(_0710_),
    .A2(_0712_),
    .B1(_0733_),
    .B2(_0574_),
    .ZN(_0734_));
 NOR3_X2 _1491_ (.A1(_0696_),
    .A2(_0716_),
    .A3(_0734_),
    .ZN(_0735_));
 NOR2_X1 _1492_ (.A1(_0673_),
    .A2(_0735_),
    .ZN(_0736_));
 XOR2_X2 _1493_ (.A(_0732_),
    .B(_0736_),
    .Z(_1215_));
 AND3_X1 _1494_ (.A1(_0579_),
    .A2(_0620_),
    .A3(_0666_),
    .ZN(_0737_));
 AOI22_X4 _1495_ (.A1(_0645_),
    .A2(_0664_),
    .B1(_0737_),
    .B2(_0646_),
    .ZN(_0738_));
 NOR2_X1 _1496_ (.A1(_0717_),
    .A2(_0734_),
    .ZN(_0739_));
 AOI21_X1 _1497_ (.A(_0654_),
    .B1(_0732_),
    .B2(_0739_),
    .ZN(_0740_));
 XOR2_X2 _1498_ (.A(_0738_),
    .B(_0740_),
    .Z(_1218_));
 AND2_X1 _1499_ (.A1(_0732_),
    .A2(_0738_),
    .ZN(_0741_));
 AOI21_X2 _1500_ (.A(_0654_),
    .B1(_0735_),
    .B2(_0741_),
    .ZN(_0742_));
 AND2_X1 _1501_ (.A1(_0583_),
    .A2(_0592_),
    .ZN(_0743_));
 NAND2_X1 _1502_ (.A1(_0626_),
    .A2(_0743_),
    .ZN(_0744_));
 XOR2_X2 _1503_ (.A(_0742_),
    .B(_0744_),
    .Z(_1221_));
 NOR2_X1 _1504_ (.A1(_0677_),
    .A2(_0678_),
    .ZN(_0745_));
 NAND2_X2 _1505_ (.A1(_0583_),
    .A2(_0592_),
    .ZN(_0746_));
 NOR2_X1 _1506_ (.A1(_0745_),
    .A2(_0746_),
    .ZN(_0747_));
 OAI221_X2 _1507_ (.A(_0738_),
    .B1(_0746_),
    .B2(_0627_),
    .C1(_0651_),
    .C2(_0574_),
    .ZN(_0748_));
 NOR3_X1 _1508_ (.A1(_0717_),
    .A2(_0734_),
    .A3(_0748_),
    .ZN(_0749_));
 NOR2_X1 _1509_ (.A1(_0673_),
    .A2(_0749_),
    .ZN(_0750_));
 XNOR2_X1 _1510_ (.A(_0747_),
    .B(_0750_),
    .ZN(_1224_));
 AND3_X1 _1511_ (.A1(_0592_),
    .A2(_0618_),
    .A3(_0666_),
    .ZN(_0751_));
 NAND2_X1 _1512_ (.A1(_0622_),
    .A2(_0751_),
    .ZN(_0752_));
 NAND2_X1 _1513_ (.A1(_0694_),
    .A2(_0743_),
    .ZN(_0753_));
 AOI21_X1 _1514_ (.A(_0753_),
    .B1(_0745_),
    .B2(_0627_),
    .ZN(_0754_));
 OR2_X1 _1515_ (.A1(_0742_),
    .A2(_0754_),
    .ZN(_0755_));
 XOR2_X2 _1516_ (.A(_0752_),
    .B(_0755_),
    .Z(_1227_));
 MUX2_X1 _1517_ (.A(\y[10] ),
    .B(\y[11] ),
    .S(_0578_),
    .Z(_0756_));
 OR3_X1 _1518_ (.A1(_0625_),
    .A2(_0570_),
    .A3(_0756_),
    .ZN(_0757_));
 CLKBUF_X3 _1519_ (.A(\y[15] ),
    .Z(_0758_));
 MUX2_X2 _1520_ (.A(\y[14] ),
    .B(_0758_),
    .S(_0577_),
    .Z(_0759_));
 OR3_X1 _1521_ (.A1(_0624_),
    .A2(_0571_),
    .A3(_0759_),
    .ZN(_0760_));
 MUX2_X1 _1522_ (.A(\y[8] ),
    .B(\y[9] ),
    .S(_0578_),
    .Z(_0761_));
 OR3_X2 _1523_ (.A1(_0552_),
    .A2(_0570_),
    .A3(_0761_),
    .ZN(_0762_));
 MUX2_X1 _1524_ (.A(\y[12] ),
    .B(\y[13] ),
    .S(_0578_),
    .Z(_0763_));
 OR3_X2 _1525_ (.A1(_0552_),
    .A2(_0571_),
    .A3(_0763_),
    .ZN(_0764_));
 AND4_X2 _1526_ (.A1(_0757_),
    .A2(_0760_),
    .A3(_0762_),
    .A4(_0764_),
    .ZN(_0765_));
 MUX2_X1 _1527_ (.A(\y[6] ),
    .B(\y[7] ),
    .S(_0578_),
    .Z(_0766_));
 MUX2_X1 _1528_ (.A(\y[4] ),
    .B(\y[5] ),
    .S(_0578_),
    .Z(_0767_));
 MUX2_X1 _1529_ (.A(_0766_),
    .B(_0767_),
    .S(_0624_),
    .Z(_0768_));
 MUX2_X1 _1530_ (.A(\y[2] ),
    .B(\y[3] ),
    .S(net2),
    .Z(_0769_));
 MUX2_X1 _1531_ (.A(\y[0] ),
    .B(\y[1] ),
    .S(net2),
    .Z(_0770_));
 MUX2_X1 _1532_ (.A(_0769_),
    .B(_0770_),
    .S(_0625_),
    .Z(_0771_));
 MUX2_X1 _1533_ (.A(_0768_),
    .B(_0771_),
    .S(_0572_),
    .Z(_0772_));
 MUX2_X1 _1534_ (.A(_0765_),
    .B(_0772_),
    .S(_0619_),
    .Z(_1230_));
 NAND2_X1 _1535_ (.A1(_0714_),
    .A2(_1236_),
    .ZN(_0773_));
 MUX2_X1 _1536_ (.A(\y[13] ),
    .B(\y[14] ),
    .S(net3),
    .Z(_0774_));
 AND2_X1 _1537_ (.A1(_0624_),
    .A2(_0774_),
    .ZN(_0775_));
 AND3_X1 _1538_ (.A1(_0552_),
    .A2(_0579_),
    .A3(_0758_),
    .ZN(_0776_));
 NOR3_X2 _1539_ (.A1(_0618_),
    .A2(_0775_),
    .A3(_0776_),
    .ZN(_0777_));
 MUX2_X1 _1540_ (.A(\y[7] ),
    .B(\y[8] ),
    .S(net3),
    .Z(_0778_));
 MUX2_X1 _1541_ (.A(\y[5] ),
    .B(\y[6] ),
    .S(net1),
    .Z(_0779_));
 OAI22_X2 _1542_ (.A1(_0681_),
    .A2(_0778_),
    .B1(_0779_),
    .B2(_0680_),
    .ZN(_0780_));
 NOR3_X2 _1543_ (.A1(_0572_),
    .A2(_0777_),
    .A3(_0780_),
    .ZN(_0781_));
 MUX2_X1 _1544_ (.A(\y[11] ),
    .B(\y[12] ),
    .S(net3),
    .Z(_0782_));
 NOR2_X1 _1545_ (.A1(_0643_),
    .A2(_0782_),
    .ZN(_0783_));
 MUX2_X1 _1546_ (.A(\y[9] ),
    .B(\y[10] ),
    .S(net3),
    .Z(_0784_));
 NOR2_X1 _1547_ (.A1(_0553_),
    .A2(_0784_),
    .ZN(_0785_));
 MUX2_X1 _1548_ (.A(\y[3] ),
    .B(\y[4] ),
    .S(net1),
    .Z(_0786_));
 NOR2_X1 _1549_ (.A1(_0643_),
    .A2(_0786_),
    .ZN(_0787_));
 MUX2_X1 _1550_ (.A(\y[1] ),
    .B(\y[2] ),
    .S(_0585_),
    .Z(_0788_));
 NOR2_X1 _1551_ (.A1(_0553_),
    .A2(_0788_),
    .ZN(_0789_));
 OAI33_X1 _1552_ (.A1(_0661_),
    .A2(_0783_),
    .A3(_0785_),
    .B1(_0787_),
    .B2(_0789_),
    .B3(_0657_),
    .ZN(_0790_));
 NOR2_X1 _1553_ (.A1(_0781_),
    .A2(_0790_),
    .ZN(_1233_));
 OAI21_X1 _1554_ (.A(_0773_),
    .B1(_1233_),
    .B2(_0025_),
    .ZN(_1237_));
 INV_X1 _1555_ (.A(_1237_),
    .ZN(_1116_));
 NAND2_X1 _1556_ (.A1(_0549_),
    .A2(_0567_),
    .ZN(_0791_));
 NOR2_X1 _1557_ (.A1(_0575_),
    .A2(_0791_),
    .ZN(_0007_));
 BUF_X4 _1558_ (.A(_0549_),
    .Z(_0792_));
 BUF_X2 _1559_ (.A(_0792_),
    .Z(_0793_));
 AND3_X1 _1560_ (.A1(_0793_),
    .A2(\state[0] ),
    .A3(net4),
    .ZN(_0006_));
 INV_X1 _1561_ (.A(_1231_),
    .ZN(_1115_));
 NOR2_X1 _1562_ (.A1(_0683_),
    .A2(_0689_),
    .ZN(_1185_));
 MUX2_X2 _1563_ (.A(_0774_),
    .B(_0782_),
    .S(_0624_),
    .Z(_0794_));
 NAND2_X1 _1564_ (.A1(_0645_),
    .A2(_0794_),
    .ZN(_0795_));
 NAND3_X1 _1565_ (.A1(_0579_),
    .A2(_0666_),
    .A3(_0758_),
    .ZN(_0796_));
 OAI21_X2 _1566_ (.A(_0795_),
    .B1(_0796_),
    .B2(_0698_),
    .ZN(_0797_));
 MUX2_X1 _1567_ (.A(_0765_),
    .B(_0772_),
    .S(_0583_),
    .Z(_0798_));
 MUX2_X2 _1568_ (.A(net105),
    .B(_0756_),
    .S(_0625_),
    .Z(_0799_));
 MUX2_X1 _1569_ (.A(_0767_),
    .B(_0769_),
    .S(_0625_),
    .Z(_0800_));
 OAI22_X2 _1570_ (.A1(_0661_),
    .A2(_0799_),
    .B1(_0800_),
    .B2(_0657_),
    .ZN(_0801_));
 AND3_X1 _1571_ (.A1(_0637_),
    .A2(_0573_),
    .A3(_0759_),
    .ZN(_0802_));
 MUX2_X1 _1572_ (.A(_0761_),
    .B(_0766_),
    .S(_0625_),
    .Z(_0803_));
 AOI21_X2 _1573_ (.A(_0802_),
    .B1(_0803_),
    .B2(_0618_),
    .ZN(_0804_));
 AOI21_X4 _1574_ (.A(_0801_),
    .B1(_0804_),
    .B2(_0584_),
    .ZN(_0805_));
 NOR4_X4 _1575_ (.A1(_0798_),
    .A2(_0790_),
    .A3(_0781_),
    .A4(_0805_),
    .ZN(_0806_));
 AOI22_X2 _1576_ (.A1(_0646_),
    .A2(_0799_),
    .B1(_0803_),
    .B2(_0645_),
    .ZN(_0807_));
 NAND3_X1 _1577_ (.A1(_0592_),
    .A2(_0666_),
    .A3(_0759_),
    .ZN(_0808_));
 OAI21_X2 _1578_ (.A(_0807_),
    .B1(_0808_),
    .B2(_0619_),
    .ZN(_0809_));
 NAND2_X1 _1579_ (.A1(_0645_),
    .A2(_0768_),
    .ZN(_0810_));
 MUX2_X1 _1580_ (.A(_0763_),
    .B(_0759_),
    .S(_0553_),
    .Z(_0811_));
 INV_X1 _1581_ (.A(_0811_),
    .ZN(_0812_));
 MUX2_X1 _1582_ (.A(_0761_),
    .B(_0756_),
    .S(_0553_),
    .Z(_0813_));
 INV_X1 _1583_ (.A(_0813_),
    .ZN(_0814_));
 OAI221_X2 _1584_ (.A(_0810_),
    .B1(_0812_),
    .B2(_0661_),
    .C1(_0698_),
    .C2(_0814_),
    .ZN(_0815_));
 MUX2_X1 _1585_ (.A(_0779_),
    .B(_0786_),
    .S(_0637_),
    .Z(_0816_));
 OAI22_X2 _1586_ (.A1(_0661_),
    .A2(_0794_),
    .B1(_0816_),
    .B2(_0657_),
    .ZN(_0817_));
 AND4_X1 _1587_ (.A1(_0579_),
    .A2(_0573_),
    .A3(_0666_),
    .A4(_0758_),
    .ZN(_0818_));
 MUX2_X1 _1588_ (.A(_0778_),
    .B(_0784_),
    .S(_0552_),
    .Z(_0819_));
 AOI21_X2 _1589_ (.A(_0818_),
    .B1(_0819_),
    .B2(_0618_),
    .ZN(_0820_));
 AOI21_X4 _1590_ (.A(_0817_),
    .B1(_0820_),
    .B2(_0584_),
    .ZN(_0821_));
 OAI33_X1 _1591_ (.A1(_0584_),
    .A2(_0777_),
    .A3(_0780_),
    .B1(_0783_),
    .B2(_0785_),
    .B3(_0698_),
    .ZN(_0822_));
 NOR4_X2 _1592_ (.A1(_0809_),
    .A2(_0815_),
    .A3(_0821_),
    .A4(_0822_),
    .ZN(_0823_));
 AND2_X2 _1593_ (.A1(net134),
    .A2(_0823_),
    .ZN(_0824_));
 NAND2_X1 _1594_ (.A1(_0645_),
    .A2(_0799_),
    .ZN(_0825_));
 NAND2_X1 _1595_ (.A1(_0643_),
    .A2(_0759_),
    .ZN(_0826_));
 OAI21_X4 _1596_ (.A(_0825_),
    .B1(_0826_),
    .B2(_0698_),
    .ZN(_0827_));
 NOR3_X2 _1597_ (.A1(_0553_),
    .A2(_0570_),
    .A3(_0784_),
    .ZN(_0828_));
 NOR3_X2 _1598_ (.A1(_0637_),
    .A2(_0570_),
    .A3(_0782_),
    .ZN(_0829_));
 NOR3_X2 _1599_ (.A1(_0571_),
    .A2(_0775_),
    .A3(_0776_),
    .ZN(_0830_));
 NOR4_X4 _1600_ (.A1(_0573_),
    .A2(_0828_),
    .A3(_0829_),
    .A4(_0830_),
    .ZN(_0831_));
 AND4_X1 _1601_ (.A1(_0592_),
    .A2(_0573_),
    .A3(_0758_),
    .A4(_0708_),
    .ZN(_0832_));
 AOI221_X2 _1602_ (.A(_0832_),
    .B1(_0794_),
    .B2(_0646_),
    .C1(_0645_),
    .C2(_0819_),
    .ZN(_0833_));
 NAND4_X1 _1603_ (.A1(_0757_),
    .A2(_0760_),
    .A3(_0762_),
    .A4(_0764_),
    .ZN(_0834_));
 OAI21_X2 _1604_ (.A(_0833_),
    .B1(_0834_),
    .B2(_0573_),
    .ZN(_0835_));
 NOR3_X1 _1605_ (.A1(_0827_),
    .A2(_0831_),
    .A3(_0835_),
    .ZN(_0836_));
 AOI21_X1 _1606_ (.A(_0654_),
    .B1(_0824_),
    .B2(_0836_),
    .ZN(_0837_));
 XOR2_X2 _1607_ (.A(_0797_),
    .B(_0837_),
    .Z(_1267_));
 NAND2_X1 _1608_ (.A1(_0751_),
    .A2(_0759_),
    .ZN(_0838_));
 INV_X2 _1609_ (.A(_1235_),
    .ZN(_0839_));
 NOR2_X4 _1610_ (.A1(_0805_),
    .A2(_0839_),
    .ZN(_0840_));
 AND2_X1 _1611_ (.A1(_0823_),
    .A2(_0840_),
    .ZN(_0841_));
 OR2_X1 _1612_ (.A1(_0775_),
    .A2(_0776_),
    .ZN(_0842_));
 OAI21_X1 _1613_ (.A(_0743_),
    .B1(_0842_),
    .B2(_0811_),
    .ZN(_0843_));
 NOR4_X4 _1614_ (.A1(_0797_),
    .A2(_0827_),
    .A3(_0831_),
    .A4(_0835_),
    .ZN(_0844_));
 NAND3_X1 _1615_ (.A1(_0841_),
    .A2(_0843_),
    .A3(_0844_),
    .ZN(_0845_));
 NAND2_X1 _1616_ (.A1(_0714_),
    .A2(_0845_),
    .ZN(_0846_));
 XOR2_X2 _1617_ (.A(_0838_),
    .B(_0846_),
    .Z(_1276_));
 NAND2_X1 _1618_ (.A1(_0714_),
    .A2(_1139_),
    .ZN(_0847_));
 OAI21_X2 _1619_ (.A(_0847_),
    .B1(_0714_),
    .B2(_1137_),
    .ZN(_1107_));
 OR2_X1 _1620_ (.A1(_1138_),
    .A2(_0615_),
    .ZN(_0848_));
 AOI21_X1 _1621_ (.A(_0655_),
    .B1(_0616_),
    .B2(_0848_),
    .ZN(_0849_));
 CLKBUF_X3 _1622_ (.A(_0655_),
    .Z(_0850_));
 AOI21_X1 _1623_ (.A(_0849_),
    .B1(_0013_),
    .B2(_0850_),
    .ZN(_1142_));
 BUF_X4 _1624_ (.A(_0654_),
    .Z(_0851_));
 INV_X1 _1625_ (.A(_1136_),
    .ZN(_0852_));
 NOR3_X4 _1626_ (.A1(_0999_),
    .A2(_0998_),
    .A3(_0852_),
    .ZN(_0853_));
 XNOR2_X1 _1627_ (.A(_0609_),
    .B(_0853_),
    .ZN(_0854_));
 NOR2_X1 _1628_ (.A1(_0851_),
    .A2(_0854_),
    .ZN(_0855_));
 AOI21_X1 _1629_ (.A(_0855_),
    .B1(_0014_),
    .B2(_0850_),
    .ZN(_1145_));
 NOR2_X1 _1630_ (.A1(_0609_),
    .A2(_0616_),
    .ZN(_0856_));
 XNOR2_X1 _1631_ (.A(_1001_),
    .B(_0856_),
    .ZN(_0857_));
 NOR2_X1 _1632_ (.A1(_0851_),
    .A2(_0857_),
    .ZN(_0858_));
 AOI21_X1 _1633_ (.A(_0858_),
    .B1(_0015_),
    .B2(_0850_),
    .ZN(_1148_));
 INV_X1 _1634_ (.A(_0853_),
    .ZN(_0859_));
 NOR3_X1 _1635_ (.A1(_0609_),
    .A2(_1001_),
    .A3(_0859_),
    .ZN(_0860_));
 XNOR2_X1 _1636_ (.A(_1002_),
    .B(_0860_),
    .ZN(_0861_));
 NOR2_X1 _1637_ (.A1(_0851_),
    .A2(_0861_),
    .ZN(_0862_));
 AOI21_X1 _1638_ (.A(_0862_),
    .B1(_0016_),
    .B2(_0850_),
    .ZN(_1151_));
 NOR4_X1 _1639_ (.A1(_0609_),
    .A2(_1001_),
    .A3(_1002_),
    .A4(_0616_),
    .ZN(_0863_));
 XNOR2_X1 _1640_ (.A(_1003_),
    .B(_0863_),
    .ZN(_0864_));
 NOR2_X1 _1641_ (.A1(_0851_),
    .A2(_0864_),
    .ZN(_0865_));
 AOI21_X1 _1642_ (.A(_0865_),
    .B1(_0017_),
    .B2(_0850_),
    .ZN(_1154_));
 NOR2_X1 _1643_ (.A1(_0610_),
    .A2(_0859_),
    .ZN(_0866_));
 XNOR2_X1 _1644_ (.A(_1004_),
    .B(_0866_),
    .ZN(_0867_));
 NOR2_X1 _1645_ (.A1(_0655_),
    .A2(_0867_),
    .ZN(_0868_));
 AOI21_X1 _1646_ (.A(_0868_),
    .B1(_0018_),
    .B2(_0850_),
    .ZN(_1157_));
 NOR2_X1 _1647_ (.A1(_0611_),
    .A2(_0616_),
    .ZN(_0869_));
 XNOR2_X1 _1648_ (.A(_0608_),
    .B(_0869_),
    .ZN(_0870_));
 NOR2_X1 _1649_ (.A1(_0655_),
    .A2(_0870_),
    .ZN(_0871_));
 AOI21_X1 _1650_ (.A(_0871_),
    .B1(_0019_),
    .B2(_0850_),
    .ZN(_1160_));
 NOR3_X1 _1651_ (.A1(_0608_),
    .A2(_0611_),
    .A3(_0859_),
    .ZN(_0872_));
 XNOR2_X1 _1652_ (.A(_1006_),
    .B(_0872_),
    .ZN(_0873_));
 NOR2_X1 _1653_ (.A1(_0655_),
    .A2(_0873_),
    .ZN(_0874_));
 AOI21_X1 _1654_ (.A(_0874_),
    .B1(_0020_),
    .B2(_0850_),
    .ZN(_1163_));
 NOR4_X1 _1655_ (.A1(_0608_),
    .A2(_1006_),
    .A3(_0611_),
    .A4(_0616_),
    .ZN(_0875_));
 XNOR2_X1 _1656_ (.A(_0994_),
    .B(_0875_),
    .ZN(_0876_));
 NOR2_X1 _1657_ (.A1(_0655_),
    .A2(_0876_),
    .ZN(_0877_));
 AOI21_X1 _1658_ (.A(_0877_),
    .B1(_0021_),
    .B2(_0850_),
    .ZN(_1166_));
 NAND2_X1 _1659_ (.A1(_0612_),
    .A2(_0853_),
    .ZN(_0878_));
 XNOR2_X1 _1660_ (.A(_0607_),
    .B(_0878_),
    .ZN(_0879_));
 NOR2_X1 _1661_ (.A1(_0655_),
    .A2(_0879_),
    .ZN(_0880_));
 AOI21_X1 _1662_ (.A(_0880_),
    .B1(_0022_),
    .B2(_0850_),
    .ZN(_1169_));
 NOR2_X1 _1663_ (.A1(_0613_),
    .A2(_0616_),
    .ZN(_0881_));
 XNOR2_X1 _1664_ (.A(_0996_),
    .B(_0881_),
    .ZN(_0882_));
 NOR2_X1 _1665_ (.A1(_0655_),
    .A2(_0882_),
    .ZN(_0883_));
 AOI21_X1 _1666_ (.A(_0883_),
    .B1(_0023_),
    .B2(_0851_),
    .ZN(_1172_));
 NAND2_X1 _1667_ (.A1(_0614_),
    .A2(_0853_),
    .ZN(_0884_));
 XOR2_X1 _1668_ (.A(_0997_),
    .B(_0884_),
    .Z(_0885_));
 NOR2_X1 _1669_ (.A1(_0655_),
    .A2(_0885_),
    .ZN(_0886_));
 AOI21_X1 _1670_ (.A(_0886_),
    .B1(_0024_),
    .B2(_0851_),
    .ZN(_1175_));
 NOR2_X1 _1671_ (.A1(_0714_),
    .A2(_1185_),
    .ZN(_0887_));
 AOI21_X2 _1672_ (.A(_0887_),
    .B1(_1188_),
    .B2(_0714_),
    .ZN(_1111_));
 INV_X2 _1673_ (.A(_1230_),
    .ZN(_1234_));
 NAND2_X1 _1674_ (.A1(_0606_),
    .A2(_0805_),
    .ZN(_0888_));
 XNOR2_X1 _1675_ (.A(_0839_),
    .B(_0805_),
    .ZN(_0889_));
 OAI21_X1 _1676_ (.A(_0888_),
    .B1(_0889_),
    .B2(_0851_),
    .ZN(_1240_));
 INV_X1 _1677_ (.A(_0821_),
    .ZN(_0890_));
 XNOR2_X1 _1678_ (.A(net134),
    .B(_0890_),
    .ZN(_0891_));
 OAI22_X2 _1679_ (.A1(_0025_),
    .A2(_0890_),
    .B1(_0891_),
    .B2(_0851_),
    .ZN(_1243_));
 NAND2_X1 _1680_ (.A1(_0606_),
    .A2(_0815_),
    .ZN(_0892_));
 NAND2_X2 _1681_ (.A1(_0840_),
    .A2(_0890_),
    .ZN(_0893_));
 XNOR2_X2 _1682_ (.A(_0893_),
    .B(_0815_),
    .ZN(_0894_));
 OAI21_X2 _1683_ (.A(_0892_),
    .B1(_0851_),
    .B2(_0894_),
    .ZN(_1246_));
 NOR2_X1 _1684_ (.A1(_0815_),
    .A2(_0821_),
    .ZN(_0895_));
 AOI21_X2 _1685_ (.A(_0654_),
    .B1(_0895_),
    .B2(_0806_),
    .ZN(_0896_));
 XOR2_X2 _1686_ (.A(_0822_),
    .B(_0896_),
    .Z(_1249_));
 NOR3_X1 _1687_ (.A1(_0815_),
    .A2(_0821_),
    .A3(_0822_),
    .ZN(_0897_));
 AOI21_X4 _1688_ (.A(_0654_),
    .B1(_0897_),
    .B2(_0840_),
    .ZN(_0898_));
 XOR2_X2 _1689_ (.A(_0809_),
    .B(_0898_),
    .Z(_1252_));
 NOR2_X1 _1690_ (.A1(_0673_),
    .A2(_0824_),
    .ZN(_0899_));
 XNOR2_X1 _1691_ (.A(_0899_),
    .B(_0833_),
    .ZN(_1255_));
 NAND2_X1 _1692_ (.A1(_0619_),
    .A2(_0765_),
    .ZN(_0900_));
 AOI21_X1 _1693_ (.A(_0673_),
    .B1(_0833_),
    .B2(_0841_),
    .ZN(_0901_));
 XNOR2_X1 _1694_ (.A(_0900_),
    .B(_0901_),
    .ZN(_1258_));
 INV_X1 _1695_ (.A(_0824_),
    .ZN(_0902_));
 OAI21_X1 _1696_ (.A(_0714_),
    .B1(_0902_),
    .B2(_0835_),
    .ZN(_0903_));
 XNOR2_X1 _1697_ (.A(_0831_),
    .B(_0903_),
    .ZN(_1261_));
 NOR2_X1 _1698_ (.A1(_0831_),
    .A2(_0835_),
    .ZN(_0904_));
 AOI21_X1 _1699_ (.A(_0654_),
    .B1(_0904_),
    .B2(_0841_),
    .ZN(_0905_));
 XOR2_X2 _1700_ (.A(_0827_),
    .B(_0905_),
    .Z(_1264_));
 NAND2_X1 _1701_ (.A1(_0743_),
    .A2(_0811_),
    .ZN(_0906_));
 AOI21_X1 _1702_ (.A(_0673_),
    .B1(_0841_),
    .B2(_0844_),
    .ZN(_0907_));
 XNOR2_X1 _1703_ (.A(_0906_),
    .B(_0907_),
    .ZN(_1270_));
 NAND3_X1 _1704_ (.A1(net135),
    .A2(_0823_),
    .A3(_0844_),
    .ZN(_0908_));
 OAI21_X1 _1705_ (.A(_0714_),
    .B1(_0811_),
    .B2(_0908_),
    .ZN(_0909_));
 NAND3_X1 _1706_ (.A1(_0743_),
    .A2(_0842_),
    .A3(_0909_),
    .ZN(_0910_));
 NAND3_X1 _1707_ (.A1(_0824_),
    .A2(_0844_),
    .A3(_0906_),
    .ZN(_0911_));
 NOR2_X1 _1708_ (.A1(_0775_),
    .A2(_0776_),
    .ZN(_0912_));
 AOI22_X1 _1709_ (.A1(_0746_),
    .A2(_0908_),
    .B1(_0911_),
    .B2(_0912_),
    .ZN(_0913_));
 OAI21_X1 _1710_ (.A(_0910_),
    .B1(_0913_),
    .B2(_0851_),
    .ZN(_1273_));
 NAND2_X2 _1711_ (.A1(_0591_),
    .A2(_0596_),
    .ZN(_0914_));
 NOR3_X1 _1712_ (.A1(_1121_),
    .A2(_1122_),
    .A3(_0914_),
    .ZN(_0027_));
 NOR2_X1 _1713_ (.A1(_0602_),
    .A2(_0914_),
    .ZN(_0028_));
 INV_X1 _1714_ (.A(_1128_),
    .ZN(_0915_));
 NOR2_X1 _1715_ (.A1(_0915_),
    .A2(_0914_),
    .ZN(_0029_));
 NOR3_X1 _1716_ (.A1(_1130_),
    .A2(_1125_),
    .A3(_0914_),
    .ZN(_0030_));
 NOR2_X1 _1717_ (.A1(_0582_),
    .A2(_0596_),
    .ZN(_0916_));
 NOR2_X1 _1718_ (.A1(_1124_),
    .A2(net144),
    .ZN(_0917_));
 NOR3_X1 _1719_ (.A1(_0039_),
    .A2(_0916_),
    .A3(_0917_),
    .ZN(_0031_));
 AOI21_X1 _1720_ (.A(_0916_),
    .B1(_0596_),
    .B2(_1124_),
    .ZN(_0918_));
 NOR2_X1 _1721_ (.A1(_0039_),
    .A2(_0918_),
    .ZN(_0032_));
 AOI21_X1 _1722_ (.A(_0595_),
    .B1(net144),
    .B2(_1128_),
    .ZN(_0919_));
 NOR2_X1 _1723_ (.A1(_0039_),
    .A2(_0919_),
    .ZN(_0033_));
 OAI21_X1 _1724_ (.A(_0600_),
    .B1(_0914_),
    .B2(_0915_),
    .ZN(_0034_));
 AOI21_X1 _1725_ (.A(_0561_),
    .B1(_0563_),
    .B2(net53),
    .ZN(_0920_));
 NOR2_X1 _1726_ (.A1(_0564_),
    .A2(_0920_),
    .ZN(_0035_));
 NAND2_X1 _1727_ (.A1(_0585_),
    .A2(_0555_),
    .ZN(_0921_));
 AOI21_X1 _1728_ (.A(_0559_),
    .B1(_0580_),
    .B2(_0921_),
    .ZN(_0036_));
 INV_X1 _1729_ (.A(_1121_),
    .ZN(_0037_));
 INV_X1 _1730_ (.A(_0567_),
    .ZN(_0922_));
 BUF_X4 _1731_ (.A(_0922_),
    .Z(_0923_));
 BUF_X4 _1732_ (.A(_0923_),
    .Z(_0924_));
 NOR2_X1 _1733_ (.A1(_0924_),
    .A2(_1232_),
    .ZN(_0925_));
 BUF_X4 _1734_ (.A(_0567_),
    .Z(_0926_));
 BUF_X4 _1735_ (.A(_0565_),
    .Z(_0927_));
 MUX2_X1 _1736_ (.A(\x[0] ),
    .B(net5),
    .S(_0927_),
    .Z(_0928_));
 NOR2_X1 _1737_ (.A1(_0926_),
    .A2(_0928_),
    .ZN(_0929_));
 NOR3_X1 _1738_ (.A1(_0564_),
    .A2(_0925_),
    .A3(_0929_),
    .ZN(_0040_));
 CLKBUF_X3 _1739_ (.A(_0792_),
    .Z(_0930_));
 MUX2_X1 _1740_ (.A(\x[10] ),
    .B(net6),
    .S(_0927_),
    .Z(_0931_));
 OAI21_X1 _1741_ (.A(_0930_),
    .B1(_0569_),
    .B2(_0931_),
    .ZN(_0932_));
 INV_X1 _1742_ (.A(_1262_),
    .ZN(_0933_));
 OR2_X1 _1743_ (.A1(_1256_),
    .A2(_1259_),
    .ZN(_0934_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 NOR3_X1 _1745_ (.A1(_1247_),
    .A2(_1250_),
    .A3(_1253_),
    .ZN(_0936_));
 INV_X1 _1746_ (.A(_1241_),
    .ZN(_0937_));
 INV_X1 _1747_ (.A(_1242_),
    .ZN(_0938_));
 OAI21_X1 _1748_ (.A(_0937_),
    .B1(_0938_),
    .B2(_1117_),
    .ZN(_0939_));
 AOI21_X2 _1749_ (.A(_1244_),
    .B1(_0939_),
    .B2(net141),
    .ZN(_0940_));
 BUF_X1 _1750_ (.A(_1248_),
    .Z(_0941_));
 INV_X1 _1751_ (.A(_0941_),
    .ZN(_0942_));
 OAI21_X1 _1752_ (.A(_0936_),
    .B1(_0940_),
    .B2(_0942_),
    .ZN(_0943_));
 INV_X1 _1753_ (.A(_1257_),
    .ZN(_0944_));
 INV_X1 _1754_ (.A(_1253_),
    .ZN(_0945_));
 BUF_X1 _1755_ (.A(_1251_),
    .Z(_0946_));
 OAI21_X1 _1756_ (.A(_1254_),
    .B1(_1250_),
    .B2(_0946_),
    .ZN(_0947_));
 AOI21_X4 _1757_ (.A(_0944_),
    .B1(_0945_),
    .B2(_0947_),
    .ZN(_0948_));
 AOI21_X2 _1758_ (.A(_0934_),
    .B1(_0943_),
    .B2(_0948_),
    .ZN(_0949_));
 OAI21_X2 _1759_ (.A(_1263_),
    .B1(_1259_),
    .B2(_1260_),
    .ZN(_0950_));
 OAI21_X1 _1760_ (.A(_0933_),
    .B1(_0949_),
    .B2(_0950_),
    .ZN(_0951_));
 XNOR2_X1 _1761_ (.A(_1266_),
    .B(_0951_),
    .ZN(_0952_));
 CLKBUF_X3 _1762_ (.A(_0568_),
    .Z(_0953_));
 AOI21_X1 _1763_ (.A(_0932_),
    .B1(_0952_),
    .B2(_0953_),
    .ZN(_0041_));
 MUX2_X1 _1764_ (.A(\x[11] ),
    .B(net7),
    .S(_0927_),
    .Z(_0954_));
 OAI21_X1 _1765_ (.A(_0930_),
    .B1(_0569_),
    .B2(_0954_),
    .ZN(_0955_));
 OAI21_X1 _1766_ (.A(_1245_),
    .B1(_1241_),
    .B2(_1242_),
    .ZN(_0956_));
 NOR2_X1 _1767_ (.A1(_1238_),
    .A2(_1241_),
    .ZN(_0957_));
 NAND2_X1 _1768_ (.A1(_1231_),
    .A2(_1239_),
    .ZN(_0958_));
 AOI21_X2 _1769_ (.A(_0956_),
    .B1(_0957_),
    .B2(_0958_),
    .ZN(_0959_));
 OR3_X4 _1770_ (.A1(_1253_),
    .A2(_1250_),
    .A3(_1247_),
    .ZN(_0960_));
 OR2_X4 _1771_ (.A1(_0960_),
    .A2(_1244_),
    .ZN(_0961_));
 OAI221_X2 _1772_ (.A(_0948_),
    .B1(_0961_),
    .B2(_0959_),
    .C1(_0960_),
    .C2(_0941_),
    .ZN(_0962_));
 NOR2_X1 _1773_ (.A1(_1262_),
    .A2(_0934_),
    .ZN(_0963_));
 AOI22_X2 _1774_ (.A1(_0933_),
    .A2(_0950_),
    .B1(_0963_),
    .B2(_0962_),
    .ZN(_0964_));
 AOI21_X1 _1775_ (.A(_1265_),
    .B1(_0964_),
    .B2(_1266_),
    .ZN(_0965_));
 XOR2_X1 _1776_ (.A(_1269_),
    .B(_0965_),
    .Z(_0966_));
 AOI21_X1 _1777_ (.A(_0955_),
    .B1(_0966_),
    .B2(_0953_),
    .ZN(_0042_));
 BUF_X1 _1778_ (.A(_1272_),
    .Z(_0967_));
 NOR3_X1 _1779_ (.A1(_1262_),
    .A2(_1265_),
    .A3(_1268_),
    .ZN(_0968_));
 OAI21_X2 _1780_ (.A(_0968_),
    .B1(_0950_),
    .B2(_0949_),
    .ZN(_0969_));
 NOR3_X1 _1781_ (.A1(_1266_),
    .A2(_1265_),
    .A3(_1268_),
    .ZN(_0970_));
 NOR2_X1 _1782_ (.A1(_1269_),
    .A2(_1268_),
    .ZN(_0971_));
 NOR2_X1 _1783_ (.A1(_0970_),
    .A2(_0971_),
    .ZN(_0972_));
 AOI21_X1 _1784_ (.A(_0967_),
    .B1(_0969_),
    .B2(_0972_),
    .ZN(_0973_));
 AND3_X1 _1785_ (.A1(_0967_),
    .A2(_0969_),
    .A3(_0972_),
    .ZN(_0974_));
 OR3_X1 _1786_ (.A1(_0923_),
    .A2(_0973_),
    .A3(_0974_),
    .ZN(_0975_));
 MUX2_X1 _1787_ (.A(\x[12] ),
    .B(net8),
    .S(_0566_),
    .Z(_0976_));
 NAND2_X1 _1788_ (.A1(_0924_),
    .A2(_0976_),
    .ZN(_0977_));
 AOI21_X1 _1789_ (.A(_0559_),
    .B1(_0975_),
    .B2(_0977_),
    .ZN(_0043_));
 BUF_X1 _1790_ (.A(_1275_),
    .Z(_0978_));
 INV_X1 _1791_ (.A(_1271_),
    .ZN(_0979_));
 AND3_X1 _1792_ (.A1(_1269_),
    .A2(_0967_),
    .A3(_1265_),
    .ZN(_0980_));
 AND3_X1 _1793_ (.A1(_1266_),
    .A2(_1269_),
    .A3(_0967_),
    .ZN(_0981_));
 AOI221_X2 _1794_ (.A(_0980_),
    .B1(_0964_),
    .B2(_0981_),
    .C1(_0967_),
    .C2(_1268_),
    .ZN(_0982_));
 NAND2_X1 _1795_ (.A1(_0982_),
    .A2(_0979_),
    .ZN(_0983_));
 XOR2_X1 _1796_ (.A(_0983_),
    .B(_0978_),
    .Z(_0984_));
 NOR2_X1 _1797_ (.A1(_0984_),
    .A2(_0924_),
    .ZN(_0985_));
 MUX2_X1 _1798_ (.A(\x[13] ),
    .B(net9),
    .S(_0927_),
    .Z(_0986_));
 NOR2_X1 _1799_ (.A1(_0926_),
    .A2(_0986_),
    .ZN(_0987_));
 NOR3_X1 _1800_ (.A1(_0985_),
    .A2(_0564_),
    .A3(_0987_),
    .ZN(_0044_));
 NAND2_X1 _1801_ (.A1(_0568_),
    .A2(_1278_),
    .ZN(_0988_));
 AOI21_X1 _1802_ (.A(_1274_),
    .B1(_1271_),
    .B2(_0978_),
    .ZN(_0989_));
 NAND4_X1 _1803_ (.A1(_0967_),
    .A2(_0978_),
    .A3(_0969_),
    .A4(_0972_),
    .ZN(_0990_));
 AOI21_X1 _1804_ (.A(_0988_),
    .B1(_0989_),
    .B2(_0990_),
    .ZN(_0991_));
 INV_X1 _1805_ (.A(_1278_),
    .ZN(_0992_));
 AND4_X1 _1806_ (.A1(_0568_),
    .A2(_0992_),
    .A3(_0990_),
    .A4(_0989_),
    .ZN(_0993_));
 BUF_X4 _1807_ (.A(_0567_),
    .Z(_0136_));
 MUX2_X1 _1808_ (.A(\x[14] ),
    .B(net10),
    .S(_0565_),
    .Z(_0137_));
 OAI21_X1 _1809_ (.A(_0792_),
    .B1(_0136_),
    .B2(_0137_),
    .ZN(_0138_));
 NOR3_X1 _1810_ (.A1(_0991_),
    .A2(_0993_),
    .A3(_0138_),
    .ZN(_0045_));
 NOR3_X1 _1811_ (.A1(_1277_),
    .A2(_0978_),
    .A3(_1274_),
    .ZN(_0139_));
 NOR3_X1 _1812_ (.A1(_1277_),
    .A2(_1271_),
    .A3(_1274_),
    .ZN(_0140_));
 INV_X1 _1813_ (.A(_1277_),
    .ZN(_0141_));
 AOI221_X2 _1814_ (.A(_0139_),
    .B1(_0982_),
    .B2(_0140_),
    .C1(_0141_),
    .C2(_0992_),
    .ZN(_0142_));
 NAND2_X1 _1815_ (.A1(_0142_),
    .A2(_0567_),
    .ZN(_0143_));
 NAND4_X2 _1816_ (.A1(_0592_),
    .A2(_0619_),
    .A3(_0758_),
    .A4(_0708_),
    .ZN(_0144_));
 XNOR2_X2 _1817_ (.A(_0620_),
    .B(_0144_),
    .ZN(_0145_));
 NOR2_X1 _1818_ (.A1(_0653_),
    .A2(_0145_),
    .ZN(_0146_));
 INV_X1 _1819_ (.A(_0146_),
    .ZN(_0147_));
 AOI21_X1 _1820_ (.A(_0147_),
    .B1(_0844_),
    .B2(_0843_),
    .ZN(_0148_));
 AND2_X1 _1821_ (.A1(_0653_),
    .A2(_0145_),
    .ZN(_0149_));
 NOR3_X1 _1822_ (.A1(_0653_),
    .A2(_0838_),
    .A3(_0145_),
    .ZN(_0150_));
 NOR3_X1 _1823_ (.A1(_0148_),
    .A2(_0149_),
    .A3(_0150_),
    .ZN(_0151_));
 NAND4_X1 _1824_ (.A1(_0838_),
    .A2(_0843_),
    .A3(_0844_),
    .A4(_0145_),
    .ZN(_0152_));
 MUX2_X1 _1825_ (.A(_0147_),
    .B(_0152_),
    .S(_0824_),
    .Z(_0153_));
 AOI21_X2 _1826_ (.A(_0143_),
    .B1(_0151_),
    .B2(_0153_),
    .ZN(_0154_));
 MUX2_X1 _1827_ (.A(_0620_),
    .B(net11),
    .S(_0554_),
    .Z(_0155_));
 OAI21_X1 _1828_ (.A(_0792_),
    .B1(_0567_),
    .B2(_0155_),
    .ZN(_0156_));
 AND2_X1 _1829_ (.A1(_0153_),
    .A2(_0151_),
    .ZN(_0157_));
 NOR2_X1 _1830_ (.A1(_0923_),
    .A2(_0142_),
    .ZN(_0158_));
 AOI211_X2 _1831_ (.A(_0156_),
    .B(_0154_),
    .C1(_0157_),
    .C2(_0158_),
    .ZN(_0046_));
 NAND2_X1 _1832_ (.A1(_0568_),
    .A2(_1118_),
    .ZN(_0159_));
 MUX2_X1 _1833_ (.A(\x[1] ),
    .B(net12),
    .S(_0566_),
    .Z(_0160_));
 OAI21_X1 _1834_ (.A(_0159_),
    .B1(_0160_),
    .B2(_0569_),
    .ZN(_0161_));
 NOR2_X1 _1835_ (.A1(_0564_),
    .A2(_0161_),
    .ZN(_0047_));
 XNOR2_X1 _1836_ (.A(_1117_),
    .B(_1242_),
    .ZN(_0162_));
 NOR2_X1 _1837_ (.A1(_0924_),
    .A2(_0162_),
    .ZN(_0163_));
 BUF_X4 _1838_ (.A(_0554_),
    .Z(_0164_));
 MUX2_X1 _1839_ (.A(\x[2] ),
    .B(net13),
    .S(_0164_),
    .Z(_0165_));
 NOR2_X1 _1840_ (.A1(_0926_),
    .A2(_0165_),
    .ZN(_0166_));
 NOR3_X1 _1841_ (.A1(_0564_),
    .A2(_0163_),
    .A3(_0166_),
    .ZN(_0048_));
 AOI21_X1 _1842_ (.A(_1238_),
    .B1(_1239_),
    .B2(_1231_),
    .ZN(_0167_));
 OAI21_X1 _1843_ (.A(_0937_),
    .B1(_0167_),
    .B2(_0938_),
    .ZN(_0168_));
 NOR2_X1 _1844_ (.A1(net142),
    .A2(_0168_),
    .ZN(_0169_));
 OAI21_X1 _1845_ (.A(_0568_),
    .B1(_0959_),
    .B2(_0169_),
    .ZN(_0170_));
 MUX2_X1 _1846_ (.A(\x[3] ),
    .B(net14),
    .S(_0566_),
    .Z(_0171_));
 OAI21_X1 _1847_ (.A(_0170_),
    .B1(_0171_),
    .B2(_0569_),
    .ZN(_0172_));
 NOR2_X1 _1848_ (.A1(_0564_),
    .A2(_0172_),
    .ZN(_0049_));
 XNOR2_X1 _1849_ (.A(_0941_),
    .B(_0940_),
    .ZN(_0173_));
 NOR2_X1 _1850_ (.A1(_0924_),
    .A2(_0173_),
    .ZN(_0174_));
 MUX2_X1 _1851_ (.A(\x[4] ),
    .B(net15),
    .S(_0164_),
    .Z(_0175_));
 NOR2_X1 _1852_ (.A1(_0926_),
    .A2(_0175_),
    .ZN(_0176_));
 NOR3_X1 _1853_ (.A1(_0564_),
    .A2(_0174_),
    .A3(_0176_),
    .ZN(_0050_));
 BUF_X2 _1854_ (.A(_0792_),
    .Z(_0177_));
 MUX2_X1 _1855_ (.A(\x[5] ),
    .B(net16),
    .S(_0565_),
    .Z(_0178_));
 NAND2_X1 _1856_ (.A1(_0923_),
    .A2(_0178_),
    .ZN(_0179_));
 INV_X1 _1857_ (.A(_1247_),
    .ZN(_0180_));
 OAI21_X1 _1858_ (.A(_0941_),
    .B1(_1244_),
    .B2(_0959_),
    .ZN(_0181_));
 NAND2_X1 _1859_ (.A1(_0180_),
    .A2(_0181_),
    .ZN(_0182_));
 XNOR2_X1 _1860_ (.A(_0946_),
    .B(_0182_),
    .ZN(_0183_));
 BUF_X4 _1861_ (.A(_0923_),
    .Z(_0184_));
 OAI21_X1 _1862_ (.A(_0179_),
    .B1(_0183_),
    .B2(_0184_),
    .ZN(_0185_));
 AND2_X1 _1863_ (.A1(_0177_),
    .A2(_0185_),
    .ZN(_0051_));
 BUF_X4 _1864_ (.A(_0559_),
    .Z(_0186_));
 OAI21_X1 _1865_ (.A(_0180_),
    .B1(_0940_),
    .B2(_0942_),
    .ZN(_0187_));
 AOI21_X1 _1866_ (.A(_1250_),
    .B1(_0187_),
    .B2(_0946_),
    .ZN(_0188_));
 XNOR2_X1 _1867_ (.A(_1254_),
    .B(_0188_),
    .ZN(_0189_));
 NOR2_X1 _1868_ (.A1(_0924_),
    .A2(_0189_),
    .ZN(_0190_));
 MUX2_X1 _1869_ (.A(\x[6] ),
    .B(net17),
    .S(_0164_),
    .Z(_0191_));
 NOR2_X1 _1870_ (.A1(_0926_),
    .A2(_0191_),
    .ZN(_0192_));
 NOR3_X1 _1871_ (.A1(_0186_),
    .A2(_0190_),
    .A3(_0192_),
    .ZN(_0052_));
 NOR2_X1 _1872_ (.A1(_1257_),
    .A2(_1253_),
    .ZN(_0193_));
 AOI21_X1 _1873_ (.A(_1250_),
    .B1(_0182_),
    .B2(_0946_),
    .ZN(_0194_));
 INV_X1 _1874_ (.A(_1254_),
    .ZN(_0195_));
 OAI21_X1 _1875_ (.A(_0193_),
    .B1(_0194_),
    .B2(_0195_),
    .ZN(_0196_));
 AOI21_X1 _1876_ (.A(_0184_),
    .B1(net102),
    .B2(_0196_),
    .ZN(_0197_));
 MUX2_X1 _1877_ (.A(\x[7] ),
    .B(net18),
    .S(_0164_),
    .Z(_0198_));
 NOR2_X1 _1878_ (.A1(_0926_),
    .A2(_0198_),
    .ZN(_0199_));
 NOR3_X1 _1879_ (.A1(_0186_),
    .A2(_0197_),
    .A3(_0199_),
    .ZN(_0053_));
 INV_X1 _1880_ (.A(_1256_),
    .ZN(_0200_));
 NAND2_X1 _1881_ (.A1(_0948_),
    .A2(_0943_),
    .ZN(_0201_));
 AND3_X1 _1882_ (.A1(_1260_),
    .A2(_0200_),
    .A3(_0201_),
    .ZN(_0202_));
 AOI21_X1 _1883_ (.A(_1260_),
    .B1(_0200_),
    .B2(_0201_),
    .ZN(_0203_));
 NOR3_X1 _1884_ (.A1(_0184_),
    .A2(_0202_),
    .A3(_0203_),
    .ZN(_0204_));
 MUX2_X1 _1885_ (.A(\x[8] ),
    .B(net19),
    .S(_0164_),
    .Z(_0205_));
 NOR2_X1 _1886_ (.A1(_0926_),
    .A2(_0205_),
    .ZN(_0206_));
 NOR3_X1 _1887_ (.A1(_0186_),
    .A2(_0204_),
    .A3(_0206_),
    .ZN(_0054_));
 CLKBUF_X3 _1888_ (.A(_0923_),
    .Z(_0207_));
 NAND2_X1 _1889_ (.A1(_0200_),
    .A2(net102),
    .ZN(_0208_));
 AOI21_X1 _1890_ (.A(_1259_),
    .B1(_0208_),
    .B2(_1260_),
    .ZN(_0209_));
 XNOR2_X1 _1891_ (.A(_1263_),
    .B(_0209_),
    .ZN(_0210_));
 NOR2_X1 _1892_ (.A1(_0207_),
    .A2(_0210_),
    .ZN(_0211_));
 CLKBUF_X3 _1893_ (.A(_0567_),
    .Z(_0212_));
 MUX2_X1 _1894_ (.A(\x[9] ),
    .B(net20),
    .S(_0164_),
    .Z(_0213_));
 NOR2_X1 _1895_ (.A1(_0212_),
    .A2(_0213_),
    .ZN(_0214_));
 NOR3_X1 _1896_ (.A1(_0186_),
    .A2(_0211_),
    .A3(_0214_),
    .ZN(_0055_));
 MUX2_X1 _1897_ (.A(net54),
    .B(\x[0] ),
    .S(_0561_),
    .Z(_0215_));
 AND2_X1 _1898_ (.A1(_0177_),
    .A2(_0215_),
    .ZN(_0056_));
 MUX2_X1 _1899_ (.A(net55),
    .B(\x[10] ),
    .S(_0561_),
    .Z(_0216_));
 AND2_X1 _1900_ (.A1(_0177_),
    .A2(_0216_),
    .ZN(_0057_));
 MUX2_X1 _1901_ (.A(net56),
    .B(\x[11] ),
    .S(_0561_),
    .Z(_0217_));
 AND2_X1 _1902_ (.A1(_0177_),
    .A2(_0217_),
    .ZN(_0058_));
 MUX2_X1 _1903_ (.A(net57),
    .B(\x[12] ),
    .S(_0561_),
    .Z(_0218_));
 AND2_X1 _1904_ (.A1(_0177_),
    .A2(_0218_),
    .ZN(_0059_));
 MUX2_X1 _1905_ (.A(net58),
    .B(\x[13] ),
    .S(_0561_),
    .Z(_0219_));
 AND2_X1 _1906_ (.A1(_0177_),
    .A2(_0219_),
    .ZN(_0060_));
 MUX2_X1 _1907_ (.A(net59),
    .B(\x[14] ),
    .S(_0561_),
    .Z(_0220_));
 AND2_X1 _1908_ (.A1(_0177_),
    .A2(_0220_),
    .ZN(_0061_));
 MUX2_X1 _1909_ (.A(net60),
    .B(_0620_),
    .S(_0561_),
    .Z(_0221_));
 AND2_X1 _1910_ (.A1(_0177_),
    .A2(_0221_),
    .ZN(_0062_));
 MUX2_X1 _1911_ (.A(net61),
    .B(\x[1] ),
    .S(_0561_),
    .Z(_0222_));
 AND2_X1 _1912_ (.A1(_0177_),
    .A2(_0222_),
    .ZN(_0063_));
 CLKBUF_X3 _1913_ (.A(_0560_),
    .Z(_0223_));
 MUX2_X1 _1914_ (.A(net62),
    .B(\x[2] ),
    .S(_0223_),
    .Z(_0224_));
 AND2_X1 _1915_ (.A1(_0177_),
    .A2(_0224_),
    .ZN(_0064_));
 BUF_X2 _1916_ (.A(_0792_),
    .Z(_0225_));
 MUX2_X1 _1917_ (.A(net63),
    .B(\x[3] ),
    .S(_0223_),
    .Z(_0226_));
 AND2_X1 _1918_ (.A1(_0225_),
    .A2(_0226_),
    .ZN(_0065_));
 MUX2_X1 _1919_ (.A(net64),
    .B(\x[4] ),
    .S(_0223_),
    .Z(_0227_));
 AND2_X1 _1920_ (.A1(_0225_),
    .A2(_0227_),
    .ZN(_0066_));
 MUX2_X1 _1921_ (.A(net65),
    .B(\x[5] ),
    .S(_0223_),
    .Z(_0228_));
 AND2_X1 _1922_ (.A1(_0225_),
    .A2(_0228_),
    .ZN(_0067_));
 MUX2_X1 _1923_ (.A(net66),
    .B(\x[6] ),
    .S(_0223_),
    .Z(_0229_));
 AND2_X1 _1924_ (.A1(_0225_),
    .A2(_0229_),
    .ZN(_0068_));
 MUX2_X1 _1925_ (.A(net67),
    .B(\x[7] ),
    .S(_0223_),
    .Z(_0230_));
 AND2_X1 _1926_ (.A1(_0225_),
    .A2(_0230_),
    .ZN(_0069_));
 MUX2_X1 _1927_ (.A(net68),
    .B(\x[8] ),
    .S(_0223_),
    .Z(_0231_));
 AND2_X1 _1928_ (.A1(_0225_),
    .A2(_0231_),
    .ZN(_0070_));
 MUX2_X1 _1929_ (.A(net69),
    .B(\x[9] ),
    .S(_0223_),
    .Z(_0232_));
 AND2_X1 _1930_ (.A1(_0225_),
    .A2(_0232_),
    .ZN(_0071_));
 NAND2_X1 _1931_ (.A1(_0568_),
    .A2(_1184_),
    .ZN(_0233_));
 MUX2_X1 _1932_ (.A(\y[0] ),
    .B(net21),
    .S(_0566_),
    .Z(_0234_));
 OAI21_X1 _1933_ (.A(_0233_),
    .B1(_0234_),
    .B2(_0569_),
    .ZN(_0235_));
 NOR2_X1 _1934_ (.A1(_0564_),
    .A2(_0235_),
    .ZN(_0072_));
 BUF_X1 _1935_ (.A(_1217_),
    .Z(_0236_));
 BUF_X8 clone2 (.A(_0577_),
    .Z(net2));
 BUF_X4 clone1 (.A(net139),
    .Z(net1));
 OR3_X4 _1938_ (.A1(_1198_),
    .A2(_1201_),
    .A3(_1204_),
    .ZN(_0239_));
 INV_X1 _1939_ (.A(_1195_),
    .ZN(_0240_));
 BUF_X1 _1940_ (.A(_1193_),
    .Z(_0241_));
 AOI21_X1 _1941_ (.A(_1192_),
    .B1(_0241_),
    .B2(_1112_),
    .ZN(_0242_));
 INV_X1 _1942_ (.A(_1196_),
    .ZN(_0243_));
 OAI21_X2 _1943_ (.A(_0240_),
    .B1(_0242_),
    .B2(_0243_),
    .ZN(_0244_));
 AOI21_X4 _1944_ (.A(_0239_),
    .B1(_0244_),
    .B2(net146),
    .ZN(_0245_));
 INV_X1 _1945_ (.A(_1202_),
    .ZN(_0246_));
 INV_X1 _1946_ (.A(_1201_),
    .ZN(_0247_));
 NAND2_X1 _1947_ (.A1(_0246_),
    .A2(_0247_),
    .ZN(_0248_));
 AOI21_X1 _1948_ (.A(_1204_),
    .B1(_0248_),
    .B2(_1205_),
    .ZN(_0249_));
 BUF_X2 _1949_ (.A(_1214_),
    .Z(_0250_));
 NAND3_X2 _1950_ (.A1(_0250_),
    .A2(_1211_),
    .A3(net150),
    .ZN(_0251_));
 OR3_X4 _1951_ (.A1(_0251_),
    .A2(_0249_),
    .A3(_0245_),
    .ZN(_0252_));
 NAND2_X1 _1952_ (.A1(_0250_),
    .A2(_1210_),
    .ZN(_0253_));
 NAND3_X1 _1953_ (.A1(_1211_),
    .A2(_0250_),
    .A3(_1207_),
    .ZN(_0254_));
 NAND3_X4 _1954_ (.A1(_0252_),
    .A2(_0253_),
    .A3(_0254_),
    .ZN(_0255_));
 NOR2_X4 _1955_ (.A1(_1213_),
    .A2(_0255_),
    .ZN(_0256_));
 XNOR2_X2 _1956_ (.A(_0236_),
    .B(_0256_),
    .ZN(_0257_));
 NOR2_X2 _1957_ (.A1(_0207_),
    .A2(_0257_),
    .ZN(_0258_));
 MUX2_X1 _1958_ (.A(\y[10] ),
    .B(net22),
    .S(_0164_),
    .Z(_0259_));
 NOR2_X1 _1959_ (.A1(_0212_),
    .A2(_0259_),
    .ZN(_0260_));
 NOR3_X1 _1960_ (.A1(_0258_),
    .A2(_0186_),
    .A3(_0260_),
    .ZN(_0073_));
 INV_X1 _1961_ (.A(_1220_),
    .ZN(_0261_));
 INV_X1 _1962_ (.A(_1216_),
    .ZN(_0262_));
 INV_X1 _1963_ (.A(_1211_),
    .ZN(_0263_));
 INV_X1 _1964_ (.A(_1207_),
    .ZN(_0264_));
 OAI21_X1 _1965_ (.A(_1208_),
    .B1(_1205_),
    .B2(_1204_),
    .ZN(_0265_));
 AOI21_X1 _1966_ (.A(_0263_),
    .B1(_0264_),
    .B2(_0265_),
    .ZN(_0266_));
 OR2_X2 _1967_ (.A1(_1210_),
    .A2(_0266_),
    .ZN(_0267_));
 NOR3_X1 _1968_ (.A1(_1204_),
    .A2(_1207_),
    .A3(_1210_),
    .ZN(_0268_));
 OR3_X4 _1969_ (.A1(_1195_),
    .A2(_1198_),
    .A3(_1201_),
    .ZN(_0269_));
 OAI21_X1 _1970_ (.A(_1196_),
    .B1(_1192_),
    .B2(_0241_),
    .ZN(_0270_));
 INV_X1 _1971_ (.A(_0270_),
    .ZN(_0271_));
 NOR2_X1 _1972_ (.A1(_1189_),
    .A2(_1192_),
    .ZN(_0272_));
 INV_X1 _1973_ (.A(_1190_),
    .ZN(_0273_));
 OAI21_X1 _1974_ (.A(_0272_),
    .B1(_0273_),
    .B2(_1183_),
    .ZN(_0274_));
 AOI21_X4 _1975_ (.A(_0269_),
    .B1(_0271_),
    .B2(_0274_),
    .ZN(_0275_));
 OAI21_X1 _1976_ (.A(_1202_),
    .B1(_1198_),
    .B2(_1199_),
    .ZN(_0276_));
 AND2_X1 _1977_ (.A1(_0247_),
    .A2(_0276_),
    .ZN(_0277_));
 OAI21_X2 _1978_ (.A(_0268_),
    .B1(_0275_),
    .B2(_0277_),
    .ZN(_0278_));
 AND3_X4 _1979_ (.A1(_0267_),
    .A2(_0250_),
    .A3(_0278_),
    .ZN(_0279_));
 OAI21_X1 _1980_ (.A(_0236_),
    .B1(_1213_),
    .B2(_0279_),
    .ZN(_0280_));
 NAND3_X1 _1981_ (.A1(_0261_),
    .A2(_0262_),
    .A3(_0280_),
    .ZN(_0281_));
 OR2_X1 _1982_ (.A1(_1213_),
    .A2(_1216_),
    .ZN(_0282_));
 OAI221_X2 _1983_ (.A(_1220_),
    .B1(_0282_),
    .B2(_0279_),
    .C1(_1216_),
    .C2(_0236_),
    .ZN(_0283_));
 AOI21_X2 _1984_ (.A(_0923_),
    .B1(_0281_),
    .B2(_0283_),
    .ZN(_0284_));
 MUX2_X1 _1985_ (.A(\y[11] ),
    .B(net23),
    .S(_0164_),
    .Z(_0285_));
 NOR2_X1 _1986_ (.A1(_0212_),
    .A2(_0285_),
    .ZN(_0286_));
 NOR3_X1 _1987_ (.A1(_0284_),
    .A2(_0186_),
    .A3(_0286_),
    .ZN(_0074_));
 BUF_X1 _1988_ (.A(_1223_),
    .Z(_0287_));
 INV_X1 _1989_ (.A(_1219_),
    .ZN(_0288_));
 NOR2_X1 _1990_ (.A1(_0236_),
    .A2(_1216_),
    .ZN(_0289_));
 OAI21_X1 _1991_ (.A(_0288_),
    .B1(_0289_),
    .B2(_0261_),
    .ZN(_0290_));
 OR2_X1 _1992_ (.A1(_1219_),
    .A2(_0282_),
    .ZN(_0291_));
 OAI21_X4 _1993_ (.A(_0290_),
    .B1(_0291_),
    .B2(_0255_),
    .ZN(_0292_));
 XNOR2_X2 _1994_ (.A(_0292_),
    .B(_0287_),
    .ZN(_0293_));
 NOR2_X2 _1995_ (.A1(_0293_),
    .A2(_0207_),
    .ZN(_0294_));
 MUX2_X1 _1996_ (.A(\y[12] ),
    .B(net24),
    .S(_0164_),
    .Z(_0295_));
 NOR2_X1 _1997_ (.A1(_0212_),
    .A2(_0295_),
    .ZN(_0296_));
 NOR3_X1 _1998_ (.A1(_0294_),
    .A2(_0186_),
    .A3(_0296_),
    .ZN(_0075_));
 INV_X1 _1999_ (.A(_1226_),
    .ZN(_0297_));
 NOR2_X1 _2000_ (.A1(_0923_),
    .A2(_0297_),
    .ZN(_0298_));
 INV_X1 _2001_ (.A(_0287_),
    .ZN(_0299_));
 AOI21_X2 _2002_ (.A(_0299_),
    .B1(_0283_),
    .B2(_0288_),
    .ZN(_0300_));
 OAI21_X1 _2003_ (.A(_0298_),
    .B1(_0300_),
    .B2(_1222_),
    .ZN(_0301_));
 OR4_X4 _2004_ (.A1(_0300_),
    .A2(_1226_),
    .A3(_1222_),
    .A4(_0922_),
    .ZN(_0302_));
 MUX2_X1 _2005_ (.A(\y[13] ),
    .B(net25),
    .S(_0565_),
    .Z(_0303_));
 OR2_X1 _2006_ (.A1(_0568_),
    .A2(_0303_),
    .ZN(_0304_));
 AND4_X4 _2007_ (.A1(_0302_),
    .A2(_0301_),
    .A3(_0930_),
    .A4(_0304_),
    .ZN(_0076_));
 MUX2_X1 _2008_ (.A(\y[14] ),
    .B(net26),
    .S(_0927_),
    .Z(_0305_));
 OAI21_X1 _2009_ (.A(_0930_),
    .B1(_0569_),
    .B2(_0305_),
    .ZN(_0306_));
 INV_X1 _2010_ (.A(_1225_),
    .ZN(_0307_));
 NAND2_X1 _2011_ (.A1(_0287_),
    .A2(_1226_),
    .ZN(_0308_));
 INV_X1 _2012_ (.A(_1222_),
    .ZN(_0309_));
 OAI221_X2 _2013_ (.A(_0307_),
    .B1(_0292_),
    .B2(_0308_),
    .C1(_0309_),
    .C2(_0297_),
    .ZN(_0310_));
 XNOR2_X1 _2014_ (.A(_0310_),
    .B(_1229_),
    .ZN(_0311_));
 AOI21_X1 _2015_ (.A(_0306_),
    .B1(_0311_),
    .B2(_0953_),
    .ZN(_0077_));
 MUX2_X1 _2016_ (.A(_0758_),
    .B(net27),
    .S(_0927_),
    .Z(_0312_));
 OAI21_X1 _2017_ (.A(_0930_),
    .B1(_0569_),
    .B2(_0312_),
    .ZN(_0313_));
 NAND4_X2 _2018_ (.A1(_0592_),
    .A2(_0619_),
    .A3(_0620_),
    .A4(_0708_),
    .ZN(_0314_));
 XOR2_X2 _2019_ (.A(_0758_),
    .B(_0314_),
    .Z(_0315_));
 OAI21_X1 _2020_ (.A(_0752_),
    .B1(_0746_),
    .B2(_0745_),
    .ZN(_0316_));
 OR3_X1 _2021_ (.A1(_0748_),
    .A2(_0315_),
    .A3(_0316_),
    .ZN(_0317_));
 OR4_X1 _2022_ (.A1(_0715_),
    .A2(_0716_),
    .A3(_0734_),
    .A4(_0317_),
    .ZN(_0318_));
 AND2_X1 _2023_ (.A1(_0694_),
    .A2(_0315_),
    .ZN(_0319_));
 OAI21_X1 _2024_ (.A(_0319_),
    .B1(_0716_),
    .B2(_0715_),
    .ZN(_0320_));
 NAND2_X1 _2025_ (.A1(_0734_),
    .A2(_0319_),
    .ZN(_0321_));
 NOR2_X1 _2026_ (.A1(_0694_),
    .A2(_0315_),
    .ZN(_0322_));
 AND2_X1 _2027_ (.A1(_0315_),
    .A2(_0316_),
    .ZN(_0323_));
 AOI221_X2 _2028_ (.A(_0322_),
    .B1(_0323_),
    .B2(_0694_),
    .C1(_0748_),
    .C2(_0319_),
    .ZN(_0324_));
 NAND4_X1 _2029_ (.A1(_0318_),
    .A2(_0320_),
    .A3(_0321_),
    .A4(_0324_),
    .ZN(_0325_));
 AOI21_X1 _2030_ (.A(_1222_),
    .B1(_1219_),
    .B2(_0287_),
    .ZN(_0326_));
 OAI21_X1 _2031_ (.A(_0307_),
    .B1(_0326_),
    .B2(_0297_),
    .ZN(_0327_));
 AOI21_X1 _2032_ (.A(_1228_),
    .B1(_0327_),
    .B2(_1229_),
    .ZN(_0328_));
 NAND3_X1 _2033_ (.A1(_0287_),
    .A2(_1226_),
    .A3(_1229_),
    .ZN(_0329_));
 OAI21_X2 _2034_ (.A(_0328_),
    .B1(net149),
    .B2(_0329_),
    .ZN(_0330_));
 XOR2_X1 _2035_ (.A(_0325_),
    .B(_0330_),
    .Z(_0331_));
 AOI21_X1 _2036_ (.A(_0313_),
    .B1(_0953_),
    .B2(_0331_),
    .ZN(_0078_));
 NOR2_X1 _2037_ (.A1(_0207_),
    .A2(_1113_),
    .ZN(_0332_));
 MUX2_X1 _2038_ (.A(\y[1] ),
    .B(net28),
    .S(_0164_),
    .Z(_0333_));
 NOR2_X1 _2039_ (.A1(_0212_),
    .A2(_0333_),
    .ZN(_0334_));
 NOR3_X1 _2040_ (.A1(_0186_),
    .A2(_0332_),
    .A3(_0334_),
    .ZN(_0079_));
 XOR2_X1 _2041_ (.A(_1112_),
    .B(_0241_),
    .Z(_0335_));
 NOR2_X1 _2042_ (.A1(_0207_),
    .A2(_0335_),
    .ZN(_0336_));
 BUF_X4 _2043_ (.A(_0554_),
    .Z(_0337_));
 MUX2_X1 _2044_ (.A(\y[2] ),
    .B(net29),
    .S(_0337_),
    .Z(_0338_));
 NOR2_X1 _2045_ (.A1(_0212_),
    .A2(_0338_),
    .ZN(_0339_));
 NOR3_X1 _2046_ (.A1(_0186_),
    .A2(_0336_),
    .A3(_0339_),
    .ZN(_0080_));
 INV_X1 _2047_ (.A(_1189_),
    .ZN(_0340_));
 OAI21_X1 _2048_ (.A(_0340_),
    .B1(_0273_),
    .B2(_1183_),
    .ZN(_0341_));
 AOI21_X1 _2049_ (.A(_1192_),
    .B1(_0341_),
    .B2(_0241_),
    .ZN(_0342_));
 XNOR2_X1 _2050_ (.A(net145),
    .B(_0342_),
    .ZN(_0343_));
 NOR2_X1 _2051_ (.A1(_0207_),
    .A2(_0343_),
    .ZN(_0344_));
 MUX2_X1 _2052_ (.A(\y[3] ),
    .B(net30),
    .S(_0337_),
    .Z(_0345_));
 NOR2_X1 _2053_ (.A1(_0212_),
    .A2(_0345_),
    .ZN(_0346_));
 NOR3_X1 _2054_ (.A1(_0186_),
    .A2(_0344_),
    .A3(_0346_),
    .ZN(_0081_));
 BUF_X4 _2055_ (.A(_0559_),
    .Z(_0347_));
 INV_X1 _2056_ (.A(_1199_),
    .ZN(_0348_));
 XNOR2_X1 _2057_ (.A(_0348_),
    .B(_0244_),
    .ZN(_0349_));
 NOR2_X1 _2058_ (.A1(_0207_),
    .A2(_0349_),
    .ZN(_0350_));
 MUX2_X1 _2059_ (.A(\y[4] ),
    .B(net31),
    .S(_0337_),
    .Z(_0351_));
 NOR2_X1 _2060_ (.A1(_0212_),
    .A2(_0351_),
    .ZN(_0352_));
 NOR3_X1 _2061_ (.A1(_0347_),
    .A2(_0350_),
    .A3(_0352_),
    .ZN(_0082_));
 AOI21_X1 _2062_ (.A(_1195_),
    .B1(_0274_),
    .B2(_0271_),
    .ZN(_0353_));
 NOR2_X1 _2063_ (.A1(_0348_),
    .A2(_0353_),
    .ZN(_0354_));
 NOR2_X1 _2064_ (.A1(_1198_),
    .A2(_0354_),
    .ZN(_0355_));
 XNOR2_X1 _2065_ (.A(_1202_),
    .B(_0355_),
    .ZN(_0356_));
 NOR2_X1 _2066_ (.A1(_0207_),
    .A2(_0356_),
    .ZN(_0357_));
 MUX2_X1 _2067_ (.A(\y[5] ),
    .B(net32),
    .S(_0337_),
    .Z(_0358_));
 NOR2_X1 _2068_ (.A1(_0212_),
    .A2(_0358_),
    .ZN(_0359_));
 NOR3_X1 _2069_ (.A1(_0347_),
    .A2(_0357_),
    .A3(_0359_),
    .ZN(_0083_));
 INV_X1 _2070_ (.A(_1205_),
    .ZN(_0360_));
 AOI21_X1 _2071_ (.A(_1198_),
    .B1(_0244_),
    .B2(_1199_),
    .ZN(_0361_));
 OAI21_X1 _2072_ (.A(_0247_),
    .B1(_0361_),
    .B2(_0246_),
    .ZN(_0362_));
 XNOR2_X1 _2073_ (.A(_0360_),
    .B(_0362_),
    .ZN(_0363_));
 NAND2_X1 _2074_ (.A1(_0953_),
    .A2(_0363_),
    .ZN(_0364_));
 MUX2_X1 _2075_ (.A(\y[6] ),
    .B(net33),
    .S(_0566_),
    .Z(_0365_));
 NAND2_X1 _2076_ (.A1(_0924_),
    .A2(_0365_),
    .ZN(_0366_));
 AOI21_X1 _2077_ (.A(_0559_),
    .B1(_0364_),
    .B2(_0366_),
    .ZN(_0084_));
 INV_X1 _2078_ (.A(net151),
    .ZN(_0367_));
 NOR3_X1 _2079_ (.A1(_0360_),
    .A2(_0277_),
    .A3(_0275_),
    .ZN(_0368_));
 OR2_X1 _2080_ (.A1(_1204_),
    .A2(_0368_),
    .ZN(_0369_));
 XNOR2_X1 _2081_ (.A(_0367_),
    .B(_0369_),
    .ZN(_0370_));
 NOR2_X1 _2082_ (.A1(_0207_),
    .A2(_0370_),
    .ZN(_0371_));
 MUX2_X1 _2083_ (.A(\y[7] ),
    .B(net34),
    .S(_0337_),
    .Z(_0372_));
 NOR2_X1 _2084_ (.A1(_0212_),
    .A2(_0372_),
    .ZN(_0373_));
 NOR3_X1 _2085_ (.A1(_0347_),
    .A2(_0371_),
    .A3(_0373_),
    .ZN(_0085_));
 MUX2_X1 _2086_ (.A(\y[8] ),
    .B(net35),
    .S(_0927_),
    .Z(_0374_));
 OAI21_X1 _2087_ (.A(_0930_),
    .B1(_0926_),
    .B2(_0374_),
    .ZN(_0375_));
 NOR3_X1 _2088_ (.A1(_0367_),
    .A2(_0245_),
    .A3(_0249_),
    .ZN(_0376_));
 NOR2_X1 _2089_ (.A1(_1207_),
    .A2(_0376_),
    .ZN(_0377_));
 XNOR2_X1 _2090_ (.A(_0263_),
    .B(_0377_),
    .ZN(_0378_));
 AOI21_X1 _2091_ (.A(_0375_),
    .B1(_0378_),
    .B2(_0953_),
    .ZN(_0086_));
 MUX2_X1 _2092_ (.A(\y[9] ),
    .B(net36),
    .S(_0565_),
    .Z(_0379_));
 OR2_X1 _2093_ (.A1(_0568_),
    .A2(_0379_),
    .ZN(_0380_));
 AOI21_X1 _2094_ (.A(_0250_),
    .B1(_0267_),
    .B2(_0278_),
    .ZN(_0381_));
 OAI21_X1 _2095_ (.A(_0136_),
    .B1(_0279_),
    .B2(_0381_),
    .ZN(_0382_));
 AND3_X1 _2096_ (.A1(_0930_),
    .A2(_0380_),
    .A3(_0382_),
    .ZN(_0087_));
 MUX2_X1 _2097_ (.A(net70),
    .B(\y[0] ),
    .S(_0223_),
    .Z(_0383_));
 AND2_X1 _2098_ (.A1(_0225_),
    .A2(_0383_),
    .ZN(_0088_));
 MUX2_X1 _2099_ (.A(net71),
    .B(\y[10] ),
    .S(_0223_),
    .Z(_0384_));
 AND2_X1 _2100_ (.A1(_0225_),
    .A2(_0384_),
    .ZN(_0089_));
 BUF_X4 _2101_ (.A(_0560_),
    .Z(_0385_));
 MUX2_X1 _2102_ (.A(net72),
    .B(\y[11] ),
    .S(_0385_),
    .Z(_0386_));
 AND2_X1 _2103_ (.A1(_0225_),
    .A2(_0386_),
    .ZN(_0090_));
 BUF_X2 _2104_ (.A(_0792_),
    .Z(_0387_));
 MUX2_X1 _2105_ (.A(net73),
    .B(\y[12] ),
    .S(_0385_),
    .Z(_0388_));
 AND2_X1 _2106_ (.A1(_0387_),
    .A2(_0388_),
    .ZN(_0091_));
 MUX2_X1 _2107_ (.A(net74),
    .B(\y[13] ),
    .S(_0385_),
    .Z(_0389_));
 AND2_X1 _2108_ (.A1(_0387_),
    .A2(_0389_),
    .ZN(_0092_));
 MUX2_X1 _2109_ (.A(net75),
    .B(\y[14] ),
    .S(_0385_),
    .Z(_0390_));
 AND2_X1 _2110_ (.A1(_0387_),
    .A2(_0390_),
    .ZN(_0093_));
 MUX2_X1 _2111_ (.A(net76),
    .B(_0758_),
    .S(_0385_),
    .Z(_0391_));
 AND2_X1 _2112_ (.A1(_0387_),
    .A2(_0391_),
    .ZN(_0094_));
 MUX2_X1 _2113_ (.A(net77),
    .B(\y[1] ),
    .S(_0385_),
    .Z(_0392_));
 AND2_X1 _2114_ (.A1(_0387_),
    .A2(_0392_),
    .ZN(_0095_));
 MUX2_X1 _2115_ (.A(net78),
    .B(\y[2] ),
    .S(_0385_),
    .Z(_0393_));
 AND2_X1 _2116_ (.A1(_0387_),
    .A2(_0393_),
    .ZN(_0096_));
 MUX2_X1 _2117_ (.A(net79),
    .B(\y[3] ),
    .S(_0385_),
    .Z(_0394_));
 AND2_X1 _2118_ (.A1(_0387_),
    .A2(_0394_),
    .ZN(_0097_));
 MUX2_X1 _2119_ (.A(net80),
    .B(\y[4] ),
    .S(_0385_),
    .Z(_0395_));
 AND2_X1 _2120_ (.A1(_0387_),
    .A2(_0395_),
    .ZN(_0098_));
 MUX2_X1 _2121_ (.A(net81),
    .B(\y[5] ),
    .S(_0385_),
    .Z(_0396_));
 AND2_X1 _2122_ (.A1(_0387_),
    .A2(_0396_),
    .ZN(_0099_));
 CLKBUF_X3 _2123_ (.A(_0560_),
    .Z(_0397_));
 MUX2_X1 _2124_ (.A(net82),
    .B(\y[6] ),
    .S(_0397_),
    .Z(_0398_));
 AND2_X1 _2125_ (.A1(_0387_),
    .A2(_0398_),
    .ZN(_0100_));
 BUF_X2 _2126_ (.A(_0792_),
    .Z(_0399_));
 MUX2_X1 _2127_ (.A(net83),
    .B(\y[7] ),
    .S(_0397_),
    .Z(_0400_));
 AND2_X1 _2128_ (.A1(_0399_),
    .A2(_0400_),
    .ZN(_0101_));
 MUX2_X1 _2129_ (.A(net84),
    .B(\y[8] ),
    .S(_0397_),
    .Z(_0401_));
 AND2_X1 _2130_ (.A1(_0399_),
    .A2(_0401_),
    .ZN(_0102_));
 MUX2_X1 _2131_ (.A(net85),
    .B(\y[9] ),
    .S(_0397_),
    .Z(_0402_));
 AND2_X1 _2132_ (.A1(_0399_),
    .A2(_0402_),
    .ZN(_0103_));
 NOR2_X1 _2133_ (.A1(_0207_),
    .A2(_1135_),
    .ZN(_0403_));
 MUX2_X1 _2134_ (.A(\z[0] ),
    .B(net37),
    .S(_0337_),
    .Z(_0404_));
 NOR2_X1 _2135_ (.A1(_0136_),
    .A2(_0404_),
    .ZN(_0405_));
 NOR3_X1 _2136_ (.A1(_0347_),
    .A2(_0403_),
    .A3(_0405_),
    .ZN(_0104_));
 INV_X1 _2137_ (.A(_1164_),
    .ZN(_0406_));
 BUF_X1 _2138_ (.A(_1162_),
    .Z(_0407_));
 CLKBUF_X2 _2139_ (.A(_1165_),
    .Z(_0408_));
 AND3_X1 _2140_ (.A1(_0407_),
    .A2(_0408_),
    .A3(_1158_),
    .ZN(_0409_));
 BUF_X1 _2141_ (.A(_1159_),
    .Z(_0410_));
 AND3_X1 _2142_ (.A1(_0410_),
    .A2(_0407_),
    .A3(_0408_),
    .ZN(_0411_));
 BUF_X1 _2143_ (.A(_1152_),
    .Z(_0412_));
 OR2_X1 _2144_ (.A1(_1153_),
    .A2(_0412_),
    .ZN(_0413_));
 BUF_X1 _2145_ (.A(_1156_),
    .Z(_0414_));
 AOI21_X1 _2146_ (.A(_1155_),
    .B1(_0413_),
    .B2(_0414_),
    .ZN(_0415_));
 BUF_X1 _2147_ (.A(_1149_),
    .Z(_0416_));
 NOR3_X1 _2148_ (.A1(_0416_),
    .A2(_0412_),
    .A3(_1155_),
    .ZN(_0417_));
 BUF_X1 _2149_ (.A(_1150_),
    .Z(_0418_));
 INV_X1 _2150_ (.A(_1146_),
    .ZN(_0419_));
 AOI21_X1 _2151_ (.A(_1143_),
    .B1(_1144_),
    .B2(_1108_),
    .ZN(_0420_));
 INV_X1 _2152_ (.A(_1147_),
    .ZN(_0421_));
 OAI21_X2 _2153_ (.A(_0419_),
    .B1(_0420_),
    .B2(_0421_),
    .ZN(_0422_));
 NAND2_X1 _2154_ (.A1(_0418_),
    .A2(_0422_),
    .ZN(_0423_));
 AOI21_X2 _2155_ (.A(_0415_),
    .B1(_0417_),
    .B2(_0423_),
    .ZN(_0424_));
 AOI221_X2 _2156_ (.A(_0409_),
    .B1(_0411_),
    .B2(_0424_),
    .C1(_0408_),
    .C2(_1161_),
    .ZN(_0425_));
 AND2_X1 _2157_ (.A1(_0406_),
    .A2(_0425_),
    .ZN(_0426_));
 XNOR2_X1 _2158_ (.A(_1168_),
    .B(_0426_),
    .ZN(_0427_));
 NOR2_X1 _2159_ (.A1(_0184_),
    .A2(_0427_),
    .ZN(_0428_));
 MUX2_X1 _2160_ (.A(\z[10] ),
    .B(net38),
    .S(_0337_),
    .Z(_0429_));
 NOR2_X1 _2161_ (.A1(_0136_),
    .A2(_0429_),
    .ZN(_0430_));
 NOR3_X1 _2162_ (.A1(_0347_),
    .A2(_0428_),
    .A3(_0430_),
    .ZN(_0105_));
 OR2_X1 _2163_ (.A1(_0408_),
    .A2(_1164_),
    .ZN(_0431_));
 AOI21_X2 _2164_ (.A(_1167_),
    .B1(_0431_),
    .B2(_1168_),
    .ZN(_0432_));
 NOR3_X2 _2165_ (.A1(_1161_),
    .A2(_1164_),
    .A3(_1167_),
    .ZN(_0433_));
 OR3_X1 _2166_ (.A1(_1146_),
    .A2(_0416_),
    .A3(_0412_),
    .ZN(_0434_));
 INV_X1 _2167_ (.A(_1143_),
    .ZN(_0435_));
 AOI21_X1 _2168_ (.A(_1140_),
    .B1(_1141_),
    .B2(_1106_),
    .ZN(_0436_));
 INV_X1 _2169_ (.A(_1144_),
    .ZN(_0437_));
 OAI21_X2 _2170_ (.A(_0435_),
    .B1(_0436_),
    .B2(_0437_),
    .ZN(_0438_));
 AOI21_X2 _2171_ (.A(_0434_),
    .B1(_0438_),
    .B2(_1147_),
    .ZN(_0439_));
 OR2_X1 _2172_ (.A1(_0418_),
    .A2(_0416_),
    .ZN(_0440_));
 AOI21_X2 _2173_ (.A(_0412_),
    .B1(_0440_),
    .B2(_1153_),
    .ZN(_0441_));
 NAND3_X1 _2174_ (.A1(_0414_),
    .A2(_0410_),
    .A3(_0407_),
    .ZN(_0442_));
 NOR3_X2 _2175_ (.A1(_0439_),
    .A2(_0441_),
    .A3(_0442_),
    .ZN(_0443_));
 NAND2_X1 _2176_ (.A1(_0407_),
    .A2(_1158_),
    .ZN(_0444_));
 NAND3_X1 _2177_ (.A1(_0410_),
    .A2(_0407_),
    .A3(_1155_),
    .ZN(_0445_));
 NAND2_X1 _2178_ (.A1(_0444_),
    .A2(_0445_),
    .ZN(_0446_));
 NOR2_X2 _2179_ (.A1(_0443_),
    .A2(_0446_),
    .ZN(_0447_));
 AOI21_X4 _2180_ (.A(_0432_),
    .B1(_0433_),
    .B2(_0447_),
    .ZN(_0448_));
 XOR2_X1 _2181_ (.A(_1171_),
    .B(_0448_),
    .Z(_0449_));
 NOR2_X1 _2182_ (.A1(_0184_),
    .A2(_0449_),
    .ZN(_0450_));
 MUX2_X1 _2183_ (.A(\z[11] ),
    .B(net39),
    .S(_0337_),
    .Z(_0451_));
 NOR2_X1 _2184_ (.A1(_0136_),
    .A2(_0451_),
    .ZN(_0452_));
 NOR3_X1 _2185_ (.A1(_0347_),
    .A2(_0450_),
    .A3(_0452_),
    .ZN(_0106_));
 OR2_X1 _2186_ (.A1(_1168_),
    .A2(_1167_),
    .ZN(_0453_));
 AOI21_X1 _2187_ (.A(_1170_),
    .B1(_0453_),
    .B2(_1171_),
    .ZN(_0454_));
 NOR3_X1 _2188_ (.A1(_1164_),
    .A2(_1167_),
    .A3(_1170_),
    .ZN(_0455_));
 AOI21_X2 _2189_ (.A(_0454_),
    .B1(_0455_),
    .B2(_0425_),
    .ZN(_0456_));
 XOR2_X1 _2190_ (.A(_1174_),
    .B(_0456_),
    .Z(_0457_));
 NOR2_X1 _2191_ (.A1(_0184_),
    .A2(_0457_),
    .ZN(_0458_));
 MUX2_X1 _2192_ (.A(\z[12] ),
    .B(net40),
    .S(_0337_),
    .Z(_0459_));
 NOR2_X1 _2193_ (.A1(_0136_),
    .A2(_0459_),
    .ZN(_0460_));
 NOR3_X1 _2194_ (.A1(_0347_),
    .A2(_0458_),
    .A3(_0460_),
    .ZN(_0107_));
 MUX2_X1 _2195_ (.A(\z[13] ),
    .B(net41),
    .S(_0566_),
    .Z(_0461_));
 NAND3_X1 _2196_ (.A1(_0930_),
    .A2(_0924_),
    .A3(_0461_),
    .ZN(_0462_));
 CLKBUF_X2 _2197_ (.A(_1177_),
    .Z(_0463_));
 AND2_X1 _2198_ (.A1(_1171_),
    .A2(_1174_),
    .ZN(_0464_));
 AOI221_X2 _2199_ (.A(_1173_),
    .B1(_0448_),
    .B2(_0464_),
    .C1(_1170_),
    .C2(_1174_),
    .ZN(_0465_));
 XOR2_X1 _2200_ (.A(_0463_),
    .B(_0465_),
    .Z(_0466_));
 OAI21_X1 _2201_ (.A(_0462_),
    .B1(_0466_),
    .B2(_0791_),
    .ZN(_0108_));
 AND2_X1 _2202_ (.A1(_0567_),
    .A2(_1180_),
    .ZN(_0467_));
 NOR2_X1 _2203_ (.A1(_0923_),
    .A2(_1180_),
    .ZN(_0468_));
 AND2_X1 _2204_ (.A1(_1174_),
    .A2(_0463_),
    .ZN(_0469_));
 AOI221_X2 _2205_ (.A(_1176_),
    .B1(_0456_),
    .B2(_0469_),
    .C1(_1173_),
    .C2(_0463_),
    .ZN(_0470_));
 MUX2_X1 _2206_ (.A(_0467_),
    .B(_0468_),
    .S(_0470_),
    .Z(_0471_));
 MUX2_X1 _2207_ (.A(\z[14] ),
    .B(net42),
    .S(_0927_),
    .Z(_0472_));
 OAI21_X1 _2208_ (.A(_0930_),
    .B1(_0569_),
    .B2(_0472_),
    .ZN(_0473_));
 NOR2_X1 _2209_ (.A1(_0471_),
    .A2(_0473_),
    .ZN(_0109_));
 INV_X1 _2210_ (.A(_1176_),
    .ZN(_0474_));
 AND2_X1 _2211_ (.A1(_0463_),
    .A2(_0464_),
    .ZN(_0475_));
 AOI222_X2 _2212_ (.A1(_0463_),
    .A2(_1173_),
    .B1(_0448_),
    .B2(_0475_),
    .C1(_0469_),
    .C2(_1170_),
    .ZN(_0476_));
 OR4_X1 _2213_ (.A1(_0996_),
    .A2(_0997_),
    .A3(_0606_),
    .A4(_0859_),
    .ZN(_0477_));
 NOR2_X1 _2214_ (.A1(_0613_),
    .A2(_0477_),
    .ZN(_0478_));
 NOR3_X1 _2215_ (.A1(_1179_),
    .A2(_0791_),
    .A3(_0478_),
    .ZN(_0479_));
 NAND3_X1 _2216_ (.A1(_0474_),
    .A2(_0476_),
    .A3(_0479_),
    .ZN(_0480_));
 NOR2_X1 _2217_ (.A1(_1180_),
    .A2(_1179_),
    .ZN(_0481_));
 XOR2_X1 _2218_ (.A(_0481_),
    .B(_0478_),
    .Z(_0482_));
 MUX2_X1 _2219_ (.A(_0653_),
    .B(net43),
    .S(_0565_),
    .Z(_0483_));
 MUX2_X1 _2220_ (.A(_0482_),
    .B(_0483_),
    .S(_0923_),
    .Z(_0484_));
 NAND2_X1 _2221_ (.A1(_0930_),
    .A2(_0484_),
    .ZN(_0485_));
 OAI21_X1 _2222_ (.A(_0481_),
    .B1(_0477_),
    .B2(_0613_),
    .ZN(_0486_));
 AOI21_X1 _2223_ (.A(_0922_),
    .B1(_1179_),
    .B2(_0478_),
    .ZN(_0487_));
 AND4_X1 _2224_ (.A1(_0474_),
    .A2(_0476_),
    .A3(_0486_),
    .A4(_0487_),
    .ZN(_0488_));
 OAI21_X1 _2225_ (.A(_0480_),
    .B1(_0485_),
    .B2(_0488_),
    .ZN(_0110_));
 NAND2_X1 _2226_ (.A1(_0568_),
    .A2(_1109_),
    .ZN(_0489_));
 MUX2_X1 _2227_ (.A(\z[1] ),
    .B(net44),
    .S(_0566_),
    .Z(_0490_));
 OAI21_X1 _2228_ (.A(_0489_),
    .B1(_0490_),
    .B2(_0569_),
    .ZN(_0491_));
 NOR2_X1 _2229_ (.A1(_0564_),
    .A2(_0491_),
    .ZN(_0111_));
 XOR2_X1 _2230_ (.A(_1108_),
    .B(_1144_),
    .Z(_0492_));
 NOR2_X1 _2231_ (.A1(_0184_),
    .A2(_0492_),
    .ZN(_0493_));
 MUX2_X1 _2232_ (.A(\z[2] ),
    .B(net45),
    .S(_0337_),
    .Z(_0494_));
 NOR2_X1 _2233_ (.A1(_0136_),
    .A2(_0494_),
    .ZN(_0495_));
 NOR3_X1 _2234_ (.A1(_0347_),
    .A2(_0493_),
    .A3(_0495_),
    .ZN(_0112_));
 XNOR2_X1 _2235_ (.A(_0421_),
    .B(_0438_),
    .ZN(_0496_));
 NAND2_X1 _2236_ (.A1(_0953_),
    .A2(_0496_),
    .ZN(_0497_));
 MUX2_X1 _2237_ (.A(\z[3] ),
    .B(net46),
    .S(_0566_),
    .Z(_0498_));
 NAND2_X1 _2238_ (.A1(_0924_),
    .A2(_0498_),
    .ZN(_0499_));
 AOI21_X1 _2239_ (.A(_0559_),
    .B1(_0497_),
    .B2(_0499_),
    .ZN(_0113_));
 XOR2_X1 _2240_ (.A(_0418_),
    .B(_0422_),
    .Z(_0500_));
 NOR2_X1 _2241_ (.A1(_0184_),
    .A2(_0500_),
    .ZN(_0501_));
 MUX2_X1 _2242_ (.A(\z[4] ),
    .B(net47),
    .S(_0565_),
    .Z(_0502_));
 NOR2_X1 _2243_ (.A1(_0136_),
    .A2(_0502_),
    .ZN(_0503_));
 NOR3_X1 _2244_ (.A1(_0347_),
    .A2(_0501_),
    .A3(_0503_),
    .ZN(_0114_));
 AOI21_X1 _2245_ (.A(_1146_),
    .B1(_0438_),
    .B2(_1147_),
    .ZN(_0504_));
 INV_X1 _2246_ (.A(_0504_),
    .ZN(_0505_));
 AOI21_X1 _2247_ (.A(_0416_),
    .B1(_0505_),
    .B2(_0418_),
    .ZN(_0506_));
 XNOR2_X1 _2248_ (.A(_1153_),
    .B(_0506_),
    .ZN(_0507_));
 NOR2_X1 _2249_ (.A1(_0184_),
    .A2(_0507_),
    .ZN(_0508_));
 MUX2_X1 _2250_ (.A(\z[5] ),
    .B(net48),
    .S(_0565_),
    .Z(_0509_));
 NOR2_X1 _2251_ (.A1(_0136_),
    .A2(_0509_),
    .ZN(_0510_));
 NOR3_X1 _2252_ (.A1(_0347_),
    .A2(_0508_),
    .A3(_0510_),
    .ZN(_0115_));
 AOI21_X1 _2253_ (.A(_0416_),
    .B1(_0422_),
    .B2(_0418_),
    .ZN(_0511_));
 INV_X1 _2254_ (.A(_0511_),
    .ZN(_0512_));
 AOI21_X1 _2255_ (.A(_0412_),
    .B1(_0512_),
    .B2(_1153_),
    .ZN(_0513_));
 XNOR2_X1 _2256_ (.A(_0414_),
    .B(_0513_),
    .ZN(_0514_));
 NAND2_X1 _2257_ (.A1(_0953_),
    .A2(_0514_),
    .ZN(_0515_));
 MUX2_X1 _2258_ (.A(\z[6] ),
    .B(net49),
    .S(_0566_),
    .Z(_0516_));
 NAND2_X1 _2259_ (.A1(_0924_),
    .A2(_0516_),
    .ZN(_0517_));
 AOI21_X1 _2260_ (.A(_0559_),
    .B1(_0515_),
    .B2(_0517_),
    .ZN(_0116_));
 MUX2_X1 _2261_ (.A(\z[7] ),
    .B(net50),
    .S(_0927_),
    .Z(_0518_));
 OAI21_X1 _2262_ (.A(_0792_),
    .B1(_0926_),
    .B2(_0518_),
    .ZN(_0519_));
 NOR2_X1 _2263_ (.A1(_0439_),
    .A2(_0441_),
    .ZN(_0520_));
 AOI21_X1 _2264_ (.A(_1155_),
    .B1(_0520_),
    .B2(_0414_),
    .ZN(_0521_));
 XOR2_X1 _2265_ (.A(_0410_),
    .B(_0521_),
    .Z(_0522_));
 AOI21_X1 _2266_ (.A(_0519_),
    .B1(_0522_),
    .B2(_0953_),
    .ZN(_0117_));
 MUX2_X1 _2267_ (.A(\z[8] ),
    .B(net51),
    .S(_0927_),
    .Z(_0523_));
 OAI21_X1 _2268_ (.A(_0792_),
    .B1(_0926_),
    .B2(_0523_),
    .ZN(_0524_));
 AOI21_X1 _2269_ (.A(_1158_),
    .B1(_0424_),
    .B2(_0410_),
    .ZN(_0525_));
 XOR2_X1 _2270_ (.A(_0407_),
    .B(_0525_),
    .Z(_0526_));
 AOI21_X1 _2271_ (.A(_0524_),
    .B1(_0526_),
    .B2(_0953_),
    .ZN(_0118_));
 NOR3_X1 _2272_ (.A1(_1161_),
    .A2(_0443_),
    .A3(_0446_),
    .ZN(_0527_));
 XNOR2_X1 _2273_ (.A(_0408_),
    .B(_0527_),
    .ZN(_0528_));
 NOR2_X1 _2274_ (.A1(_0184_),
    .A2(_0528_),
    .ZN(_0529_));
 MUX2_X1 _2275_ (.A(\z[9] ),
    .B(net52),
    .S(_0565_),
    .Z(_0530_));
 NOR2_X1 _2276_ (.A1(_0136_),
    .A2(_0530_),
    .ZN(_0531_));
 NOR3_X1 _2277_ (.A1(_0559_),
    .A2(_0529_),
    .A3(_0531_),
    .ZN(_0119_));
 MUX2_X1 _2278_ (.A(net86),
    .B(\z[0] ),
    .S(_0397_),
    .Z(_0532_));
 AND2_X1 _2279_ (.A1(_0399_),
    .A2(_0532_),
    .ZN(_0120_));
 MUX2_X1 _2280_ (.A(net87),
    .B(\z[10] ),
    .S(_0397_),
    .Z(_0533_));
 AND2_X1 _2281_ (.A1(_0399_),
    .A2(_0533_),
    .ZN(_0121_));
 MUX2_X1 _2282_ (.A(net88),
    .B(\z[11] ),
    .S(_0397_),
    .Z(_0534_));
 AND2_X1 _2283_ (.A1(_0399_),
    .A2(_0534_),
    .ZN(_0122_));
 MUX2_X1 _2284_ (.A(net89),
    .B(\z[12] ),
    .S(_0397_),
    .Z(_0535_));
 AND2_X1 _2285_ (.A1(_0399_),
    .A2(_0535_),
    .ZN(_0123_));
 MUX2_X1 _2286_ (.A(net90),
    .B(\z[13] ),
    .S(_0397_),
    .Z(_0536_));
 AND2_X1 _2287_ (.A1(_0399_),
    .A2(_0536_),
    .ZN(_0124_));
 MUX2_X1 _2288_ (.A(net91),
    .B(\z[14] ),
    .S(_0397_),
    .Z(_0537_));
 AND2_X1 _2289_ (.A1(_0399_),
    .A2(_0537_),
    .ZN(_0125_));
 BUF_X4 _2290_ (.A(_0560_),
    .Z(_0538_));
 MUX2_X1 _2291_ (.A(net92),
    .B(_0673_),
    .S(_0538_),
    .Z(_0539_));
 AND2_X1 _2292_ (.A1(_0399_),
    .A2(_0539_),
    .ZN(_0126_));
 MUX2_X1 _2293_ (.A(net93),
    .B(\z[1] ),
    .S(_0538_),
    .Z(_0540_));
 AND2_X1 _2294_ (.A1(_0793_),
    .A2(_0540_),
    .ZN(_0127_));
 MUX2_X1 _2295_ (.A(net94),
    .B(\z[2] ),
    .S(_0538_),
    .Z(_0541_));
 AND2_X1 _2296_ (.A1(_0793_),
    .A2(_0541_),
    .ZN(_0128_));
 MUX2_X1 _2297_ (.A(net95),
    .B(\z[3] ),
    .S(_0538_),
    .Z(_0542_));
 AND2_X1 _2298_ (.A1(_0793_),
    .A2(_0542_),
    .ZN(_0129_));
 MUX2_X1 _2299_ (.A(net96),
    .B(\z[4] ),
    .S(_0538_),
    .Z(_0543_));
 AND2_X1 _2300_ (.A1(_0793_),
    .A2(_0543_),
    .ZN(_0130_));
 MUX2_X1 _2301_ (.A(net97),
    .B(\z[5] ),
    .S(_0538_),
    .Z(_0544_));
 AND2_X1 _2302_ (.A1(_0793_),
    .A2(_0544_),
    .ZN(_0131_));
 MUX2_X1 _2303_ (.A(net98),
    .B(\z[6] ),
    .S(_0538_),
    .Z(_0545_));
 AND2_X1 _2304_ (.A1(_0793_),
    .A2(_0545_),
    .ZN(_0132_));
 MUX2_X1 _2305_ (.A(net99),
    .B(\z[7] ),
    .S(_0538_),
    .Z(_0546_));
 AND2_X1 _2306_ (.A1(_0793_),
    .A2(_0546_),
    .ZN(_0133_));
 MUX2_X1 _2307_ (.A(net100),
    .B(\z[8] ),
    .S(_0538_),
    .Z(_0547_));
 AND2_X1 _2308_ (.A1(_0793_),
    .A2(_0547_),
    .ZN(_0134_));
 MUX2_X1 _2309_ (.A(net101),
    .B(\z[9] ),
    .S(_0538_),
    .Z(_0548_));
 AND2_X1 _2310_ (.A1(_0793_),
    .A2(_0548_),
    .ZN(_0135_));
 FA_X1 _2311_ (.A(\z[1] ),
    .B(_1106_),
    .CI(_1107_),
    .CO(_1108_),
    .S(_1109_));
 FA_X1 _2312_ (.A(\y[1] ),
    .B(_1110_),
    .CI(_1111_),
    .CO(_1112_),
    .S(_1113_));
 FA_X1 _2313_ (.A(_1114_),
    .B(_1115_),
    .CI(_1116_),
    .CO(_1117_),
    .S(_1118_));
 HA_X1 _2314_ (.A(net111),
    .B(\iteration[1] ),
    .CO(_1119_),
    .S(_1120_));
 HA_X1 _2315_ (.A(_1121_),
    .B(_1122_),
    .CO(_1123_),
    .S(_1124_));
 HA_X1 _2316_ (.A(_1121_),
    .B(_1125_),
    .CO(_1126_),
    .S(_1127_));
 HA_X1 _2317_ (.A(_1121_),
    .B(_1125_),
    .CO(_1128_),
    .S(_1129_));
 HA_X1 _2318_ (.A(_1130_),
    .B(_1122_),
    .CO(_1131_),
    .S(_1132_));
 HA_X1 _2319_ (.A(_1130_),
    .B(_1125_),
    .CO(_1133_),
    .S(_1134_));
 HA_X1 _2320_ (.A(\z[0] ),
    .B(_1007_),
    .CO(_1106_),
    .S(_1135_));
 HA_X1 _2321_ (.A(_1136_),
    .B(_1137_),
    .CO(_1138_),
    .S(_1139_));
 HA_X1 _2322_ (.A(\z[1] ),
    .B(_1107_),
    .CO(_1140_),
    .S(_1141_));
 HA_X1 _2323_ (.A(\z[2] ),
    .B(_1142_),
    .CO(_1143_),
    .S(_1144_));
 HA_X1 _2324_ (.A(\z[3] ),
    .B(_1145_),
    .CO(_1146_),
    .S(_1147_));
 HA_X1 _2325_ (.A(\z[4] ),
    .B(_1148_),
    .CO(_1149_),
    .S(_1150_));
 HA_X1 _2326_ (.A(\z[5] ),
    .B(_1151_),
    .CO(_1152_),
    .S(_1153_));
 HA_X1 _2327_ (.A(\z[6] ),
    .B(_1154_),
    .CO(_1155_),
    .S(_1156_));
 HA_X1 _2328_ (.A(\z[7] ),
    .B(_1157_),
    .CO(_1158_),
    .S(_1159_));
 HA_X1 _2329_ (.A(\z[8] ),
    .B(_1160_),
    .CO(_1161_),
    .S(_1162_));
 HA_X1 _2330_ (.A(\z[9] ),
    .B(_1163_),
    .CO(_1164_),
    .S(_1165_));
 HA_X1 _2331_ (.A(\z[10] ),
    .B(_1166_),
    .CO(_1167_),
    .S(_1168_));
 HA_X1 _2332_ (.A(\z[11] ),
    .B(_1169_),
    .CO(_1170_),
    .S(_1171_));
 HA_X1 _2333_ (.A(\z[12] ),
    .B(_1172_),
    .CO(_1173_),
    .S(_1174_));
 HA_X1 _2334_ (.A(\z[13] ),
    .B(_1175_),
    .CO(_1176_),
    .S(_1177_));
 HA_X1 _2335_ (.A(\z[14] ),
    .B(_1178_),
    .CO(_1179_),
    .S(_1180_));
 HA_X1 _2336_ (.A(_1181_),
    .B(_1182_),
    .CO(_1183_),
    .S(_1184_));
 HA_X1 _2337_ (.A(_1185_),
    .B(_1186_),
    .CO(_1187_),
    .S(_1188_));
 HA_X1 _2338_ (.A(\y[1] ),
    .B(_1111_),
    .CO(_1189_),
    .S(_1190_));
 HA_X1 _2339_ (.A(\y[2] ),
    .B(_1191_),
    .CO(_1192_),
    .S(_1193_));
 HA_X1 _2340_ (.A(_1194_),
    .B(\y[3] ),
    .CO(_1195_),
    .S(_1196_));
 HA_X1 _2341_ (.A(\y[4] ),
    .B(_1197_),
    .CO(_1198_),
    .S(_1199_));
 HA_X1 _2342_ (.A(\y[5] ),
    .B(_1200_),
    .CO(_1201_),
    .S(_1202_));
 HA_X1 _2343_ (.A(_1203_),
    .B(\y[6] ),
    .CO(_1204_),
    .S(_1205_));
 HA_X1 _2344_ (.A(\y[7] ),
    .B(_1206_),
    .CO(_1207_),
    .S(_1208_));
 HA_X1 _2345_ (.A(_1209_),
    .B(\y[8] ),
    .CO(_1210_),
    .S(_1211_));
 HA_X1 _2346_ (.A(\y[9] ),
    .B(_1212_),
    .CO(_1213_),
    .S(_1214_));
 HA_X1 _2347_ (.A(\y[10] ),
    .B(_1215_),
    .CO(_1216_),
    .S(_1217_));
 HA_X1 _2348_ (.A(\y[11] ),
    .B(_1218_),
    .CO(_1219_),
    .S(_1220_));
 HA_X1 _2349_ (.A(\y[12] ),
    .B(_1221_),
    .CO(_1222_),
    .S(_1223_));
 HA_X1 _2350_ (.A(\y[13] ),
    .B(_1224_),
    .CO(_1225_),
    .S(_1226_));
 HA_X1 _2351_ (.A(\y[14] ),
    .B(_1227_),
    .CO(_1228_),
    .S(_1229_));
 HA_X1 _2352_ (.A(\x[0] ),
    .B(net103),
    .CO(_1231_),
    .S(_1232_));
 HA_X1 _2353_ (.A(_1233_),
    .B(_1234_),
    .CO(_1235_),
    .S(_1236_));
 HA_X1 _2354_ (.A(\x[1] ),
    .B(_1237_),
    .CO(_1238_),
    .S(_1239_));
 HA_X1 _2355_ (.A(\x[2] ),
    .B(_1240_),
    .CO(_1241_),
    .S(_1242_));
 HA_X1 _2356_ (.A(_1243_),
    .B(\x[3] ),
    .CO(_1244_),
    .S(_1245_));
 HA_X1 _2357_ (.A(_1246_),
    .B(\x[4] ),
    .CO(_1247_),
    .S(_1248_));
 HA_X1 _2358_ (.A(\x[5] ),
    .B(_1249_),
    .CO(_1250_),
    .S(_1251_));
 HA_X1 _2359_ (.A(_1252_),
    .B(\x[6] ),
    .CO(_1253_),
    .S(_1254_));
 HA_X1 _2360_ (.A(_1255_),
    .B(\x[7] ),
    .CO(_1256_),
    .S(_1257_));
 HA_X1 _2361_ (.A(\x[8] ),
    .B(_1258_),
    .CO(_1259_),
    .S(_1260_));
 HA_X1 _2362_ (.A(\x[9] ),
    .B(_1261_),
    .CO(_1262_),
    .S(_1263_));
 HA_X1 _2363_ (.A(\x[10] ),
    .B(_1264_),
    .CO(_1265_),
    .S(_1266_));
 HA_X1 _2364_ (.A(_1267_),
    .B(\x[11] ),
    .CO(_1268_),
    .S(_1269_));
 HA_X1 _2365_ (.A(\x[12] ),
    .B(_1270_),
    .CO(_1271_),
    .S(_1272_));
 HA_X1 _2366_ (.A(\x[13] ),
    .B(_1273_),
    .CO(_1274_),
    .S(_1275_));
 HA_X1 _2367_ (.A(_1276_),
    .B(\x[14] ),
    .CO(_1277_),
    .S(_1278_));
 DFF_X1 _2368_ (.D(_0027_),
    .CK(clknet_4_7_0_clk),
    .Q(_0994_),
    .QN(_0021_));
 DFF_X1 _2369_ (.D(_0028_),
    .CK(clknet_4_13_0_clk),
    .Q(_0995_),
    .QN(_0022_));
 DFF_X1 _2370_ (.D(_0029_),
    .CK(clknet_4_13_0_clk),
    .Q(_0996_),
    .QN(_0023_));
 DFF_X1 _2371_ (.D(_0030_),
    .CK(clknet_4_12_0_clk),
    .Q(_0997_),
    .QN(_0024_));
 DFF_X1 _2372_ (.D(_0031_),
    .CK(clknet_4_7_0_clk),
    .Q(_1003_),
    .QN(_0017_));
 DFF_X1 _2373_ (.D(_0032_),
    .CK(clknet_4_7_0_clk),
    .Q(_1004_),
    .QN(_0018_));
 DFF_X1 _2374_ (.D(_0033_),
    .CK(clknet_4_7_0_clk),
    .Q(_1005_),
    .QN(_0019_));
 DFF_X1 _2375_ (.D(_0034_),
    .CK(clknet_4_7_0_clk),
    .Q(_1006_),
    .QN(_0020_));
 DFF_X1 _2376_ (.D(_0000_),
    .CK(clknet_4_12_0_clk),
    .Q(_1007_),
    .QN(_1136_));
 DFF_X1 _2377_ (.D(_0001_),
    .CK(clknet_4_6_0_clk),
    .Q(_0998_),
    .QN(_1137_));
 DFF_X1 _2378_ (.D(_0002_),
    .CK(clknet_4_6_0_clk),
    .Q(_0999_),
    .QN(_0013_));
 DFF_X1 _2379_ (.D(_0003_),
    .CK(clknet_4_7_0_clk),
    .Q(_1000_),
    .QN(_0014_));
 DFF_X1 _2380_ (.D(_0004_),
    .CK(clknet_4_7_0_clk),
    .Q(_1001_),
    .QN(_0015_));
 DFF_X1 _2381_ (.D(_0005_),
    .CK(clknet_4_7_0_clk),
    .Q(_1002_),
    .QN(_0016_));
 DFF_X1 \done$_SDFFE_PN0P_  (.D(_0035_),
    .CK(clknet_4_4_0_clk),
    .Q(net53),
    .QN(_1102_));
 DFF_X2 \iteration[0]$_SDFFE_PN0N_  (.D(_0036_),
    .CK(clknet_4_6_0_clk),
    .Q(\iteration[0] ),
    .QN(_0012_));
 DFF_X1 \iteration[1]$_SDFFE_PN0N_  (.D(_0037_),
    .CK(clknet_4_6_0_clk),
    .Q(\iteration[1] ),
    .QN(_0026_));
 DFF_X1 \iteration[2]$_SDFFE_PN0N_  (.D(net144),
    .CK(clknet_4_6_0_clk),
    .Q(\iteration[2] ),
    .QN(_0011_));
 DFF_X2 \iteration[3]$_SDFFE_PN0N_  (.D(_0039_),
    .CK(clknet_4_6_0_clk),
    .Q(\iteration[3] ),
    .QN(_0010_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_0008_),
    .CK(clknet_4_4_0_clk),
    .Q(\state[0] ),
    .QN(_1103_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_0009_),
    .CK(clknet_4_12_0_clk),
    .Q(\state[1] ),
    .QN(_1104_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_0006_),
    .CK(clknet_4_4_0_clk),
    .Q(\state[2] ),
    .QN(_1105_));
 DFF_X1 \state[3]$_DFF_P_  (.D(_0007_),
    .CK(clknet_4_12_0_clk),
    .Q(\state[3] ),
    .QN(_1101_));
 DFF_X2 \x[0]$_SDFFE_PN0N_  (.D(_0040_),
    .CK(clknet_4_3_0_clk),
    .Q(\x[0] ),
    .QN(_1100_));
 DFF_X2 \x[10]$_SDFFE_PN0N_  (.D(_0041_),
    .CK(clknet_4_3_0_clk),
    .Q(\x[10] ),
    .QN(_1099_));
 DFF_X2 \x[11]$_SDFFE_PN0N_  (.D(_0042_),
    .CK(clknet_4_1_0_clk),
    .Q(\x[11] ),
    .QN(_1098_));
 DFF_X2 \x[12]$_SDFFE_PN0N_  (.D(_0043_),
    .CK(clknet_4_1_0_clk),
    .Q(\x[12] ),
    .QN(_1097_));
 DFF_X2 \x[13]$_SDFFE_PN0N_  (.D(_0044_),
    .CK(clknet_4_1_0_clk),
    .Q(\x[13] ),
    .QN(_1096_));
 DFF_X2 \x[14]$_SDFFE_PN0N_  (.D(_0045_),
    .CK(clknet_4_1_0_clk),
    .Q(\x[14] ),
    .QN(_1095_));
 DFF_X1 \x[15]$_SDFFE_PN0N_  (.D(_0046_),
    .CK(clknet_4_6_0_clk),
    .Q(\x[15] ),
    .QN(_1094_));
 DFF_X2 \x[1]$_SDFFE_PN0N_  (.D(_0047_),
    .CK(clknet_4_0_0_clk),
    .Q(\x[1] ),
    .QN(_1114_));
 DFF_X2 \x[2]$_SDFFE_PN0N_  (.D(_0048_),
    .CK(clknet_4_0_0_clk),
    .Q(\x[2] ),
    .QN(_1093_));
 DFF_X2 \x[3]$_SDFFE_PN0N_  (.D(_0049_),
    .CK(clknet_4_0_0_clk),
    .Q(\x[3] ),
    .QN(_1092_));
 DFF_X2 \x[4]$_SDFFE_PN0N_  (.D(_0050_),
    .CK(clknet_4_2_0_clk),
    .Q(\x[4] ),
    .QN(_1091_));
 DFF_X2 \x[5]$_SDFFE_PN0N_  (.D(_0051_),
    .CK(clknet_4_3_0_clk),
    .Q(\x[5] ),
    .QN(_1090_));
 DFF_X2 \x[6]$_SDFFE_PN0N_  (.D(_0052_),
    .CK(clknet_4_2_0_clk),
    .Q(\x[6] ),
    .QN(_1089_));
 DFF_X2 \x[7]$_SDFFE_PN0N_  (.D(_0053_),
    .CK(clknet_4_2_0_clk),
    .Q(\x[7] ),
    .QN(_1088_));
 DFF_X2 \x[8]$_SDFFE_PN0N_  (.D(_0054_),
    .CK(clknet_4_2_0_clk),
    .Q(\x[8] ),
    .QN(_1087_));
 DFF_X2 \x[9]$_SDFFE_PN0N_  (.D(_0055_),
    .CK(clknet_4_8_0_clk),
    .Q(\x[9] ),
    .QN(_1086_));
 DFF_X1 \x_out[0]$_SDFFE_PN0P_  (.D(_0056_),
    .CK(clknet_4_0_0_clk),
    .Q(net54),
    .QN(_1085_));
 DFF_X1 \x_out[10]$_SDFFE_PN0P_  (.D(_0057_),
    .CK(clknet_4_1_0_clk),
    .Q(net55),
    .QN(_1084_));
 DFF_X1 \x_out[11]$_SDFFE_PN0P_  (.D(_0058_),
    .CK(clknet_4_1_0_clk),
    .Q(net56),
    .QN(_1083_));
 DFF_X1 \x_out[12]$_SDFFE_PN0P_  (.D(_0059_),
    .CK(clknet_4_1_0_clk),
    .Q(net57),
    .QN(_1082_));
 DFF_X1 \x_out[13]$_SDFFE_PN0P_  (.D(_0060_),
    .CK(clknet_4_1_0_clk),
    .Q(net58),
    .QN(_1081_));
 DFF_X1 \x_out[14]$_SDFFE_PN0P_  (.D(_0061_),
    .CK(clknet_4_4_0_clk),
    .Q(net59),
    .QN(_1080_));
 DFF_X1 \x_out[15]$_SDFFE_PN0P_  (.D(_0062_),
    .CK(clknet_4_4_0_clk),
    .Q(net60),
    .QN(_1079_));
 DFF_X1 \x_out[1]$_SDFFE_PN0P_  (.D(_0063_),
    .CK(clknet_4_0_0_clk),
    .Q(net61),
    .QN(_1078_));
 DFF_X1 \x_out[2]$_SDFFE_PN0P_  (.D(_0064_),
    .CK(clknet_4_0_0_clk),
    .Q(net62),
    .QN(_1077_));
 DFF_X1 \x_out[3]$_SDFFE_PN0P_  (.D(_0065_),
    .CK(clknet_4_0_0_clk),
    .Q(net63),
    .QN(_1076_));
 DFF_X1 \x_out[4]$_SDFFE_PN0P_  (.D(_0066_),
    .CK(clknet_4_2_0_clk),
    .Q(net64),
    .QN(_1075_));
 DFF_X1 \x_out[5]$_SDFFE_PN0P_  (.D(_0067_),
    .CK(clknet_4_3_0_clk),
    .Q(net65),
    .QN(_1074_));
 DFF_X1 \x_out[6]$_SDFFE_PN0P_  (.D(_0068_),
    .CK(clknet_4_2_0_clk),
    .Q(net66),
    .QN(_1073_));
 DFF_X1 \x_out[7]$_SDFFE_PN0P_  (.D(_0069_),
    .CK(clknet_4_2_0_clk),
    .Q(net67),
    .QN(_1072_));
 DFF_X1 \x_out[8]$_SDFFE_PN0P_  (.D(_0070_),
    .CK(clknet_4_9_0_clk),
    .Q(net68),
    .QN(_1071_));
 DFF_X1 \x_out[9]$_SDFFE_PN0P_  (.D(_0071_),
    .CK(clknet_4_8_0_clk),
    .Q(net69),
    .QN(_1070_));
 DFF_X1 \y[0]$_SDFFE_PN0N_  (.D(_0072_),
    .CK(clknet_4_9_0_clk),
    .Q(\y[0] ),
    .QN(_1181_));
 DFF_X2 \y[10]$_SDFFE_PN0N_  (.D(_0073_),
    .CK(clknet_4_11_0_clk),
    .Q(\y[10] ),
    .QN(_1069_));
 DFF_X2 \y[11]$_SDFFE_PN0N_  (.D(_0074_),
    .CK(clknet_4_11_0_clk),
    .Q(\y[11] ),
    .QN(_1068_));
 DFF_X2 \y[12]$_SDFFE_PN0N_  (.D(_0075_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[12] ),
    .QN(_1067_));
 DFF_X2 \y[13]$_SDFFE_PN0N_  (.D(_0076_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[13] ),
    .QN(_1066_));
 DFF_X2 \y[14]$_SDFFE_PN0N_  (.D(_0077_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[14] ),
    .QN(_1065_));
 DFF_X1 \y[15]$_SDFFE_PN0N_  (.D(_0078_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[15] ),
    .QN(_1064_));
 DFF_X2 \y[1]$_SDFFE_PN0N_  (.D(_0079_),
    .CK(clknet_4_9_0_clk),
    .Q(\y[1] ),
    .QN(_1063_));
 DFF_X2 \y[2]$_SDFFE_PN0N_  (.D(_0080_),
    .CK(clknet_4_10_0_clk),
    .Q(\y[2] ),
    .QN(_1062_));
 DFF_X2 \y[3]$_SDFFE_PN0N_  (.D(_0081_),
    .CK(clknet_4_10_0_clk),
    .Q(\y[3] ),
    .QN(_1061_));
 DFF_X2 \y[4]$_SDFFE_PN0N_  (.D(_0082_),
    .CK(clknet_4_10_0_clk),
    .Q(\y[4] ),
    .QN(_1060_));
 DFF_X2 \y[5]$_SDFFE_PN0N_  (.D(_0083_),
    .CK(clknet_4_10_0_clk),
    .Q(\y[5] ),
    .QN(_1059_));
 DFF_X2 \y[6]$_SDFFE_PN0N_  (.D(_0084_),
    .CK(clknet_4_12_0_clk),
    .Q(\y[6] ),
    .QN(_1058_));
 DFF_X2 \y[7]$_SDFFE_PN0N_  (.D(_0085_),
    .CK(clknet_4_11_0_clk),
    .Q(\y[7] ),
    .QN(_1057_));
 DFF_X2 \y[8]$_SDFFE_PN0N_  (.D(_0086_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[8] ),
    .QN(_1056_));
 DFF_X2 \y[9]$_SDFFE_PN0N_  (.D(_0087_),
    .CK(clknet_4_14_0_clk),
    .Q(\y[9] ),
    .QN(_1055_));
 DFF_X1 \y_out[0]$_SDFFE_PN0P_  (.D(_0088_),
    .CK(clknet_4_8_0_clk),
    .Q(net70),
    .QN(_1054_));
 DFF_X1 \y_out[10]$_SDFFE_PN0P_  (.D(_0089_),
    .CK(clknet_4_8_0_clk),
    .Q(net71),
    .QN(_1053_));
 DFF_X1 \y_out[11]$_SDFFE_PN0P_  (.D(_0090_),
    .CK(clknet_4_9_0_clk),
    .Q(net72),
    .QN(_1052_));
 DFF_X1 \y_out[12]$_SDFFE_PN0P_  (.D(_0091_),
    .CK(clknet_4_11_0_clk),
    .Q(net73),
    .QN(_1051_));
 DFF_X1 \y_out[13]$_SDFFE_PN0P_  (.D(_0092_),
    .CK(clknet_4_14_0_clk),
    .Q(net74),
    .QN(_1050_));
 DFF_X1 \y_out[14]$_SDFFE_PN0P_  (.D(_0093_),
    .CK(clknet_4_14_0_clk),
    .Q(net75),
    .QN(_1049_));
 DFF_X1 \y_out[15]$_SDFFE_PN0P_  (.D(_0094_),
    .CK(clknet_4_11_0_clk),
    .Q(net76),
    .QN(_1048_));
 DFF_X1 \y_out[1]$_SDFFE_PN0P_  (.D(_0095_),
    .CK(clknet_4_9_0_clk),
    .Q(net77),
    .QN(_1047_));
 DFF_X1 \y_out[2]$_SDFFE_PN0P_  (.D(_0096_),
    .CK(clknet_4_10_0_clk),
    .Q(net78),
    .QN(_1046_));
 DFF_X1 \y_out[3]$_SDFFE_PN0P_  (.D(_0097_),
    .CK(clknet_4_10_0_clk),
    .Q(net79),
    .QN(_1045_));
 DFF_X1 \y_out[4]$_SDFFE_PN0P_  (.D(_0098_),
    .CK(clknet_4_10_0_clk),
    .Q(net80),
    .QN(_1044_));
 DFF_X1 \y_out[5]$_SDFFE_PN0P_  (.D(_0099_),
    .CK(clknet_4_11_0_clk),
    .Q(net81),
    .QN(_1043_));
 DFF_X1 \y_out[6]$_SDFFE_PN0P_  (.D(_0100_),
    .CK(clknet_4_14_0_clk),
    .Q(net82),
    .QN(_1042_));
 DFF_X1 \y_out[7]$_SDFFE_PN0P_  (.D(_0101_),
    .CK(clknet_4_15_0_clk),
    .Q(net83),
    .QN(_1041_));
 DFF_X1 \y_out[8]$_SDFFE_PN0P_  (.D(_0102_),
    .CK(clknet_4_15_0_clk),
    .Q(net84),
    .QN(_1040_));
 DFF_X1 \y_out[9]$_SDFFE_PN0P_  (.D(_0103_),
    .CK(clknet_4_14_0_clk),
    .Q(net85),
    .QN(_1039_));
 DFF_X1 \z[0]$_SDFFE_PN0N_  (.D(_0104_),
    .CK(clknet_4_15_0_clk),
    .Q(\z[0] ),
    .QN(_1038_));
 DFF_X1 \z[10]$_SDFFE_PN0N_  (.D(_0105_),
    .CK(clknet_4_13_0_clk),
    .Q(\z[10] ),
    .QN(_1037_));
 DFF_X1 \z[11]$_SDFFE_PN0N_  (.D(_0106_),
    .CK(clknet_4_13_0_clk),
    .Q(\z[11] ),
    .QN(_1036_));
 DFF_X1 \z[12]$_SDFFE_PN0N_  (.D(_0107_),
    .CK(clknet_4_13_0_clk),
    .Q(\z[12] ),
    .QN(_1035_));
 DFF_X1 \z[13]$_SDFFE_PN0N_  (.D(_0108_),
    .CK(clknet_4_13_0_clk),
    .Q(\z[13] ),
    .QN(_1034_));
 DFF_X1 \z[14]$_SDFFE_PN0N_  (.D(_0109_),
    .CK(clknet_4_13_0_clk),
    .Q(\z[14] ),
    .QN(_1033_));
 DFF_X2 \z[15]$_SDFFE_PN0N_  (.D(_0110_),
    .CK(clknet_4_12_0_clk),
    .Q(\z[15] ),
    .QN(_0025_));
 DFF_X2 \z[1]$_SDFFE_PN0N_  (.D(_0111_),
    .CK(clknet_4_4_0_clk),
    .Q(\z[1] ),
    .QN(_1032_));
 DFF_X1 \z[2]$_SDFFE_PN0N_  (.D(_0112_),
    .CK(clknet_4_4_0_clk),
    .Q(\z[2] ),
    .QN(_1031_));
 DFF_X1 \z[3]$_SDFFE_PN0N_  (.D(_0113_),
    .CK(clknet_4_4_0_clk),
    .Q(\z[3] ),
    .QN(_1030_));
 DFF_X1 \z[4]$_SDFFE_PN0N_  (.D(_0114_),
    .CK(clknet_4_5_0_clk),
    .Q(\z[4] ),
    .QN(_1029_));
 DFF_X1 \z[5]$_SDFFE_PN0N_  (.D(_0115_),
    .CK(clknet_4_5_0_clk),
    .Q(\z[5] ),
    .QN(_1028_));
 DFF_X1 \z[6]$_SDFFE_PN0N_  (.D(_0116_),
    .CK(clknet_4_5_0_clk),
    .Q(\z[6] ),
    .QN(_1027_));
 DFF_X1 \z[7]$_SDFFE_PN0N_  (.D(_0117_),
    .CK(clknet_4_5_0_clk),
    .Q(\z[7] ),
    .QN(_1026_));
 DFF_X1 \z[8]$_SDFFE_PN0N_  (.D(_0118_),
    .CK(clknet_4_7_0_clk),
    .Q(\z[8] ),
    .QN(_1025_));
 DFF_X1 \z[9]$_SDFFE_PN0N_  (.D(_0119_),
    .CK(clknet_4_7_0_clk),
    .Q(\z[9] ),
    .QN(_1024_));
 DFF_X1 \z_out[0]$_SDFFE_PN0P_  (.D(_0120_),
    .CK(clknet_4_15_0_clk),
    .Q(net86),
    .QN(_1023_));
 DFF_X1 \z_out[10]$_SDFFE_PN0P_  (.D(_0121_),
    .CK(clknet_4_13_0_clk),
    .Q(net87),
    .QN(_1022_));
 DFF_X1 \z_out[11]$_SDFFE_PN0P_  (.D(_0122_),
    .CK(clknet_4_15_0_clk),
    .Q(net88),
    .QN(_1021_));
 DFF_X1 \z_out[12]$_SDFFE_PN0P_  (.D(_0123_),
    .CK(clknet_4_15_0_clk),
    .Q(net89),
    .QN(_1020_));
 DFF_X1 \z_out[13]$_SDFFE_PN0P_  (.D(_0124_),
    .CK(clknet_4_13_0_clk),
    .Q(net90),
    .QN(_1019_));
 DFF_X1 \z_out[14]$_SDFFE_PN0P_  (.D(_0125_),
    .CK(clknet_4_15_0_clk),
    .Q(net91),
    .QN(_1018_));
 DFF_X1 \z_out[15]$_SDFFE_PN0P_  (.D(_0126_),
    .CK(clknet_4_15_0_clk),
    .Q(net92),
    .QN(_1017_));
 DFF_X1 \z_out[1]$_SDFFE_PN0P_  (.D(_0127_),
    .CK(clknet_4_4_0_clk),
    .Q(net93),
    .QN(_1016_));
 DFF_X1 \z_out[2]$_SDFFE_PN0P_  (.D(_0128_),
    .CK(clknet_4_4_0_clk),
    .Q(net94),
    .QN(_1015_));
 DFF_X1 \z_out[3]$_SDFFE_PN0P_  (.D(_0129_),
    .CK(clknet_4_4_0_clk),
    .Q(net95),
    .QN(_1014_));
 DFF_X1 \z_out[4]$_SDFFE_PN0P_  (.D(_0130_),
    .CK(clknet_4_5_0_clk),
    .Q(net96),
    .QN(_1013_));
 DFF_X1 \z_out[5]$_SDFFE_PN0P_  (.D(_0131_),
    .CK(clknet_4_5_0_clk),
    .Q(net97),
    .QN(_1012_));
 DFF_X1 \z_out[6]$_SDFFE_PN0P_  (.D(_0132_),
    .CK(clknet_4_5_0_clk),
    .Q(net98),
    .QN(_1011_));
 DFF_X1 \z_out[7]$_SDFFE_PN0P_  (.D(_0133_),
    .CK(clknet_4_5_0_clk),
    .Q(net99),
    .QN(_1010_));
 DFF_X1 \z_out[8]$_SDFFE_PN0P_  (.D(_0134_),
    .CK(clknet_4_5_0_clk),
    .Q(net100),
    .QN(_1009_));
 DFF_X1 \z_out[9]$_SDFFE_PN0P_  (.D(_0135_),
    .CK(clknet_4_5_0_clk),
    .Q(net101),
    .QN(_1008_));
 BUF_X4 clone3 (.A(\iteration[0] ),
    .Z(net3));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_85 ();
 BUF_X1 input1 (.A(start),
    .Z(net4));
 BUF_X1 input2 (.A(x_in[0]),
    .Z(net5));
 BUF_X1 input3 (.A(x_in[10]),
    .Z(net6));
 BUF_X1 input4 (.A(x_in[11]),
    .Z(net7));
 BUF_X1 input5 (.A(x_in[12]),
    .Z(net8));
 BUF_X1 input6 (.A(x_in[13]),
    .Z(net9));
 BUF_X1 input7 (.A(x_in[14]),
    .Z(net10));
 BUF_X1 input8 (.A(x_in[15]),
    .Z(net11));
 BUF_X1 input9 (.A(x_in[1]),
    .Z(net12));
 BUF_X1 input10 (.A(x_in[2]),
    .Z(net13));
 BUF_X1 input11 (.A(x_in[3]),
    .Z(net14));
 BUF_X1 input12 (.A(x_in[4]),
    .Z(net15));
 BUF_X1 input13 (.A(x_in[5]),
    .Z(net16));
 BUF_X1 input14 (.A(x_in[6]),
    .Z(net17));
 BUF_X1 input15 (.A(x_in[7]),
    .Z(net18));
 BUF_X1 input16 (.A(x_in[8]),
    .Z(net19));
 BUF_X1 input17 (.A(x_in[9]),
    .Z(net20));
 BUF_X1 input18 (.A(y_in[0]),
    .Z(net21));
 BUF_X1 input19 (.A(y_in[10]),
    .Z(net22));
 BUF_X1 input20 (.A(y_in[11]),
    .Z(net23));
 BUF_X1 input21 (.A(y_in[12]),
    .Z(net24));
 BUF_X1 input22 (.A(y_in[13]),
    .Z(net25));
 BUF_X1 input23 (.A(y_in[14]),
    .Z(net26));
 BUF_X1 input24 (.A(y_in[15]),
    .Z(net27));
 BUF_X1 input25 (.A(y_in[1]),
    .Z(net28));
 BUF_X1 input26 (.A(y_in[2]),
    .Z(net29));
 BUF_X1 input27 (.A(y_in[3]),
    .Z(net30));
 BUF_X1 input28 (.A(y_in[4]),
    .Z(net31));
 BUF_X1 input29 (.A(y_in[5]),
    .Z(net32));
 BUF_X1 input30 (.A(y_in[6]),
    .Z(net33));
 BUF_X1 input31 (.A(y_in[7]),
    .Z(net34));
 BUF_X1 input32 (.A(y_in[8]),
    .Z(net35));
 BUF_X1 input33 (.A(y_in[9]),
    .Z(net36));
 BUF_X1 input34 (.A(z_in[0]),
    .Z(net37));
 BUF_X1 input35 (.A(z_in[10]),
    .Z(net38));
 BUF_X1 input36 (.A(z_in[11]),
    .Z(net39));
 BUF_X1 input37 (.A(z_in[12]),
    .Z(net40));
 BUF_X1 input38 (.A(z_in[13]),
    .Z(net41));
 BUF_X1 input39 (.A(z_in[14]),
    .Z(net42));
 BUF_X1 input40 (.A(z_in[15]),
    .Z(net43));
 BUF_X1 input41 (.A(z_in[1]),
    .Z(net44));
 BUF_X1 input42 (.A(z_in[2]),
    .Z(net45));
 BUF_X1 input43 (.A(z_in[3]),
    .Z(net46));
 BUF_X1 input44 (.A(z_in[4]),
    .Z(net47));
 BUF_X1 input45 (.A(z_in[5]),
    .Z(net48));
 BUF_X1 input46 (.A(z_in[6]),
    .Z(net49));
 BUF_X1 input47 (.A(z_in[7]),
    .Z(net50));
 BUF_X1 input48 (.A(z_in[8]),
    .Z(net51));
 BUF_X1 input49 (.A(z_in[9]),
    .Z(net52));
 BUF_X1 output50 (.A(net53),
    .Z(done));
 BUF_X1 output51 (.A(net54),
    .Z(x_out[0]));
 BUF_X1 output52 (.A(net55),
    .Z(x_out[10]));
 BUF_X1 output53 (.A(net56),
    .Z(x_out[11]));
 BUF_X1 output54 (.A(net57),
    .Z(x_out[12]));
 BUF_X1 output55 (.A(net58),
    .Z(x_out[13]));
 BUF_X1 output56 (.A(net59),
    .Z(x_out[14]));
 BUF_X1 output57 (.A(net60),
    .Z(x_out[15]));
 BUF_X1 output58 (.A(net61),
    .Z(x_out[1]));
 BUF_X1 output59 (.A(net62),
    .Z(x_out[2]));
 BUF_X1 output60 (.A(net63),
    .Z(x_out[3]));
 BUF_X1 output61 (.A(net64),
    .Z(x_out[4]));
 BUF_X1 output62 (.A(net65),
    .Z(x_out[5]));
 BUF_X1 output63 (.A(net66),
    .Z(x_out[6]));
 BUF_X1 output64 (.A(net67),
    .Z(x_out[7]));
 BUF_X1 output65 (.A(net68),
    .Z(x_out[8]));
 BUF_X1 output66 (.A(net69),
    .Z(x_out[9]));
 BUF_X1 output67 (.A(net70),
    .Z(y_out[0]));
 BUF_X1 output68 (.A(net71),
    .Z(y_out[10]));
 BUF_X1 output69 (.A(net72),
    .Z(y_out[11]));
 BUF_X1 output70 (.A(net73),
    .Z(y_out[12]));
 BUF_X1 output71 (.A(net74),
    .Z(y_out[13]));
 BUF_X1 output72 (.A(net75),
    .Z(y_out[14]));
 BUF_X1 output73 (.A(net76),
    .Z(y_out[15]));
 BUF_X1 output74 (.A(net77),
    .Z(y_out[1]));
 BUF_X1 output75 (.A(net78),
    .Z(y_out[2]));
 BUF_X1 output76 (.A(net79),
    .Z(y_out[3]));
 BUF_X1 output77 (.A(net80),
    .Z(y_out[4]));
 BUF_X1 output78 (.A(net81),
    .Z(y_out[5]));
 BUF_X1 output79 (.A(net82),
    .Z(y_out[6]));
 BUF_X1 output80 (.A(net83),
    .Z(y_out[7]));
 BUF_X1 output81 (.A(net84),
    .Z(y_out[8]));
 BUF_X1 output82 (.A(net85),
    .Z(y_out[9]));
 BUF_X1 output83 (.A(net86),
    .Z(z_out[0]));
 BUF_X1 output84 (.A(net87),
    .Z(z_out[10]));
 BUF_X1 output85 (.A(net88),
    .Z(z_out[11]));
 BUF_X1 output86 (.A(net89),
    .Z(z_out[12]));
 BUF_X1 output87 (.A(net90),
    .Z(z_out[13]));
 BUF_X1 output88 (.A(net91),
    .Z(z_out[14]));
 BUF_X1 output89 (.A(net92),
    .Z(z_out[15]));
 BUF_X1 output90 (.A(net93),
    .Z(z_out[1]));
 BUF_X1 output91 (.A(net94),
    .Z(z_out[2]));
 BUF_X1 output92 (.A(net95),
    .Z(z_out[3]));
 BUF_X1 output93 (.A(net96),
    .Z(z_out[4]));
 BUF_X1 output94 (.A(net97),
    .Z(z_out[5]));
 BUF_X1 output95 (.A(net98),
    .Z(z_out[6]));
 BUF_X1 output96 (.A(net99),
    .Z(z_out[7]));
 BUF_X1 output97 (.A(net100),
    .Z(z_out[8]));
 BUF_X1 output98 (.A(net101),
    .Z(z_out[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X2 clkload1 (.A(clknet_4_1_0_clk));
 INV_X2 clkload2 (.A(clknet_4_2_0_clk));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk));
 CLKBUF_X1 clkload4 (.A(clknet_4_5_0_clk));
 INV_X2 clkload5 (.A(clknet_4_6_0_clk));
 CLKBUF_X1 clkload6 (.A(clknet_4_7_0_clk));
 INV_X4 clkload7 (.A(clknet_4_8_0_clk));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_10_0_clk));
 INV_X4 clkload10 (.A(clknet_4_11_0_clk));
 INV_X4 clkload11 (.A(clknet_4_12_0_clk));
 INV_X1 clkload12 (.A(clknet_4_13_0_clk));
 CLKBUF_X1 clkload13 (.A(clknet_4_14_0_clk));
 INV_X2 clkload14 (.A(clknet_4_15_0_clk));
 BUF_X1 rebuffer1 (.A(_0962_),
    .Z(net102));
 BUF_X1 rebuffer2 (.A(_1230_),
    .Z(net103));
 BUF_X1 rebuffer5 (.A(net141),
    .Z(net142));
 BUF_X1 rebuffer4 (.A(_0763_),
    .Z(net105));
 BUF_X1 rebuffer3 (.A(_1245_),
    .Z(net141));
 BUF_X1 rebuffer47 (.A(net150),
    .Z(net151));
 BUF_X4 rebuffer42 (.A(\iteration[0] ),
    .Z(net148));
 BUF_X2 rebuffer46 (.A(_1208_),
    .Z(net150));
 BUF_X2 rebuffer43 (.A(_0283_),
    .Z(net149));
 BUF_X2 rebuffer10 (.A(net112),
    .Z(net111));
 BUF_X1 rebuffer11 (.A(net113),
    .Z(net112));
 BUF_X1 rebuffer12 (.A(net114),
    .Z(net113));
 BUF_X1 rebuffer13 (.A(net115),
    .Z(net114));
 BUF_X1 rebuffer14 (.A(net116),
    .Z(net115));
 BUF_X1 rebuffer15 (.A(net117),
    .Z(net116));
 BUF_X1 rebuffer16 (.A(net118),
    .Z(net117));
 BUF_X1 rebuffer17 (.A(net119),
    .Z(net118));
 BUF_X1 rebuffer18 (.A(net120),
    .Z(net119));
 BUF_X1 rebuffer19 (.A(net121),
    .Z(net120));
 BUF_X1 rebuffer20 (.A(net122),
    .Z(net121));
 BUF_X1 rebuffer21 (.A(net123),
    .Z(net122));
 BUF_X1 rebuffer22 (.A(net124),
    .Z(net123));
 BUF_X1 rebuffer23 (.A(net125),
    .Z(net124));
 BUF_X1 rebuffer24 (.A(net126),
    .Z(net125));
 BUF_X1 rebuffer25 (.A(net127),
    .Z(net126));
 BUF_X1 rebuffer26 (.A(net128),
    .Z(net127));
 BUF_X1 rebuffer27 (.A(net129),
    .Z(net128));
 BUF_X1 rebuffer28 (.A(net130),
    .Z(net129));
 BUF_X1 rebuffer29 (.A(net131),
    .Z(net130));
 BUF_X1 rebuffer30 (.A(net132),
    .Z(net131));
 BUF_X4 rebuffer31 (.A(net133),
    .Z(net132));
 BUF_X4 rebuffer32 (.A(net148),
    .Z(net133));
 BUF_X2 rebuffer33 (.A(_0806_),
    .Z(net134));
 BUF_X1 rebuffer34 (.A(net134),
    .Z(net135));
 BUF_X1 rebuffer35 (.A(_0638_),
    .Z(net136));
 BUF_X1 rebuffer36 (.A(_0623_),
    .Z(net137));
 BUF_X4 rebuffer37 (.A(_0689_),
    .Z(net138));
 BUF_X8 rebuffer38 (.A(_0577_),
    .Z(net139));
 BUF_X1 rebuffer44 (.A(_1196_),
    .Z(net145));
 BUF_X1 rebuffer45 (.A(_1199_),
    .Z(net146));
 BUF_X2 max_cap1 (.A(_0699_),
    .Z(net140));
 BUF_X2 rebuffer39 (.A(_0676_),
    .Z(net143));
 NOR2_X2 clone40 (.A1(net147),
    .A2(_0558_),
    .ZN(net144));
 BUF_X2 rebuffer41 (.A(_0594_),
    .Z(net147));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_41 ();
 FILLCELL_X1 FILLER_0_45 ();
 FILLCELL_X4 FILLER_0_72 ();
 FILLCELL_X1 FILLER_0_76 ();
 FILLCELL_X8 FILLER_0_80 ();
 FILLCELL_X2 FILLER_0_88 ();
 FILLCELL_X1 FILLER_0_90 ();
 FILLCELL_X1 FILLER_0_98 ();
 FILLCELL_X2 FILLER_0_102 ();
 FILLCELL_X1 FILLER_0_111 ();
 FILLCELL_X2 FILLER_0_115 ();
 FILLCELL_X8 FILLER_0_127 ();
 FILLCELL_X4 FILLER_0_138 ();
 FILLCELL_X2 FILLER_0_142 ();
 FILLCELL_X1 FILLER_0_144 ();
 FILLCELL_X8 FILLER_0_148 ();
 FILLCELL_X2 FILLER_0_166 ();
 FILLCELL_X8 FILLER_0_178 ();
 FILLCELL_X4 FILLER_0_199 ();
 FILLCELL_X2 FILLER_0_203 ();
 FILLCELL_X1 FILLER_0_205 ();
 FILLCELL_X8 FILLER_0_212 ();
 FILLCELL_X8 FILLER_0_230 ();
 FILLCELL_X1 FILLER_0_238 ();
 FILLCELL_X2 FILLER_0_242 ();
 FILLCELL_X1 FILLER_0_244 ();
 FILLCELL_X8 FILLER_0_248 ();
 FILLCELL_X1 FILLER_0_256 ();
 FILLCELL_X2 FILLER_0_264 ();
 FILLCELL_X4 FILLER_0_269 ();
 FILLCELL_X2 FILLER_0_287 ();
 FILLCELL_X32 FILLER_0_292 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X1 FILLER_1_33 ();
 FILLCELL_X1 FILLER_1_55 ();
 FILLCELL_X8 FILLER_1_67 ();
 FILLCELL_X4 FILLER_1_82 ();
 FILLCELL_X2 FILLER_1_86 ();
 FILLCELL_X1 FILLER_1_88 ();
 FILLCELL_X2 FILLER_1_114 ();
 FILLCELL_X1 FILLER_1_116 ();
 FILLCELL_X4 FILLER_1_150 ();
 FILLCELL_X8 FILLER_1_211 ();
 FILLCELL_X4 FILLER_1_219 ();
 FILLCELL_X1 FILLER_1_223 ();
 FILLCELL_X1 FILLER_1_273 ();
 FILLCELL_X32 FILLER_1_291 ();
 FILLCELL_X1 FILLER_1_323 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_41 ();
 FILLCELL_X2 FILLER_2_45 ();
 FILLCELL_X16 FILLER_2_54 ();
 FILLCELL_X4 FILLER_2_70 ();
 FILLCELL_X1 FILLER_2_74 ();
 FILLCELL_X8 FILLER_2_78 ();
 FILLCELL_X2 FILLER_2_86 ();
 FILLCELL_X1 FILLER_2_88 ();
 FILLCELL_X16 FILLER_2_106 ();
 FILLCELL_X16 FILLER_2_125 ();
 FILLCELL_X2 FILLER_2_151 ();
 FILLCELL_X1 FILLER_2_153 ();
 FILLCELL_X4 FILLER_2_171 ();
 FILLCELL_X1 FILLER_2_175 ();
 FILLCELL_X8 FILLER_2_187 ();
 FILLCELL_X2 FILLER_2_195 ();
 FILLCELL_X1 FILLER_2_197 ();
 FILLCELL_X16 FILLER_2_219 ();
 FILLCELL_X1 FILLER_2_235 ();
 FILLCELL_X16 FILLER_2_243 ();
 FILLCELL_X4 FILLER_2_259 ();
 FILLCELL_X2 FILLER_2_267 ();
 FILLCELL_X32 FILLER_2_276 ();
 FILLCELL_X16 FILLER_2_308 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X4 FILLER_3_33 ();
 FILLCELL_X2 FILLER_3_37 ();
 FILLCELL_X1 FILLER_3_39 ();
 FILLCELL_X4 FILLER_3_43 ();
 FILLCELL_X2 FILLER_3_47 ();
 FILLCELL_X8 FILLER_3_56 ();
 FILLCELL_X4 FILLER_3_64 ();
 FILLCELL_X8 FILLER_3_96 ();
 FILLCELL_X2 FILLER_3_104 ();
 FILLCELL_X1 FILLER_3_106 ();
 FILLCELL_X1 FILLER_3_113 ();
 FILLCELL_X4 FILLER_3_117 ();
 FILLCELL_X1 FILLER_3_125 ();
 FILLCELL_X1 FILLER_3_149 ();
 FILLCELL_X4 FILLER_3_169 ();
 FILLCELL_X1 FILLER_3_173 ();
 FILLCELL_X8 FILLER_3_191 ();
 FILLCELL_X2 FILLER_3_199 ();
 FILLCELL_X1 FILLER_3_201 ();
 FILLCELL_X8 FILLER_3_209 ();
 FILLCELL_X4 FILLER_3_217 ();
 FILLCELL_X4 FILLER_3_228 ();
 FILLCELL_X2 FILLER_3_232 ();
 FILLCELL_X1 FILLER_3_234 ();
 FILLCELL_X8 FILLER_3_261 ();
 FILLCELL_X2 FILLER_3_269 ();
 FILLCELL_X1 FILLER_3_271 ();
 FILLCELL_X32 FILLER_3_275 ();
 FILLCELL_X16 FILLER_3_307 ();
 FILLCELL_X1 FILLER_3_323 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X2 FILLER_4_33 ();
 FILLCELL_X1 FILLER_4_35 ();
 FILLCELL_X4 FILLER_4_59 ();
 FILLCELL_X1 FILLER_4_63 ();
 FILLCELL_X4 FILLER_4_70 ();
 FILLCELL_X2 FILLER_4_74 ();
 FILLCELL_X1 FILLER_4_82 ();
 FILLCELL_X1 FILLER_4_90 ();
 FILLCELL_X1 FILLER_4_95 ();
 FILLCELL_X32 FILLER_4_121 ();
 FILLCELL_X4 FILLER_4_153 ();
 FILLCELL_X1 FILLER_4_157 ();
 FILLCELL_X16 FILLER_4_165 ();
 FILLCELL_X8 FILLER_4_181 ();
 FILLCELL_X2 FILLER_4_189 ();
 FILLCELL_X8 FILLER_4_194 ();
 FILLCELL_X4 FILLER_4_202 ();
 FILLCELL_X4 FILLER_4_210 ();
 FILLCELL_X1 FILLER_4_214 ();
 FILLCELL_X2 FILLER_4_236 ();
 FILLCELL_X1 FILLER_4_248 ();
 FILLCELL_X16 FILLER_4_251 ();
 FILLCELL_X4 FILLER_4_267 ();
 FILLCELL_X1 FILLER_4_271 ();
 FILLCELL_X8 FILLER_4_291 ();
 FILLCELL_X4 FILLER_4_299 ();
 FILLCELL_X1 FILLER_4_320 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_17 ();
 FILLCELL_X2 FILLER_5_25 ();
 FILLCELL_X1 FILLER_5_27 ();
 FILLCELL_X16 FILLER_5_31 ();
 FILLCELL_X4 FILLER_5_47 ();
 FILLCELL_X2 FILLER_5_53 ();
 FILLCELL_X1 FILLER_5_55 ();
 FILLCELL_X4 FILLER_5_60 ();
 FILLCELL_X2 FILLER_5_64 ();
 FILLCELL_X1 FILLER_5_70 ();
 FILLCELL_X2 FILLER_5_115 ();
 FILLCELL_X2 FILLER_5_125 ();
 FILLCELL_X1 FILLER_5_136 ();
 FILLCELL_X16 FILLER_5_141 ();
 FILLCELL_X4 FILLER_5_170 ();
 FILLCELL_X2 FILLER_5_174 ();
 FILLCELL_X4 FILLER_5_183 ();
 FILLCELL_X2 FILLER_5_187 ();
 FILLCELL_X4 FILLER_5_206 ();
 FILLCELL_X2 FILLER_5_223 ();
 FILLCELL_X1 FILLER_5_225 ();
 FILLCELL_X4 FILLER_5_245 ();
 FILLCELL_X1 FILLER_5_249 ();
 FILLCELL_X1 FILLER_5_269 ();
 FILLCELL_X1 FILLER_5_277 ();
 FILLCELL_X4 FILLER_5_281 ();
 FILLCELL_X4 FILLER_5_292 ();
 FILLCELL_X1 FILLER_5_296 ();
 FILLCELL_X8 FILLER_5_311 ();
 FILLCELL_X4 FILLER_5_319 ();
 FILLCELL_X1 FILLER_5_323 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_9 ();
 FILLCELL_X8 FILLER_6_13 ();
 FILLCELL_X1 FILLER_6_28 ();
 FILLCELL_X1 FILLER_6_33 ();
 FILLCELL_X1 FILLER_6_37 ();
 FILLCELL_X1 FILLER_6_44 ();
 FILLCELL_X2 FILLER_6_61 ();
 FILLCELL_X1 FILLER_6_63 ();
 FILLCELL_X2 FILLER_6_74 ();
 FILLCELL_X1 FILLER_6_95 ();
 FILLCELL_X16 FILLER_6_138 ();
 FILLCELL_X4 FILLER_6_154 ();
 FILLCELL_X1 FILLER_6_158 ();
 FILLCELL_X16 FILLER_6_194 ();
 FILLCELL_X8 FILLER_6_210 ();
 FILLCELL_X1 FILLER_6_220 ();
 FILLCELL_X32 FILLER_6_224 ();
 FILLCELL_X2 FILLER_6_256 ();
 FILLCELL_X1 FILLER_6_258 ();
 FILLCELL_X1 FILLER_6_263 ();
 FILLCELL_X1 FILLER_6_268 ();
 FILLCELL_X1 FILLER_6_278 ();
 FILLCELL_X16 FILLER_6_302 ();
 FILLCELL_X4 FILLER_6_318 ();
 FILLCELL_X2 FILLER_6_322 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_36 ();
 FILLCELL_X2 FILLER_7_40 ();
 FILLCELL_X4 FILLER_7_76 ();
 FILLCELL_X1 FILLER_7_80 ();
 FILLCELL_X2 FILLER_7_88 ();
 FILLCELL_X8 FILLER_7_96 ();
 FILLCELL_X4 FILLER_7_104 ();
 FILLCELL_X2 FILLER_7_108 ();
 FILLCELL_X1 FILLER_7_110 ();
 FILLCELL_X4 FILLER_7_113 ();
 FILLCELL_X2 FILLER_7_138 ();
 FILLCELL_X4 FILLER_7_153 ();
 FILLCELL_X2 FILLER_7_157 ();
 FILLCELL_X1 FILLER_7_180 ();
 FILLCELL_X4 FILLER_7_188 ();
 FILLCELL_X1 FILLER_7_192 ();
 FILLCELL_X16 FILLER_7_200 ();
 FILLCELL_X8 FILLER_7_216 ();
 FILLCELL_X2 FILLER_7_224 ();
 FILLCELL_X4 FILLER_7_236 ();
 FILLCELL_X2 FILLER_7_240 ();
 FILLCELL_X2 FILLER_7_244 ();
 FILLCELL_X1 FILLER_7_246 ();
 FILLCELL_X1 FILLER_7_257 ();
 FILLCELL_X1 FILLER_7_261 ();
 FILLCELL_X1 FILLER_7_266 ();
 FILLCELL_X1 FILLER_7_276 ();
 FILLCELL_X1 FILLER_7_279 ();
 FILLCELL_X8 FILLER_7_283 ();
 FILLCELL_X4 FILLER_7_291 ();
 FILLCELL_X1 FILLER_7_295 ();
 FILLCELL_X8 FILLER_7_315 ();
 FILLCELL_X1 FILLER_7_323 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_27 ();
 FILLCELL_X8 FILLER_8_43 ();
 FILLCELL_X4 FILLER_8_51 ();
 FILLCELL_X16 FILLER_8_62 ();
 FILLCELL_X2 FILLER_8_78 ();
 FILLCELL_X1 FILLER_8_80 ();
 FILLCELL_X16 FILLER_8_84 ();
 FILLCELL_X4 FILLER_8_100 ();
 FILLCELL_X2 FILLER_8_104 ();
 FILLCELL_X32 FILLER_8_115 ();
 FILLCELL_X4 FILLER_8_147 ();
 FILLCELL_X4 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_165 ();
 FILLCELL_X8 FILLER_8_176 ();
 FILLCELL_X2 FILLER_8_184 ();
 FILLCELL_X4 FILLER_8_189 ();
 FILLCELL_X2 FILLER_8_193 ();
 FILLCELL_X8 FILLER_8_209 ();
 FILLCELL_X4 FILLER_8_217 ();
 FILLCELL_X2 FILLER_8_221 ();
 FILLCELL_X1 FILLER_8_223 ();
 FILLCELL_X1 FILLER_8_255 ();
 FILLCELL_X4 FILLER_8_301 ();
 FILLCELL_X2 FILLER_8_305 ();
 FILLCELL_X1 FILLER_8_307 ();
 FILLCELL_X8 FILLER_8_315 ();
 FILLCELL_X1 FILLER_8_323 ();
 FILLCELL_X2 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_6 ();
 FILLCELL_X2 FILLER_9_14 ();
 FILLCELL_X1 FILLER_9_16 ();
 FILLCELL_X2 FILLER_9_20 ();
 FILLCELL_X1 FILLER_9_22 ();
 FILLCELL_X2 FILLER_9_30 ();
 FILLCELL_X1 FILLER_9_32 ();
 FILLCELL_X2 FILLER_9_36 ();
 FILLCELL_X1 FILLER_9_38 ();
 FILLCELL_X8 FILLER_9_43 ();
 FILLCELL_X2 FILLER_9_51 ();
 FILLCELL_X1 FILLER_9_53 ();
 FILLCELL_X4 FILLER_9_66 ();
 FILLCELL_X1 FILLER_9_70 ();
 FILLCELL_X1 FILLER_9_101 ();
 FILLCELL_X4 FILLER_9_131 ();
 FILLCELL_X2 FILLER_9_135 ();
 FILLCELL_X1 FILLER_9_159 ();
 FILLCELL_X2 FILLER_9_167 ();
 FILLCELL_X1 FILLER_9_179 ();
 FILLCELL_X4 FILLER_9_194 ();
 FILLCELL_X8 FILLER_9_205 ();
 FILLCELL_X2 FILLER_9_213 ();
 FILLCELL_X1 FILLER_9_222 ();
 FILLCELL_X2 FILLER_9_247 ();
 FILLCELL_X1 FILLER_9_249 ();
 FILLCELL_X2 FILLER_9_256 ();
 FILLCELL_X2 FILLER_9_268 ();
 FILLCELL_X4 FILLER_9_293 ();
 FILLCELL_X1 FILLER_9_297 ();
 FILLCELL_X2 FILLER_9_312 ();
 FILLCELL_X2 FILLER_9_317 ();
 FILLCELL_X1 FILLER_9_319 ();
 FILLCELL_X1 FILLER_9_323 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_17 ();
 FILLCELL_X2 FILLER_10_25 ();
 FILLCELL_X4 FILLER_10_70 ();
 FILLCELL_X1 FILLER_10_74 ();
 FILLCELL_X8 FILLER_10_78 ();
 FILLCELL_X1 FILLER_10_102 ();
 FILLCELL_X2 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_148 ();
 FILLCELL_X2 FILLER_10_158 ();
 FILLCELL_X1 FILLER_10_160 ();
 FILLCELL_X1 FILLER_10_186 ();
 FILLCELL_X2 FILLER_10_190 ();
 FILLCELL_X1 FILLER_10_199 ();
 FILLCELL_X4 FILLER_10_207 ();
 FILLCELL_X2 FILLER_10_256 ();
 FILLCELL_X1 FILLER_10_258 ();
 FILLCELL_X1 FILLER_10_292 ();
 FILLCELL_X1 FILLER_10_303 ();
 FILLCELL_X2 FILLER_10_321 ();
 FILLCELL_X1 FILLER_10_323 ();
 FILLCELL_X4 FILLER_11_29 ();
 FILLCELL_X2 FILLER_11_33 ();
 FILLCELL_X16 FILLER_11_40 ();
 FILLCELL_X8 FILLER_11_58 ();
 FILLCELL_X1 FILLER_11_66 ();
 FILLCELL_X1 FILLER_11_77 ();
 FILLCELL_X8 FILLER_11_85 ();
 FILLCELL_X1 FILLER_11_93 ();
 FILLCELL_X1 FILLER_11_106 ();
 FILLCELL_X2 FILLER_11_116 ();
 FILLCELL_X1 FILLER_11_118 ();
 FILLCELL_X2 FILLER_11_138 ();
 FILLCELL_X1 FILLER_11_140 ();
 FILLCELL_X1 FILLER_11_148 ();
 FILLCELL_X4 FILLER_11_162 ();
 FILLCELL_X2 FILLER_11_166 ();
 FILLCELL_X1 FILLER_11_177 ();
 FILLCELL_X8 FILLER_11_195 ();
 FILLCELL_X2 FILLER_11_203 ();
 FILLCELL_X1 FILLER_11_212 ();
 FILLCELL_X1 FILLER_11_220 ();
 FILLCELL_X1 FILLER_11_234 ();
 FILLCELL_X2 FILLER_11_260 ();
 FILLCELL_X1 FILLER_11_262 ();
 FILLCELL_X2 FILLER_11_272 ();
 FILLCELL_X1 FILLER_11_278 ();
 FILLCELL_X2 FILLER_11_292 ();
 FILLCELL_X1 FILLER_11_320 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_5 ();
 FILLCELL_X2 FILLER_12_9 ();
 FILLCELL_X4 FILLER_12_22 ();
 FILLCELL_X1 FILLER_12_26 ();
 FILLCELL_X4 FILLER_12_59 ();
 FILLCELL_X2 FILLER_12_63 ();
 FILLCELL_X1 FILLER_12_65 ();
 FILLCELL_X4 FILLER_12_79 ();
 FILLCELL_X2 FILLER_12_83 ();
 FILLCELL_X1 FILLER_12_85 ();
 FILLCELL_X1 FILLER_12_101 ();
 FILLCELL_X1 FILLER_12_116 ();
 FILLCELL_X2 FILLER_12_121 ();
 FILLCELL_X4 FILLER_12_137 ();
 FILLCELL_X1 FILLER_12_146 ();
 FILLCELL_X4 FILLER_12_153 ();
 FILLCELL_X2 FILLER_12_157 ();
 FILLCELL_X2 FILLER_12_166 ();
 FILLCELL_X1 FILLER_12_168 ();
 FILLCELL_X2 FILLER_12_176 ();
 FILLCELL_X4 FILLER_12_233 ();
 FILLCELL_X4 FILLER_12_256 ();
 FILLCELL_X2 FILLER_12_260 ();
 FILLCELL_X1 FILLER_12_262 ();
 FILLCELL_X1 FILLER_12_275 ();
 FILLCELL_X16 FILLER_12_289 ();
 FILLCELL_X4 FILLER_12_305 ();
 FILLCELL_X1 FILLER_12_309 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_3 ();
 FILLCELL_X4 FILLER_13_24 ();
 FILLCELL_X1 FILLER_13_28 ();
 FILLCELL_X4 FILLER_13_36 ();
 FILLCELL_X1 FILLER_13_63 ();
 FILLCELL_X4 FILLER_13_68 ();
 FILLCELL_X2 FILLER_13_72 ();
 FILLCELL_X8 FILLER_13_91 ();
 FILLCELL_X4 FILLER_13_99 ();
 FILLCELL_X2 FILLER_13_103 ();
 FILLCELL_X1 FILLER_13_105 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_134 ();
 FILLCELL_X1 FILLER_13_146 ();
 FILLCELL_X8 FILLER_13_159 ();
 FILLCELL_X4 FILLER_13_174 ();
 FILLCELL_X1 FILLER_13_178 ();
 FILLCELL_X1 FILLER_13_186 ();
 FILLCELL_X2 FILLER_13_194 ();
 FILLCELL_X2 FILLER_13_205 ();
 FILLCELL_X2 FILLER_13_216 ();
 FILLCELL_X2 FILLER_13_225 ();
 FILLCELL_X1 FILLER_13_227 ();
 FILLCELL_X4 FILLER_13_269 ();
 FILLCELL_X1 FILLER_13_273 ();
 FILLCELL_X1 FILLER_13_285 ();
 FILLCELL_X2 FILLER_13_297 ();
 FILLCELL_X2 FILLER_13_305 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_5 ();
 FILLCELL_X8 FILLER_14_9 ();
 FILLCELL_X4 FILLER_14_17 ();
 FILLCELL_X2 FILLER_14_21 ();
 FILLCELL_X4 FILLER_14_33 ();
 FILLCELL_X1 FILLER_14_37 ();
 FILLCELL_X8 FILLER_14_50 ();
 FILLCELL_X8 FILLER_14_68 ();
 FILLCELL_X1 FILLER_14_76 ();
 FILLCELL_X16 FILLER_14_88 ();
 FILLCELL_X4 FILLER_14_104 ();
 FILLCELL_X2 FILLER_14_108 ();
 FILLCELL_X8 FILLER_14_117 ();
 FILLCELL_X4 FILLER_14_125 ();
 FILLCELL_X2 FILLER_14_129 ();
 FILLCELL_X2 FILLER_14_140 ();
 FILLCELL_X4 FILLER_14_151 ();
 FILLCELL_X1 FILLER_14_155 ();
 FILLCELL_X2 FILLER_14_163 ();
 FILLCELL_X2 FILLER_14_172 ();
 FILLCELL_X8 FILLER_14_181 ();
 FILLCELL_X1 FILLER_14_189 ();
 FILLCELL_X2 FILLER_14_205 ();
 FILLCELL_X1 FILLER_14_207 ();
 FILLCELL_X2 FILLER_14_217 ();
 FILLCELL_X1 FILLER_14_219 ();
 FILLCELL_X1 FILLER_14_234 ();
 FILLCELL_X8 FILLER_14_251 ();
 FILLCELL_X4 FILLER_14_259 ();
 FILLCELL_X2 FILLER_14_263 ();
 FILLCELL_X1 FILLER_14_265 ();
 FILLCELL_X2 FILLER_14_279 ();
 FILLCELL_X1 FILLER_14_281 ();
 FILLCELL_X8 FILLER_14_313 ();
 FILLCELL_X2 FILLER_14_321 ();
 FILLCELL_X1 FILLER_14_323 ();
 FILLCELL_X4 FILLER_15_4 ();
 FILLCELL_X1 FILLER_15_8 ();
 FILLCELL_X1 FILLER_15_13 ();
 FILLCELL_X4 FILLER_15_24 ();
 FILLCELL_X2 FILLER_15_28 ();
 FILLCELL_X2 FILLER_15_60 ();
 FILLCELL_X1 FILLER_15_62 ();
 FILLCELL_X4 FILLER_15_69 ();
 FILLCELL_X16 FILLER_15_87 ();
 FILLCELL_X2 FILLER_15_103 ();
 FILLCELL_X8 FILLER_15_107 ();
 FILLCELL_X4 FILLER_15_115 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X1 FILLER_15_162 ();
 FILLCELL_X4 FILLER_15_170 ();
 FILLCELL_X2 FILLER_15_174 ();
 FILLCELL_X1 FILLER_15_176 ();
 FILLCELL_X1 FILLER_15_198 ();
 FILLCELL_X4 FILLER_15_202 ();
 FILLCELL_X1 FILLER_15_206 ();
 FILLCELL_X4 FILLER_15_248 ();
 FILLCELL_X1 FILLER_15_252 ();
 FILLCELL_X2 FILLER_15_275 ();
 FILLCELL_X8 FILLER_15_288 ();
 FILLCELL_X4 FILLER_15_319 ();
 FILLCELL_X1 FILLER_15_323 ();
 FILLCELL_X2 FILLER_16_18 ();
 FILLCELL_X1 FILLER_16_20 ();
 FILLCELL_X2 FILLER_16_24 ();
 FILLCELL_X1 FILLER_16_26 ();
 FILLCELL_X2 FILLER_16_34 ();
 FILLCELL_X2 FILLER_16_62 ();
 FILLCELL_X1 FILLER_16_64 ();
 FILLCELL_X8 FILLER_16_77 ();
 FILLCELL_X4 FILLER_16_85 ();
 FILLCELL_X2 FILLER_16_89 ();
 FILLCELL_X1 FILLER_16_117 ();
 FILLCELL_X4 FILLER_16_125 ();
 FILLCELL_X4 FILLER_16_163 ();
 FILLCELL_X2 FILLER_16_167 ();
 FILLCELL_X2 FILLER_16_185 ();
 FILLCELL_X2 FILLER_16_191 ();
 FILLCELL_X2 FILLER_16_239 ();
 FILLCELL_X2 FILLER_16_253 ();
 FILLCELL_X1 FILLER_16_255 ();
 FILLCELL_X2 FILLER_16_270 ();
 FILLCELL_X1 FILLER_16_272 ();
 FILLCELL_X2 FILLER_16_281 ();
 FILLCELL_X1 FILLER_16_299 ();
 FILLCELL_X4 FILLER_16_318 ();
 FILLCELL_X2 FILLER_16_322 ();
 FILLCELL_X1 FILLER_17_25 ();
 FILLCELL_X4 FILLER_17_30 ();
 FILLCELL_X8 FILLER_17_53 ();
 FILLCELL_X2 FILLER_17_61 ();
 FILLCELL_X16 FILLER_17_81 ();
 FILLCELL_X1 FILLER_17_97 ();
 FILLCELL_X1 FILLER_17_106 ();
 FILLCELL_X1 FILLER_17_131 ();
 FILLCELL_X2 FILLER_17_144 ();
 FILLCELL_X1 FILLER_17_146 ();
 FILLCELL_X2 FILLER_17_184 ();
 FILLCELL_X1 FILLER_17_186 ();
 FILLCELL_X1 FILLER_17_205 ();
 FILLCELL_X8 FILLER_17_250 ();
 FILLCELL_X2 FILLER_17_258 ();
 FILLCELL_X2 FILLER_17_274 ();
 FILLCELL_X1 FILLER_17_276 ();
 FILLCELL_X2 FILLER_17_292 ();
 FILLCELL_X4 FILLER_17_317 ();
 FILLCELL_X2 FILLER_17_321 ();
 FILLCELL_X1 FILLER_17_323 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_9 ();
 FILLCELL_X1 FILLER_18_11 ();
 FILLCELL_X1 FILLER_18_15 ();
 FILLCELL_X2 FILLER_18_20 ();
 FILLCELL_X1 FILLER_18_22 ();
 FILLCELL_X4 FILLER_18_30 ();
 FILLCELL_X1 FILLER_18_34 ();
 FILLCELL_X2 FILLER_18_54 ();
 FILLCELL_X1 FILLER_18_61 ();
 FILLCELL_X4 FILLER_18_71 ();
 FILLCELL_X4 FILLER_18_94 ();
 FILLCELL_X8 FILLER_18_116 ();
 FILLCELL_X4 FILLER_18_124 ();
 FILLCELL_X2 FILLER_18_128 ();
 FILLCELL_X1 FILLER_18_130 ();
 FILLCELL_X2 FILLER_18_138 ();
 FILLCELL_X4 FILLER_18_158 ();
 FILLCELL_X4 FILLER_18_169 ();
 FILLCELL_X1 FILLER_18_173 ();
 FILLCELL_X8 FILLER_18_181 ();
 FILLCELL_X1 FILLER_18_189 ();
 FILLCELL_X2 FILLER_18_194 ();
 FILLCELL_X2 FILLER_18_224 ();
 FILLCELL_X1 FILLER_18_231 ();
 FILLCELL_X4 FILLER_18_248 ();
 FILLCELL_X1 FILLER_18_252 ();
 FILLCELL_X16 FILLER_18_266 ();
 FILLCELL_X4 FILLER_18_301 ();
 FILLCELL_X2 FILLER_18_305 ();
 FILLCELL_X2 FILLER_19_4 ();
 FILLCELL_X4 FILLER_19_36 ();
 FILLCELL_X8 FILLER_19_44 ();
 FILLCELL_X4 FILLER_19_52 ();
 FILLCELL_X2 FILLER_19_56 ();
 FILLCELL_X4 FILLER_19_68 ();
 FILLCELL_X2 FILLER_19_72 ();
 FILLCELL_X8 FILLER_19_87 ();
 FILLCELL_X2 FILLER_19_95 ();
 FILLCELL_X4 FILLER_19_107 ();
 FILLCELL_X4 FILLER_19_115 ();
 FILLCELL_X1 FILLER_19_119 ();
 FILLCELL_X1 FILLER_19_136 ();
 FILLCELL_X2 FILLER_19_151 ();
 FILLCELL_X1 FILLER_19_153 ();
 FILLCELL_X8 FILLER_19_160 ();
 FILLCELL_X4 FILLER_19_168 ();
 FILLCELL_X2 FILLER_19_172 ();
 FILLCELL_X2 FILLER_19_189 ();
 FILLCELL_X2 FILLER_19_216 ();
 FILLCELL_X2 FILLER_19_247 ();
 FILLCELL_X8 FILLER_19_258 ();
 FILLCELL_X4 FILLER_19_266 ();
 FILLCELL_X1 FILLER_19_270 ();
 FILLCELL_X16 FILLER_19_281 ();
 FILLCELL_X4 FILLER_19_297 ();
 FILLCELL_X2 FILLER_19_301 ();
 FILLCELL_X4 FILLER_19_314 ();
 FILLCELL_X2 FILLER_19_318 ();
 FILLCELL_X1 FILLER_19_320 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_3 ();
 FILLCELL_X16 FILLER_20_7 ();
 FILLCELL_X4 FILLER_20_23 ();
 FILLCELL_X1 FILLER_20_27 ();
 FILLCELL_X4 FILLER_20_35 ();
 FILLCELL_X2 FILLER_20_42 ();
 FILLCELL_X1 FILLER_20_44 ();
 FILLCELL_X8 FILLER_20_49 ();
 FILLCELL_X2 FILLER_20_57 ();
 FILLCELL_X1 FILLER_20_59 ();
 FILLCELL_X4 FILLER_20_69 ();
 FILLCELL_X2 FILLER_20_73 ();
 FILLCELL_X8 FILLER_20_88 ();
 FILLCELL_X4 FILLER_20_96 ();
 FILLCELL_X1 FILLER_20_100 ();
 FILLCELL_X1 FILLER_20_114 ();
 FILLCELL_X1 FILLER_20_118 ();
 FILLCELL_X1 FILLER_20_123 ();
 FILLCELL_X2 FILLER_20_131 ();
 FILLCELL_X2 FILLER_20_140 ();
 FILLCELL_X1 FILLER_20_142 ();
 FILLCELL_X2 FILLER_20_161 ();
 FILLCELL_X2 FILLER_20_175 ();
 FILLCELL_X1 FILLER_20_187 ();
 FILLCELL_X2 FILLER_20_197 ();
 FILLCELL_X1 FILLER_20_199 ();
 FILLCELL_X1 FILLER_20_204 ();
 FILLCELL_X4 FILLER_20_219 ();
 FILLCELL_X2 FILLER_20_223 ();
 FILLCELL_X4 FILLER_20_234 ();
 FILLCELL_X2 FILLER_20_238 ();
 FILLCELL_X1 FILLER_20_240 ();
 FILLCELL_X1 FILLER_20_280 ();
 FILLCELL_X8 FILLER_20_285 ();
 FILLCELL_X2 FILLER_20_293 ();
 FILLCELL_X1 FILLER_20_298 ();
 FILLCELL_X8 FILLER_20_309 ();
 FILLCELL_X4 FILLER_20_317 ();
 FILLCELL_X2 FILLER_20_321 ();
 FILLCELL_X1 FILLER_20_323 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_6 ();
 FILLCELL_X4 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_18 ();
 FILLCELL_X2 FILLER_21_23 ();
 FILLCELL_X8 FILLER_21_32 ();
 FILLCELL_X1 FILLER_21_40 ();
 FILLCELL_X8 FILLER_21_60 ();
 FILLCELL_X2 FILLER_21_68 ();
 FILLCELL_X16 FILLER_21_75 ();
 FILLCELL_X8 FILLER_21_91 ();
 FILLCELL_X2 FILLER_21_99 ();
 FILLCELL_X16 FILLER_21_116 ();
 FILLCELL_X1 FILLER_21_132 ();
 FILLCELL_X4 FILLER_21_138 ();
 FILLCELL_X2 FILLER_21_142 ();
 FILLCELL_X1 FILLER_21_172 ();
 FILLCELL_X8 FILLER_21_207 ();
 FILLCELL_X4 FILLER_21_215 ();
 FILLCELL_X1 FILLER_21_219 ();
 FILLCELL_X4 FILLER_21_224 ();
 FILLCELL_X4 FILLER_21_232 ();
 FILLCELL_X2 FILLER_21_236 ();
 FILLCELL_X2 FILLER_21_241 ();
 FILLCELL_X8 FILLER_21_253 ();
 FILLCELL_X4 FILLER_21_261 ();
 FILLCELL_X2 FILLER_21_265 ();
 FILLCELL_X1 FILLER_21_267 ();
 FILLCELL_X1 FILLER_21_283 ();
 FILLCELL_X2 FILLER_21_307 ();
 FILLCELL_X1 FILLER_21_309 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_9 ();
 FILLCELL_X16 FILLER_22_27 ();
 FILLCELL_X4 FILLER_22_43 ();
 FILLCELL_X2 FILLER_22_47 ();
 FILLCELL_X1 FILLER_22_49 ();
 FILLCELL_X8 FILLER_22_61 ();
 FILLCELL_X2 FILLER_22_81 ();
 FILLCELL_X2 FILLER_22_85 ();
 FILLCELL_X4 FILLER_22_97 ();
 FILLCELL_X2 FILLER_22_101 ();
 FILLCELL_X1 FILLER_22_112 ();
 FILLCELL_X8 FILLER_22_116 ();
 FILLCELL_X2 FILLER_22_124 ();
 FILLCELL_X1 FILLER_22_126 ();
 FILLCELL_X1 FILLER_22_139 ();
 FILLCELL_X1 FILLER_22_147 ();
 FILLCELL_X8 FILLER_22_247 ();
 FILLCELL_X4 FILLER_22_255 ();
 FILLCELL_X4 FILLER_22_266 ();
 FILLCELL_X1 FILLER_22_270 ();
 FILLCELL_X8 FILLER_22_286 ();
 FILLCELL_X4 FILLER_22_294 ();
 FILLCELL_X2 FILLER_22_298 ();
 FILLCELL_X1 FILLER_22_300 ();
 FILLCELL_X2 FILLER_22_321 ();
 FILLCELL_X1 FILLER_22_323 ();
 FILLCELL_X2 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_3 ();
 FILLCELL_X2 FILLER_23_7 ();
 FILLCELL_X1 FILLER_23_13 ();
 FILLCELL_X2 FILLER_23_21 ();
 FILLCELL_X4 FILLER_23_26 ();
 FILLCELL_X2 FILLER_23_30 ();
 FILLCELL_X2 FILLER_23_36 ();
 FILLCELL_X8 FILLER_23_45 ();
 FILLCELL_X4 FILLER_23_53 ();
 FILLCELL_X2 FILLER_23_57 ();
 FILLCELL_X1 FILLER_23_86 ();
 FILLCELL_X4 FILLER_23_90 ();
 FILLCELL_X1 FILLER_23_94 ();
 FILLCELL_X2 FILLER_23_116 ();
 FILLCELL_X1 FILLER_23_118 ();
 FILLCELL_X4 FILLER_23_129 ();
 FILLCELL_X2 FILLER_23_133 ();
 FILLCELL_X1 FILLER_23_138 ();
 FILLCELL_X8 FILLER_23_185 ();
 FILLCELL_X1 FILLER_23_193 ();
 FILLCELL_X4 FILLER_23_215 ();
 FILLCELL_X2 FILLER_23_222 ();
 FILLCELL_X1 FILLER_23_224 ();
 FILLCELL_X1 FILLER_23_230 ();
 FILLCELL_X8 FILLER_23_234 ();
 FILLCELL_X4 FILLER_23_242 ();
 FILLCELL_X2 FILLER_23_246 ();
 FILLCELL_X4 FILLER_23_254 ();
 FILLCELL_X2 FILLER_23_277 ();
 FILLCELL_X1 FILLER_23_279 ();
 FILLCELL_X2 FILLER_23_305 ();
 FILLCELL_X8 FILLER_23_314 ();
 FILLCELL_X2 FILLER_23_322 ();
 FILLCELL_X4 FILLER_24_18 ();
 FILLCELL_X2 FILLER_24_22 ();
 FILLCELL_X1 FILLER_24_24 ();
 FILLCELL_X4 FILLER_24_45 ();
 FILLCELL_X2 FILLER_24_49 ();
 FILLCELL_X1 FILLER_24_51 ();
 FILLCELL_X16 FILLER_24_71 ();
 FILLCELL_X2 FILLER_24_87 ();
 FILLCELL_X1 FILLER_24_89 ();
 FILLCELL_X4 FILLER_24_101 ();
 FILLCELL_X8 FILLER_24_117 ();
 FILLCELL_X4 FILLER_24_125 ();
 FILLCELL_X2 FILLER_24_129 ();
 FILLCELL_X2 FILLER_24_141 ();
 FILLCELL_X8 FILLER_24_197 ();
 FILLCELL_X4 FILLER_24_205 ();
 FILLCELL_X2 FILLER_24_213 ();
 FILLCELL_X1 FILLER_24_215 ();
 FILLCELL_X1 FILLER_24_228 ();
 FILLCELL_X4 FILLER_24_245 ();
 FILLCELL_X1 FILLER_24_249 ();
 FILLCELL_X1 FILLER_24_261 ();
 FILLCELL_X1 FILLER_24_269 ();
 FILLCELL_X1 FILLER_24_282 ();
 FILLCELL_X4 FILLER_24_288 ();
 FILLCELL_X2 FILLER_24_292 ();
 FILLCELL_X4 FILLER_24_298 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_9 ();
 FILLCELL_X4 FILLER_25_16 ();
 FILLCELL_X2 FILLER_25_20 ();
 FILLCELL_X1 FILLER_25_22 ();
 FILLCELL_X4 FILLER_25_43 ();
 FILLCELL_X2 FILLER_25_47 ();
 FILLCELL_X8 FILLER_25_56 ();
 FILLCELL_X2 FILLER_25_76 ();
 FILLCELL_X1 FILLER_25_104 ();
 FILLCELL_X8 FILLER_25_110 ();
 FILLCELL_X4 FILLER_25_118 ();
 FILLCELL_X2 FILLER_25_122 ();
 FILLCELL_X1 FILLER_25_124 ();
 FILLCELL_X1 FILLER_25_142 ();
 FILLCELL_X1 FILLER_25_177 ();
 FILLCELL_X16 FILLER_25_209 ();
 FILLCELL_X8 FILLER_25_225 ();
 FILLCELL_X1 FILLER_25_233 ();
 FILLCELL_X1 FILLER_25_261 ();
 FILLCELL_X8 FILLER_25_294 ();
 FILLCELL_X8 FILLER_25_309 ();
 FILLCELL_X4 FILLER_25_317 ();
 FILLCELL_X2 FILLER_25_321 ();
 FILLCELL_X1 FILLER_25_323 ();
 FILLCELL_X2 FILLER_26_18 ();
 FILLCELL_X1 FILLER_26_20 ();
 FILLCELL_X2 FILLER_26_34 ();
 FILLCELL_X2 FILLER_26_41 ();
 FILLCELL_X1 FILLER_26_43 ();
 FILLCELL_X1 FILLER_26_75 ();
 FILLCELL_X4 FILLER_26_83 ();
 FILLCELL_X2 FILLER_26_87 ();
 FILLCELL_X2 FILLER_26_106 ();
 FILLCELL_X1 FILLER_26_108 ();
 FILLCELL_X1 FILLER_26_175 ();
 FILLCELL_X1 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_197 ();
 FILLCELL_X1 FILLER_26_205 ();
 FILLCELL_X1 FILLER_26_221 ();
 FILLCELL_X16 FILLER_26_225 ();
 FILLCELL_X4 FILLER_26_241 ();
 FILLCELL_X1 FILLER_26_245 ();
 FILLCELL_X1 FILLER_26_260 ();
 FILLCELL_X4 FILLER_26_264 ();
 FILLCELL_X2 FILLER_26_268 ();
 FILLCELL_X1 FILLER_26_274 ();
 FILLCELL_X2 FILLER_26_295 ();
 FILLCELL_X1 FILLER_26_297 ();
 FILLCELL_X2 FILLER_26_301 ();
 FILLCELL_X1 FILLER_26_303 ();
 FILLCELL_X8 FILLER_26_311 ();
 FILLCELL_X2 FILLER_26_319 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X8 FILLER_27_8 ();
 FILLCELL_X1 FILLER_27_16 ();
 FILLCELL_X1 FILLER_27_38 ();
 FILLCELL_X8 FILLER_27_46 ();
 FILLCELL_X4 FILLER_27_54 ();
 FILLCELL_X2 FILLER_27_58 ();
 FILLCELL_X16 FILLER_27_67 ();
 FILLCELL_X2 FILLER_27_83 ();
 FILLCELL_X2 FILLER_27_95 ();
 FILLCELL_X8 FILLER_27_104 ();
 FILLCELL_X4 FILLER_27_112 ();
 FILLCELL_X1 FILLER_27_116 ();
 FILLCELL_X1 FILLER_27_164 ();
 FILLCELL_X1 FILLER_27_188 ();
 FILLCELL_X1 FILLER_27_192 ();
 FILLCELL_X4 FILLER_27_197 ();
 FILLCELL_X2 FILLER_27_219 ();
 FILLCELL_X4 FILLER_27_225 ();
 FILLCELL_X2 FILLER_27_229 ();
 FILLCELL_X1 FILLER_27_231 ();
 FILLCELL_X4 FILLER_27_237 ();
 FILLCELL_X2 FILLER_27_252 ();
 FILLCELL_X8 FILLER_27_273 ();
 FILLCELL_X16 FILLER_27_285 ();
 FILLCELL_X2 FILLER_27_301 ();
 FILLCELL_X1 FILLER_27_303 ();
 FILLCELL_X2 FILLER_27_321 ();
 FILLCELL_X1 FILLER_27_323 ();
 FILLCELL_X2 FILLER_28_1 ();
 FILLCELL_X8 FILLER_28_30 ();
 FILLCELL_X2 FILLER_28_38 ();
 FILLCELL_X1 FILLER_28_40 ();
 FILLCELL_X8 FILLER_28_60 ();
 FILLCELL_X1 FILLER_28_68 ();
 FILLCELL_X1 FILLER_28_72 ();
 FILLCELL_X2 FILLER_28_93 ();
 FILLCELL_X1 FILLER_28_95 ();
 FILLCELL_X16 FILLER_28_113 ();
 FILLCELL_X8 FILLER_28_129 ();
 FILLCELL_X2 FILLER_28_137 ();
 FILLCELL_X8 FILLER_28_141 ();
 FILLCELL_X1 FILLER_28_160 ();
 FILLCELL_X4 FILLER_28_176 ();
 FILLCELL_X1 FILLER_28_180 ();
 FILLCELL_X1 FILLER_28_216 ();
 FILLCELL_X8 FILLER_28_241 ();
 FILLCELL_X2 FILLER_28_249 ();
 FILLCELL_X1 FILLER_28_251 ();
 FILLCELL_X2 FILLER_28_256 ();
 FILLCELL_X1 FILLER_28_258 ();
 FILLCELL_X4 FILLER_28_273 ();
 FILLCELL_X1 FILLER_28_296 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_8 ();
 FILLCELL_X4 FILLER_29_37 ();
 FILLCELL_X8 FILLER_29_44 ();
 FILLCELL_X4 FILLER_29_52 ();
 FILLCELL_X16 FILLER_29_79 ();
 FILLCELL_X1 FILLER_29_95 ();
 FILLCELL_X16 FILLER_29_123 ();
 FILLCELL_X4 FILLER_29_153 ();
 FILLCELL_X2 FILLER_29_170 ();
 FILLCELL_X8 FILLER_29_179 ();
 FILLCELL_X4 FILLER_29_187 ();
 FILLCELL_X2 FILLER_29_191 ();
 FILLCELL_X2 FILLER_29_196 ();
 FILLCELL_X1 FILLER_29_198 ();
 FILLCELL_X16 FILLER_29_203 ();
 FILLCELL_X1 FILLER_29_219 ();
 FILLCELL_X8 FILLER_29_232 ();
 FILLCELL_X1 FILLER_29_240 ();
 FILLCELL_X8 FILLER_29_248 ();
 FILLCELL_X4 FILLER_29_256 ();
 FILLCELL_X2 FILLER_29_260 ();
 FILLCELL_X4 FILLER_29_270 ();
 FILLCELL_X2 FILLER_29_274 ();
 FILLCELL_X1 FILLER_29_276 ();
 FILLCELL_X2 FILLER_29_307 ();
 FILLCELL_X4 FILLER_29_313 ();
 FILLCELL_X1 FILLER_29_317 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_9 ();
 FILLCELL_X32 FILLER_30_13 ();
 FILLCELL_X4 FILLER_30_45 ();
 FILLCELL_X2 FILLER_30_59 ();
 FILLCELL_X2 FILLER_30_65 ();
 FILLCELL_X2 FILLER_30_70 ();
 FILLCELL_X1 FILLER_30_72 ();
 FILLCELL_X1 FILLER_30_77 ();
 FILLCELL_X1 FILLER_30_80 ();
 FILLCELL_X8 FILLER_30_93 ();
 FILLCELL_X4 FILLER_30_101 ();
 FILLCELL_X2 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_107 ();
 FILLCELL_X1 FILLER_30_132 ();
 FILLCELL_X4 FILLER_30_143 ();
 FILLCELL_X2 FILLER_30_147 ();
 FILLCELL_X2 FILLER_30_164 ();
 FILLCELL_X2 FILLER_30_202 ();
 FILLCELL_X4 FILLER_30_230 ();
 FILLCELL_X2 FILLER_30_234 ();
 FILLCELL_X1 FILLER_30_236 ();
 FILLCELL_X8 FILLER_30_250 ();
 FILLCELL_X1 FILLER_30_258 ();
 FILLCELL_X8 FILLER_30_278 ();
 FILLCELL_X8 FILLER_30_311 ();
 FILLCELL_X4 FILLER_30_319 ();
 FILLCELL_X1 FILLER_30_323 ();
 FILLCELL_X8 FILLER_31_29 ();
 FILLCELL_X1 FILLER_31_37 ();
 FILLCELL_X1 FILLER_31_41 ();
 FILLCELL_X16 FILLER_31_59 ();
 FILLCELL_X4 FILLER_31_75 ();
 FILLCELL_X2 FILLER_31_79 ();
 FILLCELL_X1 FILLER_31_81 ();
 FILLCELL_X8 FILLER_31_89 ();
 FILLCELL_X1 FILLER_31_97 ();
 FILLCELL_X2 FILLER_31_143 ();
 FILLCELL_X4 FILLER_31_154 ();
 FILLCELL_X1 FILLER_31_161 ();
 FILLCELL_X8 FILLER_31_177 ();
 FILLCELL_X2 FILLER_31_185 ();
 FILLCELL_X8 FILLER_31_191 ();
 FILLCELL_X4 FILLER_31_199 ();
 FILLCELL_X2 FILLER_31_203 ();
 FILLCELL_X2 FILLER_31_211 ();
 FILLCELL_X1 FILLER_31_217 ();
 FILLCELL_X1 FILLER_31_222 ();
 FILLCELL_X1 FILLER_31_230 ();
 FILLCELL_X8 FILLER_31_262 ();
 FILLCELL_X4 FILLER_31_270 ();
 FILLCELL_X2 FILLER_31_274 ();
 FILLCELL_X4 FILLER_31_290 ();
 FILLCELL_X2 FILLER_31_297 ();
 FILLCELL_X1 FILLER_31_306 ();
 FILLCELL_X4 FILLER_32_1 ();
 FILLCELL_X2 FILLER_32_5 ();
 FILLCELL_X1 FILLER_32_7 ();
 FILLCELL_X16 FILLER_32_11 ();
 FILLCELL_X1 FILLER_32_27 ();
 FILLCELL_X2 FILLER_32_35 ();
 FILLCELL_X2 FILLER_32_42 ();
 FILLCELL_X1 FILLER_32_48 ();
 FILLCELL_X4 FILLER_32_52 ();
 FILLCELL_X2 FILLER_32_56 ();
 FILLCELL_X1 FILLER_32_58 ();
 FILLCELL_X1 FILLER_32_65 ();
 FILLCELL_X1 FILLER_32_68 ();
 FILLCELL_X1 FILLER_32_76 ();
 FILLCELL_X16 FILLER_32_87 ();
 FILLCELL_X4 FILLER_32_103 ();
 FILLCELL_X4 FILLER_32_135 ();
 FILLCELL_X2 FILLER_32_144 ();
 FILLCELL_X1 FILLER_32_146 ();
 FILLCELL_X16 FILLER_32_167 ();
 FILLCELL_X2 FILLER_32_183 ();
 FILLCELL_X1 FILLER_32_201 ();
 FILLCELL_X2 FILLER_32_209 ();
 FILLCELL_X1 FILLER_32_211 ();
 FILLCELL_X1 FILLER_32_218 ();
 FILLCELL_X1 FILLER_32_223 ();
 FILLCELL_X8 FILLER_32_234 ();
 FILLCELL_X4 FILLER_32_242 ();
 FILLCELL_X1 FILLER_32_246 ();
 FILLCELL_X8 FILLER_32_263 ();
 FILLCELL_X2 FILLER_32_271 ();
 FILLCELL_X4 FILLER_32_277 ();
 FILLCELL_X8 FILLER_32_309 ();
 FILLCELL_X1 FILLER_32_317 ();
 FILLCELL_X4 FILLER_33_4 ();
 FILLCELL_X2 FILLER_33_8 ();
 FILLCELL_X1 FILLER_33_24 ();
 FILLCELL_X8 FILLER_33_57 ();
 FILLCELL_X2 FILLER_33_65 ();
 FILLCELL_X1 FILLER_33_67 ();
 FILLCELL_X2 FILLER_33_74 ();
 FILLCELL_X2 FILLER_33_90 ();
 FILLCELL_X2 FILLER_33_100 ();
 FILLCELL_X8 FILLER_33_134 ();
 FILLCELL_X1 FILLER_33_152 ();
 FILLCELL_X1 FILLER_33_163 ();
 FILLCELL_X8 FILLER_33_169 ();
 FILLCELL_X4 FILLER_33_177 ();
 FILLCELL_X2 FILLER_33_181 ();
 FILLCELL_X1 FILLER_33_183 ();
 FILLCELL_X4 FILLER_33_187 ();
 FILLCELL_X2 FILLER_33_191 ();
 FILLCELL_X1 FILLER_33_193 ();
 FILLCELL_X4 FILLER_33_203 ();
 FILLCELL_X2 FILLER_33_207 ();
 FILLCELL_X1 FILLER_33_209 ();
 FILLCELL_X2 FILLER_33_226 ();
 FILLCELL_X1 FILLER_33_228 ();
 FILLCELL_X2 FILLER_33_247 ();
 FILLCELL_X16 FILLER_33_252 ();
 FILLCELL_X4 FILLER_33_268 ();
 FILLCELL_X2 FILLER_33_302 ();
 FILLCELL_X1 FILLER_33_304 ();
 FILLCELL_X8 FILLER_33_312 ();
 FILLCELL_X1 FILLER_33_320 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X2 FILLER_34_5 ();
 FILLCELL_X1 FILLER_34_7 ();
 FILLCELL_X2 FILLER_34_11 ();
 FILLCELL_X1 FILLER_34_13 ();
 FILLCELL_X16 FILLER_34_49 ();
 FILLCELL_X4 FILLER_34_65 ();
 FILLCELL_X2 FILLER_34_71 ();
 FILLCELL_X1 FILLER_34_73 ();
 FILLCELL_X8 FILLER_34_79 ();
 FILLCELL_X2 FILLER_34_87 ();
 FILLCELL_X2 FILLER_34_106 ();
 FILLCELL_X4 FILLER_34_128 ();
 FILLCELL_X1 FILLER_34_135 ();
 FILLCELL_X4 FILLER_34_158 ();
 FILLCELL_X1 FILLER_34_162 ();
 FILLCELL_X8 FILLER_34_170 ();
 FILLCELL_X2 FILLER_34_178 ();
 FILLCELL_X4 FILLER_34_203 ();
 FILLCELL_X2 FILLER_34_207 ();
 FILLCELL_X1 FILLER_34_209 ();
 FILLCELL_X1 FILLER_34_217 ();
 FILLCELL_X2 FILLER_34_222 ();
 FILLCELL_X1 FILLER_34_224 ();
 FILLCELL_X2 FILLER_34_242 ();
 FILLCELL_X1 FILLER_34_244 ();
 FILLCELL_X8 FILLER_34_273 ();
 FILLCELL_X2 FILLER_34_281 ();
 FILLCELL_X2 FILLER_34_288 ();
 FILLCELL_X2 FILLER_34_301 ();
 FILLCELL_X1 FILLER_34_303 ();
 FILLCELL_X2 FILLER_34_321 ();
 FILLCELL_X1 FILLER_34_323 ();
 FILLCELL_X4 FILLER_35_1 ();
 FILLCELL_X4 FILLER_35_8 ();
 FILLCELL_X2 FILLER_35_12 ();
 FILLCELL_X1 FILLER_35_14 ();
 FILLCELL_X2 FILLER_35_22 ();
 FILLCELL_X1 FILLER_35_24 ();
 FILLCELL_X4 FILLER_35_32 ();
 FILLCELL_X2 FILLER_35_36 ();
 FILLCELL_X1 FILLER_35_38 ();
 FILLCELL_X8 FILLER_35_43 ();
 FILLCELL_X2 FILLER_35_71 ();
 FILLCELL_X1 FILLER_35_73 ();
 FILLCELL_X2 FILLER_35_91 ();
 FILLCELL_X16 FILLER_35_99 ();
 FILLCELL_X4 FILLER_35_115 ();
 FILLCELL_X2 FILLER_35_119 ();
 FILLCELL_X1 FILLER_35_121 ();
 FILLCELL_X2 FILLER_35_129 ();
 FILLCELL_X1 FILLER_35_131 ();
 FILLCELL_X8 FILLER_35_139 ();
 FILLCELL_X4 FILLER_35_147 ();
 FILLCELL_X2 FILLER_35_151 ();
 FILLCELL_X1 FILLER_35_153 ();
 FILLCELL_X2 FILLER_35_156 ();
 FILLCELL_X1 FILLER_35_165 ();
 FILLCELL_X1 FILLER_35_169 ();
 FILLCELL_X1 FILLER_35_187 ();
 FILLCELL_X1 FILLER_35_191 ();
 FILLCELL_X1 FILLER_35_198 ();
 FILLCELL_X4 FILLER_35_202 ();
 FILLCELL_X1 FILLER_35_206 ();
 FILLCELL_X1 FILLER_35_227 ();
 FILLCELL_X2 FILLER_35_235 ();
 FILLCELL_X16 FILLER_35_248 ();
 FILLCELL_X4 FILLER_35_264 ();
 FILLCELL_X8 FILLER_35_285 ();
 FILLCELL_X4 FILLER_35_313 ();
 FILLCELL_X4 FILLER_35_320 ();
 FILLCELL_X2 FILLER_36_22 ();
 FILLCELL_X8 FILLER_36_28 ();
 FILLCELL_X1 FILLER_36_63 ();
 FILLCELL_X1 FILLER_36_66 ();
 FILLCELL_X2 FILLER_36_71 ();
 FILLCELL_X2 FILLER_36_80 ();
 FILLCELL_X2 FILLER_36_89 ();
 FILLCELL_X16 FILLER_36_104 ();
 FILLCELL_X1 FILLER_36_120 ();
 FILLCELL_X2 FILLER_36_127 ();
 FILLCELL_X1 FILLER_36_129 ();
 FILLCELL_X8 FILLER_36_151 ();
 FILLCELL_X4 FILLER_36_159 ();
 FILLCELL_X1 FILLER_36_163 ();
 FILLCELL_X1 FILLER_36_183 ();
 FILLCELL_X8 FILLER_36_187 ();
 FILLCELL_X2 FILLER_36_195 ();
 FILLCELL_X1 FILLER_36_197 ();
 FILLCELL_X4 FILLER_36_202 ();
 FILLCELL_X1 FILLER_36_206 ();
 FILLCELL_X1 FILLER_36_226 ();
 FILLCELL_X8 FILLER_36_237 ();
 FILLCELL_X32 FILLER_36_262 ();
 FILLCELL_X16 FILLER_36_294 ();
 FILLCELL_X8 FILLER_36_310 ();
 FILLCELL_X4 FILLER_36_318 ();
 FILLCELL_X2 FILLER_36_322 ();
 FILLCELL_X4 FILLER_37_1 ();
 FILLCELL_X1 FILLER_37_5 ();
 FILLCELL_X32 FILLER_37_26 ();
 FILLCELL_X4 FILLER_37_58 ();
 FILLCELL_X2 FILLER_37_62 ();
 FILLCELL_X1 FILLER_37_70 ();
 FILLCELL_X2 FILLER_37_75 ();
 FILLCELL_X2 FILLER_37_81 ();
 FILLCELL_X1 FILLER_37_83 ();
 FILLCELL_X4 FILLER_37_88 ();
 FILLCELL_X2 FILLER_37_92 ();
 FILLCELL_X8 FILLER_37_98 ();
 FILLCELL_X2 FILLER_37_123 ();
 FILLCELL_X4 FILLER_37_136 ();
 FILLCELL_X16 FILLER_37_152 ();
 FILLCELL_X8 FILLER_37_168 ();
 FILLCELL_X2 FILLER_37_176 ();
 FILLCELL_X16 FILLER_37_187 ();
 FILLCELL_X4 FILLER_37_203 ();
 FILLCELL_X2 FILLER_37_207 ();
 FILLCELL_X32 FILLER_37_238 ();
 FILLCELL_X32 FILLER_37_270 ();
 FILLCELL_X16 FILLER_37_302 ();
 FILLCELL_X4 FILLER_37_318 ();
 FILLCELL_X2 FILLER_37_322 ();
 FILLCELL_X16 FILLER_38_1 ();
 FILLCELL_X2 FILLER_38_17 ();
 FILLCELL_X1 FILLER_38_19 ();
 FILLCELL_X2 FILLER_38_23 ();
 FILLCELL_X1 FILLER_38_25 ();
 FILLCELL_X1 FILLER_38_54 ();
 FILLCELL_X1 FILLER_38_71 ();
 FILLCELL_X2 FILLER_38_83 ();
 FILLCELL_X1 FILLER_38_85 ();
 FILLCELL_X8 FILLER_38_109 ();
 FILLCELL_X2 FILLER_38_117 ();
 FILLCELL_X1 FILLER_38_119 ();
 FILLCELL_X8 FILLER_38_137 ();
 FILLCELL_X2 FILLER_38_149 ();
 FILLCELL_X4 FILLER_38_177 ();
 FILLCELL_X4 FILLER_38_188 ();
 FILLCELL_X2 FILLER_38_192 ();
 FILLCELL_X1 FILLER_38_194 ();
 FILLCELL_X2 FILLER_38_206 ();
 FILLCELL_X2 FILLER_38_218 ();
 FILLCELL_X2 FILLER_38_224 ();
 FILLCELL_X1 FILLER_38_226 ();
 FILLCELL_X2 FILLER_38_236 ();
 FILLCELL_X1 FILLER_38_238 ();
 FILLCELL_X8 FILLER_38_246 ();
 FILLCELL_X4 FILLER_38_254 ();
 FILLCELL_X32 FILLER_38_269 ();
 FILLCELL_X16 FILLER_38_301 ();
 FILLCELL_X4 FILLER_38_317 ();
 FILLCELL_X2 FILLER_38_321 ();
 FILLCELL_X1 FILLER_38_323 ();
 FILLCELL_X16 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_17 ();
 FILLCELL_X1 FILLER_39_19 ();
 FILLCELL_X8 FILLER_39_37 ();
 FILLCELL_X4 FILLER_39_45 ();
 FILLCELL_X1 FILLER_39_49 ();
 FILLCELL_X2 FILLER_39_64 ();
 FILLCELL_X1 FILLER_39_66 ();
 FILLCELL_X8 FILLER_39_79 ();
 FILLCELL_X2 FILLER_39_87 ();
 FILLCELL_X1 FILLER_39_89 ();
 FILLCELL_X4 FILLER_39_120 ();
 FILLCELL_X2 FILLER_39_124 ();
 FILLCELL_X1 FILLER_39_126 ();
 FILLCELL_X8 FILLER_39_136 ();
 FILLCELL_X2 FILLER_39_144 ();
 FILLCELL_X1 FILLER_39_146 ();
 FILLCELL_X2 FILLER_39_156 ();
 FILLCELL_X1 FILLER_39_158 ();
 FILLCELL_X1 FILLER_39_184 ();
 FILLCELL_X1 FILLER_39_198 ();
 FILLCELL_X8 FILLER_39_203 ();
 FILLCELL_X4 FILLER_39_211 ();
 FILLCELL_X8 FILLER_39_224 ();
 FILLCELL_X4 FILLER_39_256 ();
 FILLCELL_X2 FILLER_39_260 ();
 FILLCELL_X1 FILLER_39_262 ();
 FILLCELL_X32 FILLER_39_280 ();
 FILLCELL_X8 FILLER_39_312 ();
 FILLCELL_X4 FILLER_39_320 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_17 ();
 FILLCELL_X4 FILLER_40_25 ();
 FILLCELL_X8 FILLER_40_40 ();
 FILLCELL_X8 FILLER_40_55 ();
 FILLCELL_X1 FILLER_40_63 ();
 FILLCELL_X8 FILLER_40_67 ();
 FILLCELL_X2 FILLER_40_75 ();
 FILLCELL_X8 FILLER_40_80 ();
 FILLCELL_X4 FILLER_40_88 ();
 FILLCELL_X2 FILLER_40_92 ();
 FILLCELL_X1 FILLER_40_94 ();
 FILLCELL_X8 FILLER_40_104 ();
 FILLCELL_X4 FILLER_40_112 ();
 FILLCELL_X4 FILLER_40_136 ();
 FILLCELL_X2 FILLER_40_140 ();
 FILLCELL_X1 FILLER_40_142 ();
 FILLCELL_X4 FILLER_40_147 ();
 FILLCELL_X1 FILLER_40_151 ();
 FILLCELL_X4 FILLER_40_155 ();
 FILLCELL_X2 FILLER_40_159 ();
 FILLCELL_X1 FILLER_40_170 ();
 FILLCELL_X1 FILLER_40_175 ();
 FILLCELL_X1 FILLER_40_181 ();
 FILLCELL_X2 FILLER_40_193 ();
 FILLCELL_X4 FILLER_40_201 ();
 FILLCELL_X2 FILLER_40_208 ();
 FILLCELL_X4 FILLER_40_217 ();
 FILLCELL_X2 FILLER_40_221 ();
 FILLCELL_X1 FILLER_40_223 ();
 FILLCELL_X2 FILLER_40_245 ();
 FILLCELL_X1 FILLER_40_247 ();
 FILLCELL_X8 FILLER_40_252 ();
 FILLCELL_X1 FILLER_40_260 ();
 FILLCELL_X32 FILLER_40_278 ();
 FILLCELL_X8 FILLER_40_310 ();
 FILLCELL_X4 FILLER_40_318 ();
 FILLCELL_X2 FILLER_40_322 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X1 FILLER_41_17 ();
 FILLCELL_X1 FILLER_41_35 ();
 FILLCELL_X1 FILLER_41_53 ();
 FILLCELL_X1 FILLER_41_64 ();
 FILLCELL_X4 FILLER_41_69 ();
 FILLCELL_X2 FILLER_41_73 ();
 FILLCELL_X1 FILLER_41_75 ();
 FILLCELL_X4 FILLER_41_86 ();
 FILLCELL_X2 FILLER_41_90 ();
 FILLCELL_X1 FILLER_41_92 ();
 FILLCELL_X4 FILLER_41_99 ();
 FILLCELL_X16 FILLER_41_107 ();
 FILLCELL_X8 FILLER_41_123 ();
 FILLCELL_X1 FILLER_41_131 ();
 FILLCELL_X1 FILLER_41_152 ();
 FILLCELL_X1 FILLER_41_170 ();
 FILLCELL_X2 FILLER_41_185 ();
 FILLCELL_X2 FILLER_41_231 ();
 FILLCELL_X2 FILLER_41_236 ();
 FILLCELL_X32 FILLER_41_269 ();
 FILLCELL_X16 FILLER_41_301 ();
 FILLCELL_X4 FILLER_41_317 ();
 FILLCELL_X2 FILLER_41_321 ();
 FILLCELL_X1 FILLER_41_323 ();
 FILLCELL_X16 FILLER_42_1 ();
 FILLCELL_X8 FILLER_42_17 ();
 FILLCELL_X4 FILLER_42_25 ();
 FILLCELL_X1 FILLER_42_29 ();
 FILLCELL_X8 FILLER_42_33 ();
 FILLCELL_X4 FILLER_42_41 ();
 FILLCELL_X2 FILLER_42_45 ();
 FILLCELL_X1 FILLER_42_47 ();
 FILLCELL_X2 FILLER_42_51 ();
 FILLCELL_X4 FILLER_42_59 ();
 FILLCELL_X1 FILLER_42_63 ();
 FILLCELL_X4 FILLER_42_81 ();
 FILLCELL_X1 FILLER_42_85 ();
 FILLCELL_X4 FILLER_42_96 ();
 FILLCELL_X2 FILLER_42_100 ();
 FILLCELL_X4 FILLER_42_119 ();
 FILLCELL_X2 FILLER_42_123 ();
 FILLCELL_X1 FILLER_42_125 ();
 FILLCELL_X32 FILLER_42_130 ();
 FILLCELL_X4 FILLER_42_162 ();
 FILLCELL_X32 FILLER_42_170 ();
 FILLCELL_X4 FILLER_42_202 ();
 FILLCELL_X1 FILLER_42_206 ();
 FILLCELL_X2 FILLER_42_210 ();
 FILLCELL_X1 FILLER_42_212 ();
 FILLCELL_X8 FILLER_42_216 ();
 FILLCELL_X2 FILLER_42_224 ();
 FILLCELL_X1 FILLER_42_229 ();
 FILLCELL_X2 FILLER_42_243 ();
 FILLCELL_X8 FILLER_42_248 ();
 FILLCELL_X2 FILLER_42_262 ();
 FILLCELL_X1 FILLER_42_264 ();
 FILLCELL_X8 FILLER_42_269 ();
 FILLCELL_X32 FILLER_42_283 ();
 FILLCELL_X8 FILLER_42_315 ();
 FILLCELL_X1 FILLER_42_323 ();
endmodule
