module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire net1519;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire clknet_2_0_0_clk;
 wire _00943_;
 wire _00944_;
 wire net2112;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire net1676;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire net1703;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire net1704;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire clknet_leaf_30_clk_i_regs;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire net1693;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire clknet_2_0__leaf_clk_i_regs;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire clknet_leaf_2_clk;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire net1683;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire net1682;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire clknet_leaf_4_clk;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire clknet_leaf_5_clk;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire net1680;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire net1679;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire net1518;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire net1454;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire net1468;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire net1453;
 wire net1471;
 wire _03452_;
 wire net1452;
 wire net1479;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire net1481;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire net1483;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire net1451;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire net1450;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire net1449;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire net1448;
 wire _03506_;
 wire net1447;
 wire _03508_;
 wire net1446;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire net2162;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire net2163;
 wire _03520_;
 wire _03521_;
 wire net2164;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire net2165;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire net2166;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire net2167;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire net2168;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire net2169;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire net2170;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire net1445;
 wire net1444;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire net2171;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire net1443;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire net1442;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire net1441;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire net2172;
 wire _03905_;
 wire _03906_;
 wire net1440;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire net1439;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire net1438;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire net1437;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire net1436;
 wire _03943_;
 wire _03944_;
 wire net1435;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire net1434;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire net1433;
 wire _03977_;
 wire _03978_;
 wire net2173;
 wire net2174;
 wire _03981_;
 wire net1432;
 wire _03983_;
 wire _03984_;
 wire net2175;
 wire net1431;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire net2204;
 wire net1429;
 wire _03992_;
 wire net1428;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire net2176;
 wire net1427;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire net1426;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire net2177;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire net2178;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire net2179;
 wire _04046_;
 wire net2180;
 wire _04048_;
 wire _04049_;
 wire net2181;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire net2182;
 wire net2183;
 wire _04064_;
 wire _04065_;
 wire net2184;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire net1425;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire net1424;
 wire net1423;
 wire _04088_;
 wire _04089_;
 wire net1422;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire net1421;
 wire net1420;
 wire _04135_;
 wire net2185;
 wire _04137_;
 wire _04138_;
 wire net1419;
 wire net1418;
 wire net1416;
 wire net1415;
 wire net1414;
 wire net1417;
 wire net1413;
 wire _04146_;
 wire net1412;
 wire net2186;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire net2187;
 wire net2188;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire net1411;
 wire _04165_;
 wire _04166_;
 wire net2189;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire net2190;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire net1410;
 wire _04193_;
 wire _04194_;
 wire net2191;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire net2192;
 wire net1409;
 wire _04204_;
 wire _04205_;
 wire net2193;
 wire _04207_;
 wire _04208_;
 wire net1408;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire net1407;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire net2194;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire net2272;
 wire net1405;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire net1406;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire net2276;
 wire _04346_;
 wire net1404;
 wire _04348_;
 wire net1403;
 wire net1402;
 wire net2278;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire net2287;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire net2288;
 wire _04413_;
 wire net2289;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire net2290;
 wire _04433_;
 wire net2291;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire net2292;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire net2293;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire net2298;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire net2299;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire net2300;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire net1401;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire net1400;
 wire net1399;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire net2465;
 wire net2466;
 wire net2467;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire net2468;
 wire _04559_;
 wire _04560_;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2475;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire net2476;
 wire net2477;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire net2478;
 wire _04580_;
 wire _04581_;
 wire net2479;
 wire _04583_;
 wire _04584_;
 wire net2480;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire net2482;
 wire _04592_;
 wire net2493;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire net2492;
 wire net2491;
 wire _04599_;
 wire _04600_;
 wire net2484;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire net2483;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire net2495;
 wire _04614_;
 wire _04615_;
 wire net2494;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire net1398;
 wire _04651_;
 wire _04653_;
 wire _04656_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire net1397;
 wire _04672_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire net1396;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04703_;
 wire _04704_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04773_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04841_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04858_;
 wire _04860_;
 wire _04862_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire net1395;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire net1393;
 wire net1392;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire net1391;
 wire _04966_;
 wire net1394;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire net1390;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04986_;
 wire _04988_;
 wire _04989_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire net1389;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire net1388;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire net1387;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire net1386;
 wire net1385;
 wire net1384;
 wire net1383;
 wire net1382;
 wire net1380;
 wire net1379;
 wire net1381;
 wire net1378;
 wire net1377;
 wire net1376;
 wire net1375;
 wire net1374;
 wire net1372;
 wire net1371;
 wire net1370;
 wire net1369;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire net1367;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire net1366;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire net2474;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire net1364;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire net1363;
 wire net1361;
 wire net1360;
 wire net1359;
 wire net1357;
 wire net1355;
 wire net1354;
 wire _05573_;
 wire _05574_;
 wire net1353;
 wire net1352;
 wire net1351;
 wire _05578_;
 wire _05579_;
 wire net1350;
 wire net1349;
 wire net1358;
 wire net1356;
 wire _05584_;
 wire net1348;
 wire net2042;
 wire net2027;
 wire net2023;
 wire net2026;
 wire net2034;
 wire _05591_;
 wire _05592_;
 wire net2021;
 wire net2020;
 wire net2045;
 wire _05596_;
 wire clknet_leaf_23_clk_i_regs;
 wire net1959;
 wire net1958;
 wire _05600_;
 wire net1960;
 wire _05602_;
 wire net1974;
 wire net1973;
 wire net1972;
 wire _05606_;
 wire net1980;
 wire net1954;
 wire net1878;
 wire _05610_;
 wire net1863;
 wire net1926;
 wire net1805;
 wire _05614_;
 wire net2008;
 wire net1749;
 wire net1660;
 wire net1661;
 wire _05619_;
 wire net1592;
 wire net1591;
 wire net1593;
 wire _05623_;
 wire net1596;
 wire net1595;
 wire net1598;
 wire _05627_;
 wire _05628_;
 wire net1594;
 wire net1590;
 wire net2089;
 wire net2092;
 wire _05633_;
 wire _05634_;
 wire net2152;
 wire net1508;
 wire net2158;
 wire net1485;
 wire net1484;
 wire net1482;
 wire net1477;
 wire net1475;
 wire net1473;
 wire net1470;
 wire net1469;
 wire net1467;
 wire net1465;
 wire _05663_;
 wire _05664_;
 wire _05675_;
 wire _05679_;
 wire _05681_;
 wire _05685_;
 wire _05689_;
 wire _05693_;
 wire _05698_;
 wire _05702_;
 wire _05706_;
 wire _05711_;
 wire _05715_;
 wire _05719_;
 wire _05723_;
 wire _05727_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05835_;
 wire _05837_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05867_;
 wire _05868_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05874_;
 wire _05875_;
 wire _05877_;
 wire _05879_;
 wire _05880_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05888_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _06000_;
 wire _06001_;
 wire _06003_;
 wire _06004_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06460_;
 wire net154;
 wire net153;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire net152;
 wire net151;
 wire net150;
 wire _06473_;
 wire net149;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire net148;
 wire net147;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire net146;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire net145;
 wire net144;
 wire _06492_;
 wire net143;
 wire net142;
 wire net141;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire net140;
 wire _06502_;
 wire net139;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire net138;
 wire net137;
 wire net136;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire net135;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire net134;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire net133;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire net132;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire net131;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire net130;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire net129;
 wire net128;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire net127;
 wire net126;
 wire _06683_;
 wire _06684_;
 wire net125;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire net124;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire net123;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire net122;
 wire _06719_;
 wire net121;
 wire net120;
 wire _06722_;
 wire _06723_;
 wire net119;
 wire net118;
 wire _06726_;
 wire net117;
 wire _06728_;
 wire net116;
 wire net115;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire net114;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire net113;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire net112;
 wire _06840_;
 wire _06841_;
 wire net111;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire net110;
 wire _06856_;
 wire _06857_;
 wire net109;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire net108;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire net107;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire _06911_;
 wire net97;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire net96;
 wire net95;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire net94;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire net93;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire net92;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire net91;
 wire net90;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire net89;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire net88;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire net87;
 wire _07003_;
 wire _07004_;
 wire net86;
 wire net85;
 wire _07007_;
 wire _07008_;
 wire net84;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire net83;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire net82;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire net81;
 wire _07035_;
 wire _07036_;
 wire net80;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire net79;
 wire net78;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire net77;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire net76;
 wire net75;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire net66;
 wire _07089_;
 wire net65;
 wire net64;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire net63;
 wire _07104_;
 wire _07105_;
 wire net62;
 wire _07107_;
 wire _07108_;
 wire net61;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire net60;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire net59;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire net58;
 wire _07138_;
 wire net57;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire net56;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire net55;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire net54;
 wire net53;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire net52;
 wire _07407_;
 wire net51;
 wire net50;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire net49;
 wire net48;
 wire _07421_;
 wire _07422_;
 wire net47;
 wire net46;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire net45;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire net44;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire net43;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire net42;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire net1738;
 wire net1737;
 wire _07521_;
 wire net2015;
 wire _07523_;
 wire net2016;
 wire net2017;
 wire net1736;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire net2018;
 wire net1735;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire clknet_leaf_24_clk_i_regs;
 wire _07537_;
 wire clknet_leaf_25_clk_i_regs;
 wire _07539_;
 wire net1734;
 wire net1733;
 wire net1732;
 wire _07543_;
 wire _07544_;
 wire net1731;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire net1730;
 wire _07557_;
 wire net1729;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire net1728;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire net1727;
 wire _07570_;
 wire _07571_;
 wire net1726;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire net1724;
 wire _07579_;
 wire net1723;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire net1722;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire net1721;
 wire _07612_;
 wire _07613_;
 wire net1720;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire net1719;
 wire _07622_;
 wire net1718;
 wire _07624_;
 wire net1725;
 wire net1717;
 wire net1740;
 wire clknet_leaf_26_clk_i_regs;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire net1716;
 wire _07640_;
 wire net1714;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire net1712;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire net1711;
 wire net1713;
 wire net1715;
 wire net1710;
 wire net1709;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire net1708;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire net1707;
 wire _07676_;
 wire _07677_;
 wire net1706;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire net1705;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire clknet_leaf_27_clk_i_regs;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire net1702;
 wire net1701;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire net1700;
 wire _07710_;
 wire _07711_;
 wire clknet_leaf_28_clk_i_regs;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire clknet_leaf_29_clk_i_regs;
 wire _07718_;
 wire _07719_;
 wire net1699;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire net1698;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire net1697;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire net1696;
 wire net1695;
 wire _07745_;
 wire clknet_leaf_31_clk_i_regs;
 wire _07747_;
 wire _07748_;
 wire clknet_leaf_33_clk_i_regs;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire clknet_leaf_32_clk_i_regs;
 wire _07763_;
 wire clknet_0_clk_i_regs;
 wire _07765_;
 wire net1694;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire clknet_2_1__leaf_clk_i_regs;
 wire _07777_;
 wire _07778_;
 wire clknet_2_2__leaf_clk_i_regs;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire clknet_2_3__leaf_clk_i_regs;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire net1692;
 wire _07789_;
 wire net1691;
 wire net1690;
 wire _07792_;
 wire _07793_;
 wire clknet_leaf_0_clk;
 wire net1689;
 wire net1688;
 wire net1687;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire clknet_leaf_1_clk;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire net2481;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire net1685;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire net1684;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire clknet_leaf_3_clk;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire net1681;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire clknet_leaf_6_clk;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire net1678;
 wire _07999_;
 wire _08000_;
 wire net1677;
 wire clknet_leaf_7_clk;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire net1675;
 wire clknet_leaf_10_clk;
 wire net1674;
 wire net1673;
 wire _08015_;
 wire net1672;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire clknet_leaf_11_clk;
 wire net1670;
 wire _08022_;
 wire net1671;
 wire net1668;
 wire _08025_;
 wire _08026_;
 wire net1666;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire net1663;
 wire _08043_;
 wire net1662;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire net1658;
 wire net1659;
 wire net1657;
 wire _08054_;
 wire net1654;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire net1655;
 wire _08060_;
 wire net1652;
 wire _08062_;
 wire net1649;
 wire net1648;
 wire _08065_;
 wire net1647;
 wire _08067_;
 wire net1646;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire net1650;
 wire _08077_;
 wire net1644;
 wire net1642;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire net1641;
 wire _08085_;
 wire _08086_;
 wire net1640;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire net1643;
 wire _08101_;
 wire net1639;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire net1645;
 wire _08187_;
 wire net1651;
 wire net1638;
 wire net1637;
 wire _08191_;
 wire _08192_;
 wire net1636;
 wire _08194_;
 wire net1635;
 wire _08196_;
 wire _08197_;
 wire net1653;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire net1634;
 wire net1631;
 wire net1632;
 wire _08224_;
 wire net1630;
 wire net1633;
 wire _08227_;
 wire _08228_;
 wire net1629;
 wire net1656;
 wire net1627;
 wire net1625;
 wire _08233_;
 wire _08234_;
 wire net1626;
 wire net1624;
 wire _08237_;
 wire _08238_;
 wire net1628;
 wire _08240_;
 wire _08241_;
 wire net1622;
 wire _08243_;
 wire net1623;
 wire net1620;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire net1621;
 wire net1619;
 wire net1618;
 wire _08256_;
 wire _08257_;
 wire net1617;
 wire _08259_;
 wire _08260_;
 wire net1616;
 wire net1613;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire net1612;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire net1611;
 wire net1610;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire net1614;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire net1615;
 wire net1664;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire net1665;
 wire _08300_;
 wire net1608;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire net1667;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire net1609;
 wire net1606;
 wire net1602;
 wire _08321_;
 wire _08322_;
 wire net1600;
 wire _08324_;
 wire net1601;
 wire _08326_;
 wire _08327_;
 wire net1597;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire net1589;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire net1588;
 wire _08341_;
 wire net1587;
 wire net1586;
 wire _08344_;
 wire net1599;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire net1603;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire net1604;
 wire net1605;
 wire net1607;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire net1669;
 wire _08430_;
 wire net1585;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire _08434_;
 wire net1583;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire net1584;
 wire net1582;
 wire net1581;
 wire net1739;
 wire net1580;
 wire net1579;
 wire net1578;
 wire clknet_leaf_14_clk;
 wire _08518_;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire _08521_;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire _08525_;
 wire _08526_;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire net1575;
 wire net1576;
 wire _08531_;
 wire net1577;
 wire net1568;
 wire _08534_;
 wire _08535_;
 wire net1567;
 wire net1566;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire net1569;
 wire _08544_;
 wire net1570;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire net1564;
 wire net1565;
 wire net1571;
 wire net1563;
 wire net1562;
 wire net1572;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire net1573;
 wire net1574;
 wire clknet_leaf_22_clk;
 wire _08566_;
 wire clknet_leaf_23_clk;
 wire _08568_;
 wire clknet_leaf_24_clk;
 wire _08570_;
 wire _08571_;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire net1561;
 wire _08578_;
 wire net1560;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire net1559;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire net1558;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire net1557;
 wire net1556;
 wire _08632_;
 wire _08633_;
 wire clknet_leaf_27_clk;
 wire net1555;
 wire _08636_;
 wire _08637_;
 wire clknet_leaf_28_clk;
 wire net1554;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire net1553;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire net1552;
 wire _08659_;
 wire _08660_;
 wire clknet_leaf_30_clk;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire clknet_leaf_29_clk;
 wire net1551;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire clknet_leaf_31_clk;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire clknet_leaf_32_clk;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire net1550;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire clknet_leaf_33_clk;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire clknet_leaf_34_clk;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire clknet_leaf_35_clk;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire clknet_leaf_36_clk;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire clknet_leaf_37_clk;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire net1549;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire net1547;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire net1546;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire net1545;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire net1544;
 wire net1548;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire net1543;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire clknet_leaf_38_clk;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire clknet_0_clk;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire net1542;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire net1541;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire net1540;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire clknet_2_1_0_clk;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire clknet_2_2_0_clk;
 wire _09660_;
 wire clknet_2_3_0_clk;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire delaynet_0_core_clock;
 wire delaynet_1_core_clock;
 wire _09668_;
 wire delaynet_2_core_clock;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire delaynet_3_core_clock;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire delaynet_4_core_clock;
 wire net1539;
 wire net2051;
 wire net2052;
 wire net2053;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire net2054;
 wire _09702_;
 wire net2055;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire net2056;
 wire net2057;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire net2058;
 wire _09753_;
 wire net2059;
 wire _09755_;
 wire net2060;
 wire net1538;
 wire _09758_;
 wire net1537;
 wire _09760_;
 wire net2061;
 wire net2062;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire net2063;
 wire _09768_;
 wire net2064;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire net2065;
 wire _09774_;
 wire net2066;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire net2068;
 wire _09786_;
 wire _09787_;
 wire net2067;
 wire _09789_;
 wire net2069;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire net2070;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire net2071;
 wire net2072;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire net2073;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire net2074;
 wire _09809_;
 wire _09810_;
 wire net2075;
 wire net2076;
 wire _09813_;
 wire _09814_;
 wire net2077;
 wire _09816_;
 wire _09817_;
 wire net1536;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire net1535;
 wire _09823_;
 wire _09824_;
 wire net1534;
 wire _09826_;
 wire _09827_;
 wire net1533;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire net2078;
 wire _09834_;
 wire _09835_;
 wire net2079;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire net2080;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire net2081;
 wire _09848_;
 wire _09849_;
 wire net2082;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire net2083;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire net2084;
 wire _09861_;
 wire net2085;
 wire net2086;
 wire _09864_;
 wire net2087;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire net2088;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire net1532;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire net2090;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire net1531;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire net2091;
 wire _09957_;
 wire net1530;
 wire net2093;
 wire net2094;
 wire _09961_;
 wire _09962_;
 wire net1529;
 wire net2095;
 wire _09965_;
 wire net1528;
 wire net2096;
 wire net1527;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire net1526;
 wire net2097;
 wire net1525;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire net1524;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire net1523;
 wire _10014_;
 wire net1522;
 wire _10016_;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire net2103;
 wire net2104;
 wire net1521;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire net1520;
 wire _10037_;
 wire net2107;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire net2105;
 wire net2106;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire net2113;
 wire net2108;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire net2111;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire net2110;
 wire net2109;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire net2114;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire net2116;
 wire net2115;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire net2117;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire net2118;
 wire net2119;
 wire net1517;
 wire net1516;
 wire _10138_;
 wire _10139_;
 wire net2120;
 wire _10141_;
 wire net2121;
 wire net2122;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire net2123;
 wire net2124;
 wire _10152_;
 wire net2125;
 wire _10154_;
 wire _10155_;
 wire net2126;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire net2127;
 wire _10161_;
 wire _10162_;
 wire net2128;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire net2130;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire net2129;
 wire net2132;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire net2131;
 wire net2135;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire net1515;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire net2134;
 wire _10203_;
 wire net2133;
 wire net2136;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire net2138;
 wire _10211_;
 wire net2137;
 wire net1514;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire net1513;
 wire _10218_;
 wire _10219_;
 wire net2139;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire net1512;
 wire _10230_;
 wire _10231_;
 wire net2140;
 wire net2141;
 wire _10234_;
 wire net2142;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire net2143;
 wire net2145;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire net2144;
 wire _10247_;
 wire net2146;
 wire net2147;
 wire net2149;
 wire net2148;
 wire _10252_;
 wire _10253_;
 wire net1511;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire net2150;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire net1510;
 wire net1509;
 wire _10271_;
 wire net2151;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire net1507;
 wire net1505;
 wire net1504;
 wire _10279_;
 wire _10280_;
 wire net1502;
 wire _10282_;
 wire _10283_;
 wire net1501;
 wire net1503;
 wire net1500;
 wire _10287_;
 wire net1506;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire net2153;
 wire net2154;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire net2155;
 wire _10374_;
 wire net2156;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire net2157;
 wire net1499;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net2159;
 wire net1497;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire net1496;
 wire net1494;
 wire net1495;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire net1493;
 wire net1492;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire net1491;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire net1490;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire net2160;
 wire net1498;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire net1489;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire net2161;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire net1488;
 wire net1487;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire net1486;
 wire net1480;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire net1478;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire net1476;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire net1474;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire net1472;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire net1463;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire net1461;
 wire _10855_;
 wire net1460;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire net1459;
 wire _10861_;
 wire _10862_;
 wire net1458;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire net1457;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire net1462;
 wire _10958_;
 wire net1456;
 wire net1455;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire net1464;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire net1466;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire net1746;
 wire \alu_adder_result_ex[0] ;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire \alu_adder_result_ex[1] ;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net37;
 wire net9;
 wire net8;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire net155;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit_q[0] ;
 wire \cs_registers_i.mcountinhibit_q[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter_val_o[9] ;
 wire \cs_registers_i.mhpmcounter[1856] ;
 wire \cs_registers_i.mhpmcounter[1857] ;
 wire \cs_registers_i.mhpmcounter[1858] ;
 wire \cs_registers_i.mhpmcounter[1859] ;
 wire \cs_registers_i.mhpmcounter[1860] ;
 wire \cs_registers_i.mhpmcounter[1861] ;
 wire \cs_registers_i.mhpmcounter[1862] ;
 wire \cs_registers_i.mhpmcounter[1863] ;
 wire \cs_registers_i.mhpmcounter[1864] ;
 wire \cs_registers_i.mhpmcounter[1865] ;
 wire \cs_registers_i.mhpmcounter[1866] ;
 wire \cs_registers_i.mhpmcounter[1867] ;
 wire \cs_registers_i.mhpmcounter[1868] ;
 wire \cs_registers_i.mhpmcounter[1869] ;
 wire \cs_registers_i.mhpmcounter[1870] ;
 wire \cs_registers_i.mhpmcounter[1871] ;
 wire \cs_registers_i.mhpmcounter[1872] ;
 wire \cs_registers_i.mhpmcounter[1873] ;
 wire \cs_registers_i.mhpmcounter[1874] ;
 wire \cs_registers_i.mhpmcounter[1875] ;
 wire \cs_registers_i.mhpmcounter[1876] ;
 wire \cs_registers_i.mhpmcounter[1877] ;
 wire \cs_registers_i.mhpmcounter[1878] ;
 wire \cs_registers_i.mhpmcounter[1879] ;
 wire \cs_registers_i.mhpmcounter[1880] ;
 wire \cs_registers_i.mhpmcounter[1881] ;
 wire \cs_registers_i.mhpmcounter[1882] ;
 wire \cs_registers_i.mhpmcounter[1883] ;
 wire \cs_registers_i.mhpmcounter[1884] ;
 wire \cs_registers_i.mhpmcounter[1885] ;
 wire \cs_registers_i.mhpmcounter[1886] ;
 wire \cs_registers_i.mhpmcounter[1887] ;
 wire \cs_registers_i.mhpmcounter[1888] ;
 wire \cs_registers_i.mhpmcounter[1889] ;
 wire \cs_registers_i.mhpmcounter[1890] ;
 wire \cs_registers_i.mhpmcounter[1891] ;
 wire \cs_registers_i.mhpmcounter[1892] ;
 wire \cs_registers_i.mhpmcounter[1893] ;
 wire \cs_registers_i.mhpmcounter[1894] ;
 wire \cs_registers_i.mhpmcounter[1895] ;
 wire \cs_registers_i.mhpmcounter[1896] ;
 wire \cs_registers_i.mhpmcounter[1897] ;
 wire \cs_registers_i.mhpmcounter[1898] ;
 wire \cs_registers_i.mhpmcounter[1899] ;
 wire \cs_registers_i.mhpmcounter[1900] ;
 wire \cs_registers_i.mhpmcounter[1901] ;
 wire \cs_registers_i.mhpmcounter[1902] ;
 wire \cs_registers_i.mhpmcounter[1903] ;
 wire \cs_registers_i.mhpmcounter[1904] ;
 wire \cs_registers_i.mhpmcounter[1905] ;
 wire \cs_registers_i.mhpmcounter[1906] ;
 wire \cs_registers_i.mhpmcounter[1907] ;
 wire \cs_registers_i.mhpmcounter[1908] ;
 wire \cs_registers_i.mhpmcounter[1909] ;
 wire \cs_registers_i.mhpmcounter[1910] ;
 wire \cs_registers_i.mhpmcounter[1911] ;
 wire \cs_registers_i.mhpmcounter[1912] ;
 wire \cs_registers_i.mhpmcounter[1913] ;
 wire \cs_registers_i.mhpmcounter[1914] ;
 wire \cs_registers_i.mhpmcounter[1915] ;
 wire \cs_registers_i.mhpmcounter[1916] ;
 wire \cs_registers_i.mhpmcounter[1917] ;
 wire \cs_registers_i.mhpmcounter[1918] ;
 wire \cs_registers_i.mhpmcounter[1919] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mstatus_q[2] ;
 wire \cs_registers_i.mstatus_q[3] ;
 wire \cs_registers_i.mstatus_q[4] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_mode_id_o[0] ;
 wire \cs_registers_i.priv_mode_id_o[1] ;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire \ex_block_i.alu_i.imd_val_q_i[0] ;
 wire \ex_block_i.alu_i.imd_val_q_i[10] ;
 wire \ex_block_i.alu_i.imd_val_q_i[11] ;
 wire \ex_block_i.alu_i.imd_val_q_i[12] ;
 wire \ex_block_i.alu_i.imd_val_q_i[13] ;
 wire \ex_block_i.alu_i.imd_val_q_i[14] ;
 wire \ex_block_i.alu_i.imd_val_q_i[15] ;
 wire \ex_block_i.alu_i.imd_val_q_i[16] ;
 wire \ex_block_i.alu_i.imd_val_q_i[17] ;
 wire \ex_block_i.alu_i.imd_val_q_i[18] ;
 wire \ex_block_i.alu_i.imd_val_q_i[19] ;
 wire \ex_block_i.alu_i.imd_val_q_i[1] ;
 wire \ex_block_i.alu_i.imd_val_q_i[20] ;
 wire \ex_block_i.alu_i.imd_val_q_i[21] ;
 wire \ex_block_i.alu_i.imd_val_q_i[22] ;
 wire \ex_block_i.alu_i.imd_val_q_i[23] ;
 wire \ex_block_i.alu_i.imd_val_q_i[24] ;
 wire \ex_block_i.alu_i.imd_val_q_i[25] ;
 wire \ex_block_i.alu_i.imd_val_q_i[26] ;
 wire \ex_block_i.alu_i.imd_val_q_i[27] ;
 wire \ex_block_i.alu_i.imd_val_q_i[28] ;
 wire \ex_block_i.alu_i.imd_val_q_i[29] ;
 wire \ex_block_i.alu_i.imd_val_q_i[2] ;
 wire \ex_block_i.alu_i.imd_val_q_i[30] ;
 wire \ex_block_i.alu_i.imd_val_q_i[31] ;
 wire \ex_block_i.alu_i.imd_val_q_i[32] ;
 wire \ex_block_i.alu_i.imd_val_q_i[33] ;
 wire \ex_block_i.alu_i.imd_val_q_i[34] ;
 wire \ex_block_i.alu_i.imd_val_q_i[35] ;
 wire \ex_block_i.alu_i.imd_val_q_i[36] ;
 wire \ex_block_i.alu_i.imd_val_q_i[37] ;
 wire \ex_block_i.alu_i.imd_val_q_i[38] ;
 wire \ex_block_i.alu_i.imd_val_q_i[39] ;
 wire \ex_block_i.alu_i.imd_val_q_i[3] ;
 wire \ex_block_i.alu_i.imd_val_q_i[40] ;
 wire \ex_block_i.alu_i.imd_val_q_i[41] ;
 wire \ex_block_i.alu_i.imd_val_q_i[42] ;
 wire \ex_block_i.alu_i.imd_val_q_i[43] ;
 wire \ex_block_i.alu_i.imd_val_q_i[44] ;
 wire \ex_block_i.alu_i.imd_val_q_i[45] ;
 wire \ex_block_i.alu_i.imd_val_q_i[46] ;
 wire \ex_block_i.alu_i.imd_val_q_i[47] ;
 wire \ex_block_i.alu_i.imd_val_q_i[48] ;
 wire \ex_block_i.alu_i.imd_val_q_i[49] ;
 wire \ex_block_i.alu_i.imd_val_q_i[4] ;
 wire \ex_block_i.alu_i.imd_val_q_i[50] ;
 wire \ex_block_i.alu_i.imd_val_q_i[51] ;
 wire \ex_block_i.alu_i.imd_val_q_i[52] ;
 wire \ex_block_i.alu_i.imd_val_q_i[53] ;
 wire \ex_block_i.alu_i.imd_val_q_i[54] ;
 wire \ex_block_i.alu_i.imd_val_q_i[55] ;
 wire \ex_block_i.alu_i.imd_val_q_i[56] ;
 wire \ex_block_i.alu_i.imd_val_q_i[57] ;
 wire \ex_block_i.alu_i.imd_val_q_i[58] ;
 wire \ex_block_i.alu_i.imd_val_q_i[59] ;
 wire \ex_block_i.alu_i.imd_val_q_i[5] ;
 wire \ex_block_i.alu_i.imd_val_q_i[60] ;
 wire \ex_block_i.alu_i.imd_val_q_i[61] ;
 wire \ex_block_i.alu_i.imd_val_q_i[62] ;
 wire \ex_block_i.alu_i.imd_val_q_i[63] ;
 wire \ex_block_i.alu_i.imd_val_q_i[6] ;
 wire \ex_block_i.alu_i.imd_val_q_i[7] ;
 wire \ex_block_i.alu_i.imd_val_q_i[8] ;
 wire \ex_block_i.alu_i.imd_val_q_i[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_i ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_i ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[0] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[1] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[2] ;
 wire \load_store_unit_i.rdata_q[3] ;
 wire \load_store_unit_i.rdata_q[4] ;
 wire \load_store_unit_i.rdata_q[5] ;
 wire \load_store_unit_i.rdata_q[6] ;
 wire \load_store_unit_i.rdata_q[7] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net7;
 wire net6;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1747;
 wire net1748;
 wire net1786;
 wire net1750;
 wire net1751;
 wire net1780;
 wire net1765;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1787;
 wire net1794;
 wire net1792;
 wire net1790;
 wire net1788;
 wire net1789;
 wire net1791;
 wire net1793;
 wire net1795;
 wire net2007;
 wire net1813;
 wire net1796;
 wire net1797;
 wire net1812;
 wire net1798;
 wire net1799;
 wire net1808;
 wire net1800;
 wire net1803;
 wire net1801;
 wire net1802;
 wire net1804;
 wire net1806;
 wire net1807;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net2006;
 wire net1815;
 wire net1814;
 wire net2005;
 wire net2004;
 wire net2003;
 wire net1821;
 wire net1818;
 wire net1817;
 wire net1816;
 wire net1819;
 wire net1820;
 wire net2002;
 wire net2001;
 wire net2000;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1999;
 wire net1827;
 wire net1998;
 wire net1829;
 wire net1828;
 wire net1837;
 wire net1830;
 wire net1836;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1997;
 wire net1838;
 wire net1988;
 wire net1839;
 wire net1987;
 wire net1840;
 wire net1986;
 wire net1841;
 wire net1844;
 wire net1843;
 wire net1842;
 wire net1985;
 wire net1983;
 wire net1982;
 wire net1851;
 wire net1981;
 wire net1852;
 wire net1984;
 wire net1845;
 wire net1850;
 wire net1849;
 wire net1846;
 wire net1848;
 wire net1847;
 wire net1957;
 wire net1854;
 wire net1853;
 wire net1956;
 wire net1955;
 wire net1930;
 wire net1929;
 wire net1928;
 wire net1927;
 wire net1857;
 wire net1856;
 wire net1855;
 wire net1925;
 wire net1859;
 wire net1858;
 wire net1924;
 wire net1883;
 wire net1884;
 wire net1860;
 wire net1862;
 wire net1861;
 wire net1882;
 wire net1881;
 wire net1879;
 wire net1875;
 wire net1874;
 wire net1880;
 wire net1873;
 wire net1872;
 wire net1867;
 wire net1866;
 wire net1865;
 wire net1864;
 wire net1871;
 wire net1868;
 wire net1870;
 wire net1869;
 wire net1876;
 wire net1877;
 wire net1923;
 wire net1917;
 wire net1916;
 wire net1915;
 wire net1914;
 wire net1913;
 wire net1886;
 wire net1885;
 wire net1922;
 wire net1921;
 wire net1920;
 wire net1919;
 wire net1918;
 wire net1887;
 wire net1902;
 wire net1888;
 wire net1901;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1905;
 wire net1904;
 wire net1903;
 wire net1912;
 wire net1906;
 wire net1911;
 wire net1910;
 wire net1907;
 wire net1909;
 wire net1908;
 wire net1931;
 wire net1953;
 wire net1947;
 wire net1946;
 wire net1936;
 wire net1932;
 wire net1935;
 wire net1934;
 wire net1933;
 wire net1945;
 wire net1944;
 wire net1943;
 wire net1942;
 wire net1941;
 wire net1940;
 wire net1937;
 wire net1939;
 wire net1938;
 wire net1952;
 wire net1951;
 wire net1950;
 wire net1949;
 wire net1948;
 wire net1961;
 wire net1971;
 wire net1970;
 wire net1969;
 wire net1968;
 wire net1979;
 wire net1978;
 wire net1977;
 wire net1976;
 wire net1975;
 wire net1967;
 wire net1963;
 wire net1962;
 wire net1966;
 wire net1965;
 wire net1964;
 wire net1996;
 wire net1991;
 wire net1990;
 wire net1989;
 wire net1995;
 wire net1994;
 wire net1993;
 wire net1992;
 wire net2044;
 wire net2037;
 wire net2036;
 wire net2035;
 wire net2022;
 wire net2019;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_0_clk_i_regs;
 wire clknet_1_0__leaf_clk_i;
 wire net2046;
 wire clknet_0_clk_i;
 wire clk_i_regs;
 wire net2050;
 wire net2049;
 wire net2048;
 wire net2047;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire clknet_leaf_13_clk_i_regs;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire clknet_leaf_10_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire clknet_leaf_7_clk_i_regs;
 wire clknet_leaf_6_clk_i_regs;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_19_clk_i_regs;
 wire clknet_leaf_18_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_17_clk_i_regs;
 wire net2024;
 wire net2025;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2043;
 wire net2041;
 wire net2040;
 wire net2039;
 wire net2038;
 wire net1362;
 wire net1368;
 wire net1373;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11641_ (.I(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2010 (.I(net2193),
    .Z(net2009));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place2011 (.I(net2008),
    .Z(net2010));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2012 (.I(net2008),
    .Z(net2011));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2013 (.I(net2008),
    .Z(net2012));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2014 (.I(net2008),
    .Z(net2013));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place2015 (.I(net2005),
    .Z(net2014));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11648_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07516_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11649_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07517_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _11650_ (.I(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .ZN(_07518_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1739 (.I(_08034_),
    .Z(net1738));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1738 (.I(_08191_),
    .Z(net1737));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11653_ (.I0(_07516_),
    .I1(_07517_),
    .S(net1884),
    .Z(_07521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2016 (.I(net2005),
    .Z(net2015));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11655_ (.A1(net1958),
    .A2(net1959),
    .ZN(_07523_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place2017 (.I(net2015),
    .Z(net2016));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2018 (.I(net2005),
    .Z(net2017));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1737 (.I(_08448_),
    .Z(net1736));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11659_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07527_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11660_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07528_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11661_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11662_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net2001),
    .Z(_07530_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2019 (.I(net2005),
    .Z(net2018));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1736 (.I(_08486_),
    .Z(net1735));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11665_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A2(net2001),
    .Z(_07533_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11666_ (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .ZN(_07534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11667_ (.I0(_07530_),
    .I1(_07533_),
    .S(net1873),
    .Z(_07535_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_24_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11669_ (.I(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .ZN(_07537_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_25_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11671_ (.I0(_07527_),
    .I1(_07528_),
    .I2(_07529_),
    .I3(_07535_),
    .S0(net1884),
    .S1(net1867),
    .Z(_07539_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1735 (.I(_08606_),
    .Z(net1734));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1734 (.I(_08669_),
    .Z(net1733));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1733 (.I(_08810_),
    .Z(net1732));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11675_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07543_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11676_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_07544_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1732 (.I(_08870_),
    .Z(net1731));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11678_ (.I0(_07543_),
    .I1(_07544_),
    .S(net1884),
    .Z(_07546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11679_ (.A1(net1958),
    .A2(net1867),
    .ZN(_07547_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11680_ (.A1(_07546_),
    .A2(_07547_),
    .Z(_07548_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11681_ (.A1(_07521_),
    .A2(_07523_),
    .B1(_07539_),
    .B2(net1958),
    .C(_07548_),
    .ZN(_07549_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11682_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_07550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11683_ (.A1(net2081),
    .A2(_07550_),
    .ZN(_07551_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11684_ (.I(\load_store_unit_i.ls_fsm_cs[0] ),
    .ZN(_07552_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11685_ (.I(\load_store_unit_i.ls_fsm_cs[2] ),
    .ZN(_07553_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11686_ (.A1(_07552_),
    .A2(\load_store_unit_i.handle_misaligned_q ),
    .B(net2086),
    .C(_07553_),
    .ZN(_07554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11687_ (.A1(_07551_),
    .A2(_07554_),
    .ZN(_07555_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1731 (.I(_08906_),
    .Z(net1730));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11689_ (.I(net1889),
    .ZN(_07557_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1730 (.I(_08945_),
    .Z(net1729));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11691_ (.A1(net2144),
    .A2(_07557_),
    .Z(_07559_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11692_ (.I(net2133),
    .ZN(_07560_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11693_ (.A1(net1888),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_07561_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1729 (.I(_08962_),
    .Z(net1728));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11695_ (.A1(net1888),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .ZN(_07563_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11696_ (.A1(_07560_),
    .A2(_07561_),
    .B(_07563_),
    .ZN(_07564_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11697_ (.A1(_07559_),
    .A2(_07564_),
    .Z(_07565_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11698_ (.I(\id_stage_i.controller_i.instr_i[6] ),
    .ZN(_07566_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11699_ (.I(net2144),
    .ZN(_07567_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11700_ (.A1(_07566_),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .B(_07567_),
    .ZN(_07568_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1728 (.I(_08999_),
    .Z(net1727));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11702_ (.A1(net2147),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .ZN(_07570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11703_ (.A1(net1889),
    .A2(_07570_),
    .ZN(_07571_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1727 (.I(_09059_),
    .Z(net1726));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11705_ (.A1(_07568_),
    .A2(_07571_),
    .B(net2130),
    .ZN(_07573_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11706_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .ZN(_07574_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11707_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .A3(net1893),
    .ZN(_07575_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11708_ (.A1(_07560_),
    .A2(net1889),
    .A3(_07561_),
    .A4(_07575_),
    .Z(_07576_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11709_ (.A1(_07565_),
    .A2(_07573_),
    .B1(_07574_),
    .B2(_07576_),
    .ZN(_07577_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1725 (.I(_09095_),
    .Z(net1724));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 _11711_ (.I(net2019),
    .ZN(_07579_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1724 (.I(_09148_),
    .Z(net1723));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11713_ (.I(\id_stage_i.controller_i.instr_i[5] ),
    .ZN(_07581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11714_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .ZN(_07582_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _11715_ (.A1(net1893),
    .A2(net1890),
    .Z(_07583_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11716_ (.A1(_07581_),
    .A2(_07582_),
    .A3(_07583_),
    .Z(_07584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11717_ (.A1(net1888),
    .A2(net1889),
    .ZN(_07585_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11718_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .Z(_07586_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _11719_ (.A1(_07579_),
    .A2(_07584_),
    .A3(_07585_),
    .B(_07586_),
    .ZN(_07587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11720_ (.A1(net2130),
    .A2(_07570_),
    .Z(_07588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11721_ (.A1(_07559_),
    .A2(_07588_),
    .Z(_07589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11722_ (.A1(net1888),
    .A2(\id_stage_i.controller_i.instr_i[5] ),
    .Z(_07590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11723_ (.A1(_07557_),
    .A2(_07590_),
    .ZN(_07591_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11724_ (.A1(_07568_),
    .A2(_07591_),
    .B(net2132),
    .ZN(_07592_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11725_ (.A1(\id_stage_i.controller_i.instr_i[0] ),
    .A2(\id_stage_i.controller_i.instr_i[1] ),
    .A3(net1893),
    .Z(_07593_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11726_ (.A1(net2132),
    .A2(_07557_),
    .A3(_07570_),
    .A4(_07593_),
    .Z(_07594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11727_ (.I(\id_stage_i.controller_i.instr_i[12] ),
    .ZN(_07595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11728_ (.A1(_07595_),
    .A2(_07574_),
    .ZN(_07596_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11729_ (.A1(_07594_),
    .A2(net1831),
    .ZN(_07597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11730_ (.A1(_07560_),
    .A2(_07586_),
    .Z(_07598_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11731_ (.I(\id_stage_i.id_fsm_q ),
    .ZN(_07599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11732_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_07599_),
    .B(net2170),
    .C(_07563_),
    .ZN(_07600_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11733_ (.A1(_07598_),
    .A2(net2183),
    .ZN(_07601_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11734_ (.A1(_07589_),
    .A2(_07592_),
    .B(_07597_),
    .C(_07601_),
    .ZN(_07602_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11735_ (.A1(_07602_),
    .A2(_07577_),
    .A3(_07587_),
    .A4(net1817),
    .Z(_07603_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1723 (.I(_09182_),
    .Z(net1722));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11737_ (.A1(_07559_),
    .A2(_07564_),
    .ZN(_07605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11738_ (.A1(net2147),
    .A2(_07581_),
    .B(net2144),
    .ZN(_07606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11739_ (.A1(net2170),
    .A2(net2149),
    .Z(_07607_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11740_ (.A1(_07606_),
    .A2(_07607_),
    .B(_07560_),
    .ZN(_07608_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11741_ (.A1(_07574_),
    .A2(_07576_),
    .B(_07551_),
    .C(_07554_),
    .ZN(_07609_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11742_ (.A1(_07605_),
    .A2(_07608_),
    .B(_07609_),
    .C(_07587_),
    .ZN(_07610_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1722 (.I(_09239_),
    .Z(net1721));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11744_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(net2064),
    .ZN(_07612_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11745_ (.A1(_07598_),
    .A2(net2183),
    .Z(_07613_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1721 (.I(_09276_),
    .Z(net1720));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11747_ (.A1(\id_stage_i.controller_i.instr_i[2] ),
    .A2(\id_stage_i.controller_i.instr_i[3] ),
    .ZN(_07615_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11748_ (.A1(\id_stage_i.controller_i.instr_i[5] ),
    .A2(_07586_),
    .A3(_07615_),
    .Z(_07616_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11749_ (.A1(_07579_),
    .A2(_07585_),
    .ZN(_07617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11750_ (.A1(_07616_),
    .A2(_07617_),
    .B(_07582_),
    .ZN(_07618_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11751_ (.A1(_07589_),
    .A2(_07592_),
    .B(_07597_),
    .C(_07618_),
    .ZN(_07619_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11752_ (.A1(_07551_),
    .A2(_07554_),
    .Z(_07620_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1720 (.I(_09443_),
    .Z(net1719));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11754_ (.A1(_07619_),
    .A2(_07613_),
    .B(net1816),
    .ZN(_07622_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1719 (.I(_09665_),
    .Z(net1718));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11756_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net1818),
    .ZN(_07624_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _11757_ (.A1(net1803),
    .A2(net2126),
    .B1(_07612_),
    .B2(net1741),
    .C(_07624_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11758_ (.I(net1704),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1726 (.I(net1724),
    .Z(net1725));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1718 (.I(_09671_),
    .Z(net1717));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_26_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11763_ (.A1(net1889),
    .A2(net1888),
    .A3(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_07629_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11764_ (.A1(_07629_),
    .A2(_07582_),
    .A3(_07583_),
    .A4(_07581_),
    .Z(_07630_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11765_ (.A1(net2130),
    .A2(_07557_),
    .A3(_07570_),
    .Z(_07631_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11766_ (.A1(net2021),
    .A2(_07574_),
    .Z(_07632_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _11767_ (.A1(_07631_),
    .A2(_07632_),
    .B(_07600_),
    .ZN(_07633_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11768_ (.A1(net2130),
    .A2(net2147),
    .A3(_07557_),
    .Z(_07634_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11769_ (.A1(_07630_),
    .A2(_07634_),
    .Z(_07635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _11770_ (.A1(_07575_),
    .A2(net2110),
    .B1(_07635_),
    .B2(_07633_),
    .C(net2115),
    .ZN(_07636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11771_ (.I0(net1932),
    .I1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .S(net2069),
    .Z(_07637_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11772_ (.A1(_07560_),
    .A2(net2170),
    .A3(_07561_),
    .Z(_07638_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1717 (.I(_09689_),
    .Z(net1716));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11774_ (.A1(net2021),
    .A2(_07574_),
    .ZN(_07640_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1715 (.I(_09780_),
    .Z(net1714));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11776_ (.I(\id_stage_i.controller_i.instr_valid_i ),
    .ZN(_07642_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11777_ (.A1(_07642_),
    .A2(\id_stage_i.id_fsm_q ),
    .B(_07590_),
    .C(_07557_),
    .ZN(_07643_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _11778_ (.A1(_07640_),
    .A2(_07638_),
    .B(_07643_),
    .ZN(_07644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11779_ (.A1(_07557_),
    .A2(_07590_),
    .Z(_07645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11780_ (.A1(net2130),
    .A2(_07593_),
    .A3(_07645_),
    .Z(_07646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _11781_ (.A1(_07593_),
    .A2(_07644_),
    .B(_07646_),
    .C(net1817),
    .ZN(_07647_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11782_ (.A1(_07616_),
    .A2(_07585_),
    .A3(net2117),
    .ZN(_07648_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11783_ (.A1(net2144),
    .A2(_07566_),
    .A3(net1889),
    .Z(_07649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11784_ (.A1(net2081),
    .A2(_07550_),
    .Z(_07650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1713 (.I(_09831_),
    .Z(net1712));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11786_ (.I(net2086),
    .ZN(_07652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11787_ (.A1(net2099),
    .A2(_01354_),
    .B(_07652_),
    .C(net2081),
    .ZN(_07653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11788_ (.A1(_07598_),
    .A2(_07649_),
    .B(_07653_),
    .C(_07650_),
    .ZN(_07654_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11789_ (.A1(_07648_),
    .A2(net2181),
    .Z(_07655_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11790_ (.A1(net2061),
    .A2(_07655_),
    .Z(_07656_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11791_ (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .ZN(_07657_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1712 (.I(_09851_),
    .Z(net1711));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1714 (.I(_09805_),
    .Z(net1713));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1716 (.I(net1714),
    .Z(net1715));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1711 (.I(_09861_),
    .Z(net1710));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1710 (.I(_09878_),
    .Z(net1709));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11797_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .S0(net2168),
    .S1(net1903),
    .Z(_07663_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11798_ (.A1(net1860),
    .A2(net1901),
    .A3(net2104),
    .A4(_07663_),
    .Z(_07664_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11799_ (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .ZN(_07665_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11800_ (.I(net2155),
    .ZN(_07666_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1709 (.I(_09946_),
    .Z(net1708));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11802_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S0(net2168),
    .S1(net1903),
    .Z(_07668_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11803_ (.A1(net1899),
    .A2(net1858),
    .A3(net1856),
    .A4(_07668_),
    .Z(_07669_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11804_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07670_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11805_ (.A1(net1899),
    .A2(net1858),
    .A3(net2104),
    .A4(_07670_),
    .Z(_07671_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11806_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07672_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11807_ (.A1(net1860),
    .A2(net1901),
    .A3(net1856),
    .A4(_07672_),
    .Z(_07673_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11808_ (.A1(_07664_),
    .A2(_07669_),
    .A3(_07671_),
    .A4(_07673_),
    .Z(_07674_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1708 (.I(_03988_),
    .Z(net1707));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11810_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .S(net2078),
    .Z(_07676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11811_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(net2078),
    .Z(_07677_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1707 (.I(_03992_),
    .Z(net1706));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11813_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A2(net2078),
    .Z(_07679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11814_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net2078),
    .Z(_07680_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11815_ (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .ZN(_07681_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1706 (.I(_00947_),
    .Z(net1705));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11817_ (.I0(_07676_),
    .I1(_07677_),
    .I2(_07679_),
    .I3(_07680_),
    .S0(net2104),
    .S1(net1847),
    .Z(_07683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11818_ (.A1(net1861),
    .A2(net1859),
    .ZN(_07684_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11819_ (.A1(_07683_),
    .A2(net1830),
    .Z(_07685_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11820_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11821_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11822_ (.I0(_07686_),
    .I1(_07687_),
    .S(net1856),
    .Z(_07688_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11823_ (.A1(net1899),
    .A2(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .ZN(_07689_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11824_ (.A1(_07688_),
    .A2(_07689_),
    .Z(_07690_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11825_ (.A1(_07674_),
    .A2(_07685_),
    .A3(_07690_),
    .Z(_07691_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _11826_ (.A1(_07616_),
    .A2(_07585_),
    .A3(_07643_),
    .A4(net2117),
    .ZN(_07692_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _11827_ (.A1(net2483),
    .A2(_07692_),
    .ZN(_07693_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11828_ (.A1(_07637_),
    .A2(_07656_),
    .B1(net1798),
    .B2(net1797),
    .ZN(_07694_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _11829_ (.I(_07694_),
    .ZN(_07695_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1705 (.I(_01226_),
    .Z(net1704));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1704 (.I(_07694_),
    .Z(net1703));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_27_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11833_ (.A1(_07575_),
    .A2(net2110),
    .B1(_07633_),
    .B2(_07635_),
    .ZN(_07697_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11834_ (.A1(_07560_),
    .A2(_07575_),
    .A3(_07591_),
    .Z(_07698_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _11835_ (.A1(_07575_),
    .A2(_07633_),
    .B(_07698_),
    .C(net1816),
    .ZN(_07699_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11836_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_07697_),
    .A3(_07699_),
    .Z(_07700_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1703 (.I(net2299),
    .Z(net1702));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1702 (.I(net2118),
    .Z(net1701));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _11840_ (.A1(_07584_),
    .A2(net2117),
    .ZN(_07704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11841_ (.A1(_07630_),
    .A2(_07634_),
    .ZN(_07705_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _11842_ (.A1(_07593_),
    .A2(_07704_),
    .B1(_07644_),
    .B2(_07705_),
    .C(_07620_),
    .ZN(_07706_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11843_ (.A1(net1908),
    .A2(_07706_),
    .Z(_07707_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11844_ (.A1(_07700_),
    .A2(_07707_),
    .B(_07655_),
    .ZN(_07708_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1701 (.I(_01173_),
    .Z(net1700));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11846_ (.A1(net1816),
    .A2(_07692_),
    .Z(_07710_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11847_ (.A1(_07586_),
    .A2(_07615_),
    .Z(_07711_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_28_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11849_ (.A1(_07711_),
    .A2(net2183),
    .ZN(_07713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11850_ (.A1(_07654_),
    .A2(_07713_),
    .Z(_07714_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _11851_ (.A1(_07714_),
    .A2(_07636_),
    .ZN(_07715_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _11852_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A2(net2061),
    .A3(_07710_),
    .A4(_07715_),
    .ZN(_07716_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_29_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11854_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07718_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11855_ (.A1(net1860),
    .A2(net1901),
    .A3(net2104),
    .A4(_07718_),
    .Z(_07719_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1700 (.I(_07925_),
    .Z(net1699));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11857_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07721_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11858_ (.A1(net1899),
    .A2(net1858),
    .A3(net1856),
    .A4(_07721_),
    .Z(_07722_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11859_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07723_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11860_ (.A1(net1899),
    .A2(net1858),
    .A3(net2104),
    .A4(_07723_),
    .Z(_07724_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11861_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07725_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11862_ (.A1(net1860),
    .A2(net1901),
    .A3(net1856),
    .A4(_07725_),
    .Z(_07726_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _11863_ (.A1(_07719_),
    .A2(_07722_),
    .A3(_07724_),
    .A4(_07726_),
    .Z(_07727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11864_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .S(net2168),
    .Z(_07728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11865_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(net2168),
    .Z(_07729_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1699 (.I(_07946_),
    .Z(net1698));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11867_ (.A1(net2078),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .Z(_07731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11868_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net2168),
    .Z(_07732_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11869_ (.I0(_07728_),
    .I1(_07729_),
    .I2(_07731_),
    .I3(_07732_),
    .S0(net2104),
    .S1(net1847),
    .Z(_07733_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11870_ (.A1(net1830),
    .A2(_07733_),
    .Z(_07734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1698 (.I(_01208_),
    .Z(net1697));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net2168),
    .S1(net1903),
    .Z(_07736_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11873_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .S0(net1906),
    .S1(net1903),
    .Z(_07737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11874_ (.I0(_07736_),
    .I1(_07737_),
    .S(net1856),
    .Z(_07738_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11875_ (.A1(_07689_),
    .A2(_07738_),
    .Z(_07739_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11876_ (.A1(_07727_),
    .A2(_07734_),
    .A3(_07739_),
    .Z(_07740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11877_ (.A1(_07693_),
    .A2(net1796),
    .ZN(_07741_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _11878_ (.A1(_07708_),
    .A2(_07716_),
    .A3(_07741_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _11879_ (.I(_01135_),
    .ZN(_07742_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_30_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_30_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1697 (.I(_07996_),
    .Z(net1696));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1696 (.I(_01214_),
    .Z(net1695));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _11883_ (.A1(_07666_),
    .A2(net2184),
    .Z(_07745_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_31_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_31_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11885_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net1909),
    .Z(_07747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _11886_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A2(_07745_),
    .B1(_07747_),
    .B2(net2104),
    .ZN(_07748_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_33_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_33_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S0(net1931),
    .S1(net1909),
    .Z(_07750_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11889_ (.A1(net1903),
    .A2(_07750_),
    .ZN(_07751_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11890_ (.A1(net1903),
    .A2(_07748_),
    .B(_07751_),
    .ZN(_07752_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net1909),
    .S1(net1903),
    .Z(_07753_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11892_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .S0(net1909),
    .S1(net1903),
    .Z(_07754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11893_ (.I0(_07753_),
    .I1(_07754_),
    .S(net1856),
    .Z(_07755_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11894_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S0(net2152),
    .S1(net1909),
    .Z(_07756_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11895_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S0(net2152),
    .S1(net1909),
    .Z(_07757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11896_ (.I0(_07756_),
    .I1(_07757_),
    .S(net1847),
    .Z(_07758_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11897_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net1909),
    .S1(net1903),
    .Z(_07759_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11898_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .S0(net1909),
    .S1(net1903),
    .Z(_07760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11899_ (.I0(_07759_),
    .I1(_07760_),
    .S(net1856),
    .Z(_07761_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_32_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11901_ (.I0(_07752_),
    .I1(_07755_),
    .I2(_07758_),
    .I3(_07761_),
    .S0(net1901),
    .S1(net1899),
    .Z(_07763_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk_i_regs (.I(clk_i_regs),
    .Z(clknet_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _11903_ (.I(net1740),
    .ZN(_07765_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1695 (.I(_08185_),
    .Z(net1694));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11905_ (.A1(_07654_),
    .A2(_07713_),
    .ZN(_07767_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11906_ (.A1(net1848),
    .A2(net1800),
    .A3(_07767_),
    .Z(_07768_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11907_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_07706_),
    .A3(net1799),
    .A4(_07767_),
    .Z(_07769_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _11908_ (.A1(_07710_),
    .A2(_07768_),
    .A3(_07769_),
    .Z(_07770_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _11909_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(net2061),
    .A3(_07715_),
    .ZN(_07771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11910_ (.A1(net1797),
    .A2(_07765_),
    .B1(_07770_),
    .B2(_07771_),
    .ZN(_07772_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11911_ (.I(net1611),
    .ZN(_07773_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_0__f_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_2_0__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1694 (.I(_08218_),
    .Z(net1693));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11914_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A2(net1799),
    .Z(_07774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11915_ (.A1(_07648_),
    .A2(net2181),
    .ZN(_07775_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_1__f_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_2_1__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11917_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net1918),
    .S1(net1905),
    .Z(_07777_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11918_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .S0(net1918),
    .S1(net1905),
    .Z(_07778_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_2__f_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_2_2__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11920_ (.I0(_07777_),
    .I1(_07778_),
    .S(net1853),
    .Z(_07780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11921_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .S(net2184),
    .Z(_07781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11922_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net1916),
    .Z(_07782_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_3__f_clk_i_regs (.I(clknet_0_clk_i_regs),
    .Z(clknet_2_3__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11924_ (.A1(net1916),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .Z(_07784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11925_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net1916),
    .Z(_07785_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11926_ (.I0(_07781_),
    .I1(_07782_),
    .I2(_07784_),
    .I3(_07785_),
    .S0(net1957),
    .S1(net1847),
    .Z(_07786_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_4 _11927_ (.A1(_07689_),
    .A2(_07780_),
    .B1(_07786_),
    .B2(_07684_),
    .ZN(_07787_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1693 (.I(_01172_),
    .Z(net1692));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11929_ (.A1(_07657_),
    .A2(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .ZN(_07789_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1692 (.I(_01179_),
    .Z(net1691));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1691 (.I(_01186_),
    .Z(net1690));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11932_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net1927),
    .S1(net1905),
    .Z(_07792_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _11933_ (.A1(net1853),
    .A2(_07789_),
    .A3(_07792_),
    .ZN(_07793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload0 (.I(clknet_2_0__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1690 (.I(_01200_),
    .Z(net1689));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1689 (.I(_01207_),
    .Z(net1688));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1688 (.I(_08544_),
    .Z(net1687));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11938_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .S0(net1927),
    .S1(net1905),
    .Z(_07798_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _11939_ (.A1(net1860),
    .A2(net1900),
    .A3(net1939),
    .A4(_07798_),
    .ZN(_07799_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11940_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .S0(net1927),
    .S1(net1905),
    .Z(_07800_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11941_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net1927),
    .S1(net1905),
    .Z(_07801_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11942_ (.A1(_07657_),
    .A2(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .A3(_07666_),
    .Z(_07802_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _11943_ (.A1(net1939),
    .A2(_07789_),
    .A3(_07800_),
    .B1(_07801_),
    .B2(_07802_),
    .ZN(_07803_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _11944_ (.A1(_07803_),
    .A2(_07793_),
    .A3(_07799_),
    .A4(_07787_),
    .Z(_07804_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _11945_ (.A1(net2483),
    .A2(_07692_),
    .Z(_07805_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload1 (.I(clknet_2_1__leaf_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _11947_ (.A1(net1858),
    .A2(_07697_),
    .A3(_07775_),
    .B1(_07804_),
    .B2(_07805_),
    .ZN(_07807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11948_ (.A1(net2066),
    .A2(_07774_),
    .B(_07807_),
    .ZN(_07808_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_leaf_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _11950_ (.I(net1702),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11951_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(net1799),
    .Z(_07809_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11952_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S0(net2152),
    .S1(net2078),
    .Z(_07810_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11953_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S0(net2152),
    .S1(net2078),
    .Z(_07811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11954_ (.I0(_07810_),
    .I1(_07811_),
    .S(net1847),
    .Z(_07812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .S(net1909),
    .Z(_07813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11956_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(net1909),
    .Z(_07814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11957_ (.A1(net1909),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .Z(_07815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net1909),
    .Z(_07816_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11959_ (.I0(_07813_),
    .I1(_07814_),
    .I2(_07815_),
    .I3(_07816_),
    .S0(net2142),
    .S1(net1847),
    .Z(_07817_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _11960_ (.A1(_07689_),
    .A2(_07812_),
    .B1(_07817_),
    .B2(_07684_),
    .ZN(_07818_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S0(net2089),
    .S1(net1903),
    .Z(_07819_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone2482 (.I(_09844_),
    .Z(net2481));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11963_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S0(net1933),
    .S1(net1909),
    .Z(_07821_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11964_ (.A1(net1899),
    .A2(net1859),
    .A3(net1903),
    .A4(_07821_),
    .Z(_07822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _11965_ (.A1(_07802_),
    .A2(_07819_),
    .B(_07822_),
    .ZN(_07823_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1686 (.I(_01235_),
    .Z(net1685));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11967_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S0(net2142),
    .S1(net2089),
    .Z(_07825_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11968_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .S0(net1909),
    .S1(net1903),
    .Z(_07826_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _11969_ (.A1(net1861),
    .A2(net1902),
    .A3(net1934),
    .A4(_07826_),
    .Z(_07827_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _11970_ (.A1(net1847),
    .A2(_07789_),
    .A3(_07825_),
    .B(_07827_),
    .ZN(_07828_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _11971_ (.A1(_07818_),
    .A2(_07823_),
    .A3(_07828_),
    .Z(_07829_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _11972_ (.A1(net1860),
    .A2(_07697_),
    .A3(_07775_),
    .B1(net1794),
    .B2(_07805_),
    .ZN(_07830_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _11973_ (.A1(net2066),
    .A2(_07809_),
    .B(_07830_),
    .ZN(_07831_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1685 (.I(_01242_),
    .Z(net1684));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1684 (.I(_01249_),
    .Z(net1683));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11976_ (.I(net1701),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _11977_ (.I(\id_stage_i.controller_i.instr_i[25] ),
    .ZN(_07833_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11978_ (.A1(_07638_),
    .A2(_07640_),
    .B(_07634_),
    .C(_07643_),
    .ZN(_07834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _11979_ (.A1(_07593_),
    .A2(_07834_),
    .B(_07704_),
    .C(net1817),
    .ZN(_07835_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _11980_ (.A1(net1799),
    .A2(_07655_),
    .B1(_07835_),
    .B2(_07805_),
    .ZN(_07836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net1907),
    .Z(_07837_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload3 (.I(clknet_leaf_25_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _11983_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .A2(net1828),
    .B1(_07837_),
    .B2(net2112),
    .C(net1904),
    .ZN(_07839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _11984_ (.A1(net1904),
    .A2(net1935),
    .ZN(_07840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11985_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(net1907),
    .Z(_07841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11986_ (.A1(_07657_),
    .A2(_07665_),
    .Z(_07842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11987_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .S(net1907),
    .Z(_07843_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _11988_ (.A1(net1934),
    .A2(net1847),
    .A3(_07843_),
    .Z(_07844_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _11989_ (.A1(_07840_),
    .A2(_07841_),
    .B(_07842_),
    .C(_07844_),
    .ZN(_07845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _11990_ (.A1(net1860),
    .A2(net1900),
    .Z(_07846_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11991_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net1907),
    .S1(net1903),
    .Z(_07847_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11992_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S0(net1907),
    .S1(net1903),
    .Z(_07848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _11993_ (.I0(_07847_),
    .I1(_07848_),
    .S(net1857),
    .Z(_07849_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _11994_ (.A1(_07846_),
    .A2(_07849_),
    .ZN(_07850_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11995_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net2184),
    .S1(net2101),
    .Z(_07851_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11996_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .S0(net2184),
    .S1(net2101),
    .Z(_07852_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11997_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net2184),
    .S1(net2101),
    .Z(_07853_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11998_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .S0(net2184),
    .S1(net2101),
    .Z(_07854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _11999_ (.I0(_07851_),
    .I1(_07852_),
    .I2(_07853_),
    .I3(_07854_),
    .S0(net1857),
    .S1(net1859),
    .Z(_07855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12000_ (.A1(net1899),
    .A2(_07855_),
    .ZN(_07856_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12001_ (.A1(_07839_),
    .A2(_07845_),
    .B(_07850_),
    .C(_07856_),
    .ZN(_07857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12002_ (.A1(net1797),
    .A2(net1792),
    .ZN(_07858_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12003_ (.A1(_07833_),
    .A2(_07836_),
    .B(_07858_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12004_ (.I(net1700),
    .ZN(_07859_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1683 (.I(_01263_),
    .Z(net1682));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12006_ (.I(net1897),
    .ZN(_07860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12007_ (.A1(net1799),
    .A2(_07714_),
    .B(_07835_),
    .ZN(_07861_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12008_ (.A1(net1899),
    .A2(net1901),
    .Z(_07862_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12009_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net2168),
    .S1(net1903),
    .Z(_07863_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12010_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S0(net2168),
    .S1(net1903),
    .Z(_07864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12011_ (.I0(_07863_),
    .I1(_07864_),
    .S(net1857),
    .Z(_07865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12012_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S0(net2151),
    .S1(net2078),
    .Z(_07866_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12013_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S0(net2151),
    .S1(net2078),
    .Z(_07867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12014_ (.I0(_07866_),
    .I1(_07867_),
    .S(net1847),
    .Z(_07868_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12015_ (.A1(net1899),
    .A2(net1858),
    .Z(_07869_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12016_ (.A1(_07862_),
    .A2(_07865_),
    .B1(_07868_),
    .B2(_07869_),
    .ZN(_07870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12017_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .S(net2168),
    .Z(_07871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12018_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S(net2168),
    .Z(_07872_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12019_ (.A1(net2078),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .Z(_07873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12020_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net2168),
    .Z(_07874_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12021_ (.I0(_07871_),
    .I1(_07872_),
    .I2(_07873_),
    .I3(_07874_),
    .S0(net2104),
    .S1(net1847),
    .Z(_07875_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12022_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07876_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12023_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07877_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12024_ (.I0(_07876_),
    .I1(_07877_),
    .S(net1857),
    .Z(_07878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12025_ (.A1(net1827),
    .A2(_07875_),
    .B1(_07878_),
    .B2(_07846_),
    .ZN(_07879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12026_ (.A1(_07870_),
    .A2(_07879_),
    .ZN(_07880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12027_ (.A1(net1797),
    .A2(net1790),
    .ZN(_07881_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _12028_ (.A1(_07860_),
    .A2(net1797),
    .A3(_07861_),
    .B(_07881_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12029_ (.I(_01180_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1682 (.I(_01270_),
    .Z(net1681));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12031_ (.A1(net1816),
    .A2(_07692_),
    .ZN(_07883_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12032_ (.A1(_07699_),
    .A2(_07775_),
    .B1(_07883_),
    .B2(_07697_),
    .ZN(_07884_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12033_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07885_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12034_ (.A1(net1860),
    .A2(net1900),
    .A3(net1936),
    .A4(_07885_),
    .Z(_07886_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12035_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07887_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12036_ (.A1(net1899),
    .A2(net1859),
    .A3(net1854),
    .A4(_07887_),
    .Z(_07888_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12037_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07889_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12038_ (.A1(net1899),
    .A2(net1859),
    .A3(net1936),
    .A4(_07889_),
    .Z(_07890_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12039_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07891_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12040_ (.A1(net1860),
    .A2(net1900),
    .A3(net1854),
    .A4(_07891_),
    .Z(_07892_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12041_ (.A1(_07886_),
    .A2(_07888_),
    .A3(_07890_),
    .A4(_07892_),
    .Z(_07893_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12042_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07894_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12043_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_07895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12044_ (.I0(_07894_),
    .I1(_07895_),
    .S(net1854),
    .Z(_07896_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12045_ (.A1(net1846),
    .A2(_07896_),
    .Z(_07897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12046_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .S(net1914),
    .Z(_07898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12047_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(net1914),
    .Z(_07899_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12048_ (.A1(net1914),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .Z(_07900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12049_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net1914),
    .Z(_07901_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12050_ (.I0(_07898_),
    .I1(_07899_),
    .I2(_07900_),
    .I3(_07901_),
    .S0(net1936),
    .S1(net1848),
    .Z(_07902_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12051_ (.A1(_07684_),
    .A2(_07902_),
    .Z(_07903_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12052_ (.A1(_07893_),
    .A2(_07897_),
    .A3(_07903_),
    .Z(_07904_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _12053_ (.A1(net1896),
    .A2(_07884_),
    .B1(net1797),
    .B2(net1788),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12054_ (.I(net1895),
    .ZN(_07905_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12055_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07906_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12056_ (.A1(net1860),
    .A2(net1900),
    .A3(net2112),
    .A4(_07906_),
    .Z(_07907_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12057_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07908_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12058_ (.A1(net1853),
    .A2(_07789_),
    .A3(_07908_),
    .Z(_07909_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12059_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07910_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12060_ (.A1(net1939),
    .A2(_07789_),
    .A3(_07910_),
    .Z(_07911_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12061_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07912_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12062_ (.A1(_07802_),
    .A2(_07912_),
    .Z(_07913_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12063_ (.A1(_07907_),
    .A2(_07909_),
    .A3(_07911_),
    .A4(_07913_),
    .Z(_07914_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12064_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07915_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12065_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .S0(net1922),
    .S1(net1905),
    .Z(_07916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12066_ (.I0(_07915_),
    .I1(_07916_),
    .S(net1854),
    .Z(_07917_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12067_ (.A1(net1846),
    .A2(_07917_),
    .Z(_07918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12068_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net1922),
    .Z(_07919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12069_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A2(net1829),
    .B1(_07919_),
    .B2(net1936),
    .ZN(_07920_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12070_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net1936),
    .S1(net1922),
    .Z(_07921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12071_ (.A1(net1905),
    .A2(_07921_),
    .ZN(_07922_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12072_ (.A1(net1905),
    .A2(_07920_),
    .B(_07922_),
    .C(_07842_),
    .ZN(_07923_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12073_ (.A1(_07914_),
    .A2(_07918_),
    .A3(_07923_),
    .ZN(_07924_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12074_ (.A1(_07905_),
    .A2(_07836_),
    .B1(_07924_),
    .B2(net1795),
    .ZN(_07925_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload4 (.I(clknet_leaf_27_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12076_ (.I(net1699),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12077_ (.I(net1894),
    .ZN(_07926_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12078_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .S0(net2089),
    .S1(net1903),
    .Z(_07927_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12079_ (.A1(net1862),
    .A2(net1902),
    .A3(net2114),
    .A4(_07927_),
    .Z(_07928_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12080_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S0(net1912),
    .S1(net1903),
    .Z(_07929_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12081_ (.A1(net1856),
    .A2(_07789_),
    .A3(_07929_),
    .Z(_07930_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12082_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S0(net1912),
    .S1(net1903),
    .Z(_07931_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12083_ (.A1(net2114),
    .A2(_07789_),
    .A3(_07931_),
    .Z(_07932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12084_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S0(net2089),
    .S1(net1903),
    .Z(_07933_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12085_ (.A1(_07802_),
    .A2(_07933_),
    .Z(_07934_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12086_ (.A1(_07928_),
    .A2(_07930_),
    .A3(_07932_),
    .A4(_07934_),
    .Z(_07935_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12087_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net1910),
    .S1(net1903),
    .Z(_07936_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12088_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S0(net1910),
    .S1(net1903),
    .Z(_07937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12089_ (.I0(_07936_),
    .I1(_07937_),
    .S(net1856),
    .Z(_07938_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12090_ (.A1(_07689_),
    .A2(_07938_),
    .Z(_07939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12091_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net1912),
    .Z(_07940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12092_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .A2(net1829),
    .B1(_07940_),
    .B2(net1945),
    .ZN(_07941_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12093_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net1945),
    .S1(net1912),
    .Z(_07942_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12094_ (.A1(net1903),
    .A2(_07942_),
    .ZN(_07943_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12095_ (.A1(net1903),
    .A2(_07941_),
    .B(_07943_),
    .C(_07842_),
    .ZN(_07944_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12096_ (.A1(_07935_),
    .A2(_07939_),
    .A3(_07944_),
    .ZN(_07945_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12097_ (.A1(_07926_),
    .A2(_07836_),
    .B1(_07945_),
    .B2(net1795),
    .ZN(_07946_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload5 (.I(clknet_leaf_29_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12099_ (.I(net1698),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _12100_ (.I(net1892),
    .ZN(_07947_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload6 (.I(clknet_leaf_30_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12102_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .S0(net1912),
    .S1(net1905),
    .Z(_07949_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12103_ (.A1(net1862),
    .A2(net1902),
    .A3(net1951),
    .A4(_07949_),
    .Z(_07950_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12104_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S0(net1915),
    .S1(net1905),
    .Z(_07951_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12105_ (.A1(net1853),
    .A2(_07789_),
    .A3(_07951_),
    .Z(_07952_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12106_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S0(net1915),
    .S1(net1905),
    .Z(_07953_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12107_ (.A1(net1951),
    .A2(_07789_),
    .A3(_07953_),
    .Z(_07954_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12108_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S0(net1912),
    .S1(net1905),
    .Z(_07955_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12109_ (.A1(_07802_),
    .A2(_07955_),
    .Z(_07956_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12110_ (.A1(_07950_),
    .A2(_07952_),
    .A3(_07954_),
    .A4(_07956_),
    .Z(_07957_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12111_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net1917),
    .S1(net1905),
    .Z(_07958_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12112_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .S0(net1917),
    .S1(net1905),
    .Z(_07959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12113_ (.I0(_07958_),
    .I1(_07959_),
    .S(net1853),
    .Z(_07960_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12114_ (.A1(net1846),
    .A2(_07960_),
    .Z(_07961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12115_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net2179),
    .Z(_07962_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12116_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A2(net1829),
    .B1(_07962_),
    .B2(net1957),
    .ZN(_07963_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12117_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net1957),
    .S1(net1915),
    .Z(_07964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12118_ (.A1(net1905),
    .A2(_07964_),
    .ZN(_07965_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12119_ (.A1(net1905),
    .A2(_07963_),
    .B(_07965_),
    .C(_07842_),
    .ZN(_07966_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12120_ (.A1(_07957_),
    .A2(_07961_),
    .A3(_07966_),
    .ZN(_07967_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12121_ (.A1(net1845),
    .A2(_07836_),
    .B1(_07967_),
    .B2(net1795),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12122_ (.I(net1697),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12123_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .ZN(_07968_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12124_ (.A1(net1891),
    .A2(net2181),
    .A3(_07713_),
    .ZN(_07969_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12125_ (.A1(_07968_),
    .A2(net2069),
    .A3(_07714_),
    .B(_07969_),
    .ZN(_07970_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12126_ (.A1(net2061),
    .A2(_07710_),
    .Z(_07971_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12127_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S0(net1931),
    .S1(net2078),
    .Z(_07972_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12128_ (.A1(net1903),
    .A2(_07972_),
    .Z(_07973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12129_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(net2078),
    .Z(_07974_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12130_ (.A1(_07840_),
    .A2(_07974_),
    .Z(_07975_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12131_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .S(net1906),
    .Z(_07976_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12132_ (.A1(net2104),
    .A2(net1847),
    .A3(_07976_),
    .Z(_07977_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12133_ (.A1(_07869_),
    .A2(_07973_),
    .A3(_07975_),
    .A4(_07977_),
    .Z(_07978_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12134_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07979_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12135_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .S0(net2078),
    .S1(net1903),
    .Z(_07980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12136_ (.I0(_07979_),
    .I1(_07980_),
    .S(net1857),
    .Z(_07981_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12137_ (.A1(_07862_),
    .A2(_07981_),
    .Z(_07982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12138_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .S(net1906),
    .Z(_07983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12139_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S(net1906),
    .Z(_07984_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12140_ (.A1(net2078),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .Z(_07985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12141_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net1906),
    .Z(_07986_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12142_ (.I0(_07983_),
    .I1(_07984_),
    .I2(_07985_),
    .I3(_07986_),
    .S0(net2151),
    .S1(net1847),
    .Z(_07987_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12143_ (.A1(net1827),
    .A2(_07987_),
    .Z(_07988_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12144_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .S0(net1931),
    .S1(net1903),
    .Z(_07989_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12145_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S0(net1931),
    .S1(net1903),
    .Z(_07990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12146_ (.I0(_07989_),
    .I1(_07990_),
    .S(net2078),
    .Z(_07991_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12147_ (.A1(_07846_),
    .A2(_07991_),
    .Z(_07992_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12148_ (.A1(_07982_),
    .A2(_07978_),
    .A3(_07988_),
    .A4(_07992_),
    .Z(_07993_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12149_ (.A1(net1932),
    .A2(net1816),
    .A3(_07692_),
    .Z(_07994_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12150_ (.A1(_07706_),
    .A2(_07699_),
    .A3(_07714_),
    .A4(_07994_),
    .Z(_07995_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12151_ (.A1(_07970_),
    .A2(_07971_),
    .B1(net1787),
    .B2(net1797),
    .C(_07995_),
    .ZN(_07996_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12152_ (.I(_07996_),
    .ZN(_07997_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1681 (.I(_01284_),
    .Z(net1680));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1680 (.I(_01291_),
    .Z(net1679));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1679 (.I(_01298_),
    .Z(net1678));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _12156_ (.A1(_07581_),
    .A2(_07582_),
    .A3(_07583_),
    .A4(_07585_),
    .ZN(_07999_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _12157_ (.I(net2020),
    .ZN(_08000_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1678 (.I(_01305_),
    .Z(net1677));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload7 (.I(clknet_leaf_32_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12160_ (.A1(net1958),
    .A2(net1959),
    .A3(net1962),
    .A4(net1975),
    .Z(_08003_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12161_ (.A1(net2005),
    .A2(_08003_),
    .Z(_08004_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12162_ (.A1(_08000_),
    .A2(_08004_),
    .Z(_08005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12163_ (.A1(net2021),
    .A2(net1826),
    .A3(_08005_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12164_ (.I(_00946_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload8 (.I(clknet_leaf_33_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload9 (.I(clknet_leaf_1_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12167_ (.A1(net2020),
    .A2(net1826),
    .A3(_08004_),
    .Z(_08008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12168_ (.I(_08008_),
    .ZN(_08009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1677 (.I(_01333_),
    .Z(net1676));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12170_ (.I(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .ZN(_08010_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1676 (.I(_01340_),
    .Z(net1675));
 gf180mcu_fd_sc_mcu9t5v0__inv_16 clkload10 (.I(clknet_leaf_2_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1675 (.I(_09674_),
    .Z(net1674));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1674 (.I(_09678_),
    .Z(net1673));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12175_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net2004),
    .S1(net1964),
    .Z(_08015_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1673 (.I(_09682_),
    .Z(net1672));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12177_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net2004),
    .S1(net1964),
    .Z(_08017_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12178_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S0(net2004),
    .S1(net1967),
    .Z(_08018_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12179_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S0(net2018),
    .S1(net1964),
    .Z(_08019_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload11 (.I(clknet_leaf_4_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1671 (.I(_09751_),
    .Z(net1670));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12182_ (.I0(_08015_),
    .I1(_08017_),
    .I2(_08018_),
    .I3(_08019_),
    .S0(_07518_),
    .S1(net1865),
    .Z(_08022_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1672 (.I(net1670),
    .Z(net1671));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1669 (.I(_09755_),
    .Z(net1668));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12185_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S0(net2018),
    .S1(net1964),
    .Z(_08025_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12186_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S0(net2018),
    .S1(net1964),
    .Z(_08026_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1667 (.I(_09768_),
    .Z(net1666));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12188_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net2018),
    .S1(net1964),
    .Z(_08028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12189_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net2018),
    .Z(_08029_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12190_ (.A1(net2018),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .Z(_08030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12191_ (.I0(_08029_),
    .I1(_08030_),
    .S(net1869),
    .Z(_08031_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12192_ (.I0(_08025_),
    .I1(_08026_),
    .I2(_08028_),
    .I3(_08031_),
    .S0(_07518_),
    .S1(net1865),
    .Z(_08032_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12193_ (.A1(net1958),
    .A2(_08032_),
    .Z(_08033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12194_ (.A1(net1842),
    .A2(_08022_),
    .B(_08033_),
    .ZN(_08034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12195_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(net2064),
    .ZN(_08035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12196_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net2483),
    .ZN(_08036_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12197_ (.A1(net2126),
    .A2(net1738),
    .B1(_08035_),
    .B2(net2052),
    .C(_08036_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12198_ (.I(net2159),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12199_ (.I(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .ZN(_08037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12200_ (.A1(_07559_),
    .A2(_07588_),
    .ZN(_08038_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12201_ (.A1(_07606_),
    .A2(_07645_),
    .B(_07560_),
    .ZN(_08039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12202_ (.A1(_08038_),
    .A2(_08039_),
    .B1(net1831),
    .B2(_07594_),
    .C(_07587_),
    .ZN(_08040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12203_ (.A1(_08040_),
    .A2(_07601_),
    .B(net1818),
    .ZN(_08041_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1664 (.I(_09772_),
    .Z(net1663));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12205_ (.A1(net1831),
    .A2(net1826),
    .Z(_08043_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1663 (.I(_09772_),
    .Z(net1662));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12207_ (.A1(net1965),
    .A2(_08043_),
    .Z(_08045_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12208_ (.A1(_07613_),
    .A2(_07619_),
    .B(_08045_),
    .C(net1816),
    .ZN(_08046_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12209_ (.A1(\id_stage_i.controller_i.instr_i[13] ),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_08047_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12210_ (.A1(_08047_),
    .A2(_07594_),
    .B(_07650_),
    .C(_07653_),
    .ZN(_08048_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12211_ (.A1(_07565_),
    .A2(_07573_),
    .B(_07618_),
    .C(_08048_),
    .ZN(_08049_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12212_ (.A1(_08037_),
    .A2(_08041_),
    .B(_08046_),
    .C(_08049_),
    .ZN(_08050_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1659 (.I(_09782_),
    .Z(net1658));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1660 (.I(_09776_),
    .Z(net1659));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1658 (.I(_09784_),
    .Z(net1657));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12216_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S0(net2137),
    .S1(net1964),
    .Z(_08054_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1655 (.I(_09787_),
    .Z(net1654));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12218_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S0(net2137),
    .S1(net1964),
    .Z(_08056_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12219_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S0(net2137),
    .S1(net1964),
    .Z(_08057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12220_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net2002),
    .Z(_08058_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1656 (.I(net1654),
    .Z(net1655));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12222_ (.A1(net2137),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .Z(_08060_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1653 (.I(_09792_),
    .Z(net1652));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12224_ (.I0(_08058_),
    .I1(_08060_),
    .S(net1869),
    .Z(_08062_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1650 (.I(_09794_),
    .Z(net1649));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1649 (.I(_09798_),
    .Z(net1648));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12227_ (.I0(_08054_),
    .I1(_08056_),
    .I2(_08057_),
    .I3(_08062_),
    .S0(_07518_),
    .S1(net1864),
    .Z(_08065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1648 (.I(net1646),
    .Z(net1647));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12229_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08067_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1647 (.I(_09803_),
    .Z(net1646));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12231_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08069_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12232_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08070_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12233_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08071_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12234_ (.I0(_08067_),
    .I1(_08069_),
    .I2(_08070_),
    .I3(_08071_),
    .S0(_07518_),
    .S1(net1864),
    .Z(_08072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12235_ (.A1(net1842),
    .A2(_08072_),
    .Z(_08073_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12236_ (.A1(net1958),
    .A2(_08065_),
    .B(_08073_),
    .ZN(_08074_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12237_ (.A1(_07613_),
    .A2(_07619_),
    .B(\cs_registers_i.pc_id_i[1] ),
    .C(net1816),
    .ZN(_08075_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1651 (.I(net1649),
    .Z(net1650));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12239_ (.A1(net2100),
    .A2(net1786),
    .B(_08075_),
    .C(net2063),
    .ZN(_08077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12240_ (.A1(_08050_),
    .A2(_08077_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12241_ (.I(_01145_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1645 (.I(_09807_),
    .Z(net1644));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1643 (.I(_09810_),
    .Z(net1642));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12244_ (.A1(net2007),
    .A2(_08049_),
    .A3(_08043_),
    .Z(_08080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12245_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(_08049_),
    .Z(_08081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12246_ (.I0(_08080_),
    .I1(_08081_),
    .S(_07622_),
    .Z(_08082_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _12247_ (.A1(net1818),
    .A2(_07577_),
    .A3(_07587_),
    .A4(_07602_),
    .ZN(_08083_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1642 (.I(_09814_),
    .Z(net1641));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12249_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08085_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12250_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08086_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1641 (.I(_09817_),
    .Z(net1640));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12252_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08088_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12253_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08089_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12254_ (.I0(_08085_),
    .I1(_08086_),
    .I2(_08088_),
    .I3(_08089_),
    .S0(_07518_),
    .S1(net1864),
    .Z(_08090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12255_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S0(net2137),
    .S1(net1964),
    .Z(_08091_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12256_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S0(net2002),
    .S1(net1964),
    .Z(_08092_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12257_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S0(net2137),
    .S1(net1964),
    .Z(_08093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12258_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net2002),
    .Z(_08094_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12259_ (.A1(net2137),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .Z(_08095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12260_ (.I0(_08094_),
    .I1(_08095_),
    .S(net1869),
    .Z(_08096_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12261_ (.I0(_08091_),
    .I1(_08092_),
    .I2(_08093_),
    .I3(_08096_),
    .S0(_07518_),
    .S1(net1864),
    .Z(_08097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12262_ (.I0(_08090_),
    .I1(_08097_),
    .S(net1842),
    .Z(_08098_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12263_ (.A1(_08083_),
    .A2(net1784),
    .Z(_08099_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12264_ (.A1(_08082_),
    .A2(_08099_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12265_ (.I(_01139_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1644 (.I(net1642),
    .Z(net1643));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12267_ (.A1(net2022),
    .A2(net2019),
    .A3(net1845),
    .Z(_08101_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1640 (.I(_09821_),
    .Z(net1639));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12269_ (.A1(_07595_),
    .A2(_07579_),
    .A3(net1892),
    .Z(_08103_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12270_ (.A1(_08101_),
    .A2(_08103_),
    .B(_08000_),
    .ZN(_08104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12271_ (.A1(net2020),
    .A2(_07595_),
    .ZN(_08105_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12272_ (.A1(net1892),
    .A2(_08105_),
    .Z(_08106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12273_ (.A1(_07566_),
    .A2(net2189),
    .Z(_08107_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12274_ (.A1(_07616_),
    .A2(_08107_),
    .ZN(_08108_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12275_ (.A1(net1894),
    .A2(net1895),
    .A3(net1891),
    .ZN(_08109_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12276_ (.A1(net1898),
    .A2(net1896),
    .A3(net1897),
    .ZN(_08110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12277_ (.A1(_08109_),
    .A2(_08110_),
    .ZN(_08111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12278_ (.A1(_08104_),
    .A2(_08106_),
    .B(_08108_),
    .C(_08111_),
    .ZN(_08112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12279_ (.A1(net2022),
    .A2(_07579_),
    .Z(_08113_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _12280_ (.A1(_07557_),
    .A2(\id_stage_i.controller_i.instr_valid_i ),
    .A3(_07599_),
    .A4(_07590_),
    .Z(_08114_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12281_ (.A1(_07711_),
    .A2(_08114_),
    .ZN(_08115_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _12282_ (.A1(net1896),
    .A2(net1894),
    .A3(net1895),
    .A4(net1891),
    .ZN(_08116_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12283_ (.A1(_08000_),
    .A2(net2021),
    .A3(net2019),
    .A4(_07947_),
    .Z(_08117_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12284_ (.A1(net2020),
    .A2(_07595_),
    .B1(_08116_),
    .B2(_08117_),
    .ZN(_08118_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12285_ (.A1(_07557_),
    .A2(_07561_),
    .A3(_07582_),
    .A4(_07583_),
    .Z(_08119_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _12286_ (.A1(net2020),
    .A2(_08113_),
    .A3(_08115_),
    .B1(_08118_),
    .B2(_08119_),
    .ZN(_08120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12287_ (.A1(_08000_),
    .A2(net2022),
    .Z(_08121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12288_ (.A1(_07566_),
    .A2(net1889),
    .ZN(_08122_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12289_ (.A1(net2019),
    .A2(_07947_),
    .B(_08109_),
    .C(_08110_),
    .ZN(_08123_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12290_ (.A1(net1896),
    .A2(net1894),
    .A3(net1895),
    .A4(net1891),
    .Z(_08124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12291_ (.A1(net2019),
    .A2(_08124_),
    .Z(_08125_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _12292_ (.A1(_07584_),
    .A2(_08122_),
    .A3(_08123_),
    .B1(_08125_),
    .B2(_08119_),
    .ZN(_08126_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12293_ (.A1(_07711_),
    .A2(_07632_),
    .A3(_08114_),
    .Z(_08127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12294_ (.A1(_08121_),
    .A2(_08126_),
    .B(_08127_),
    .ZN(_08128_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12295_ (.A1(_08112_),
    .A2(_08120_),
    .B(_08128_),
    .ZN(_08129_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12296_ (.A1(_07567_),
    .A2(net1889),
    .A3(_07590_),
    .Z(_08130_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12297_ (.A1(net2130),
    .A2(_07570_),
    .A3(_07574_),
    .Z(_08131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12298_ (.A1(net2146),
    .A2(_07581_),
    .B(net2130),
    .ZN(_08132_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12299_ (.A1(net2130),
    .A2(net2146),
    .B(net2189),
    .ZN(_08133_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12300_ (.A1(_07586_),
    .A2(_08133_),
    .Z(_08134_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12301_ (.A1(_08130_),
    .A2(_08131_),
    .B1(_08132_),
    .B2(net2144),
    .C(_08134_),
    .ZN(_08135_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12302_ (.A1(net2020),
    .A2(_07579_),
    .ZN(_08136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12303_ (.A1(net2021),
    .A2(net2019),
    .Z(_08137_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12304_ (.A1(_08000_),
    .A2(_08124_),
    .A3(_08137_),
    .ZN(_08138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12305_ (.A1(_08136_),
    .A2(_08138_),
    .B(_08119_),
    .ZN(_08139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12306_ (.A1(_08139_),
    .A2(_08135_),
    .Z(_08140_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12307_ (.A1(net2170),
    .A2(net2021),
    .A3(net2149),
    .Z(_08141_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12308_ (.A1(_08114_),
    .A2(_08141_),
    .B(net2020),
    .C(_07711_),
    .ZN(_08142_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12309_ (.A1(net2021),
    .A2(net2019),
    .ZN(_08143_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12310_ (.A1(_07711_),
    .A2(_08114_),
    .A3(_08143_),
    .ZN(_08144_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12311_ (.A1(net1845),
    .A2(_08109_),
    .A3(_08110_),
    .ZN(_08145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12312_ (.A1(net2020),
    .A2(_08137_),
    .ZN(_08146_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12313_ (.A1(_07584_),
    .A2(_08122_),
    .A3(_08145_),
    .A4(_08146_),
    .Z(_08147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12314_ (.A1(_08142_),
    .A2(_08144_),
    .A3(_08147_),
    .ZN(_08148_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12315_ (.A1(_08000_),
    .A2(_08124_),
    .ZN(_08149_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12316_ (.A1(_07595_),
    .A2(_07579_),
    .Z(_08150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12317_ (.A1(_08137_),
    .A2(_08149_),
    .B(_08150_),
    .C(_08119_),
    .ZN(_08151_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12318_ (.A1(_08000_),
    .A2(net2022),
    .ZN(_08152_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12319_ (.A1(_08000_),
    .A2(net2022),
    .A3(_07579_),
    .Z(_08153_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12320_ (.A1(_07711_),
    .A2(_08152_),
    .A3(_08114_),
    .A4(_08153_),
    .Z(_08154_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12321_ (.A1(_08135_),
    .A2(_08151_),
    .A3(_08154_),
    .Z(_08155_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12322_ (.A1(_07616_),
    .A2(_08107_),
    .Z(_08156_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12323_ (.A1(net1898),
    .A2(_07947_),
    .Z(_08157_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12324_ (.A1(net2020),
    .A2(net2021),
    .ZN(_08158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12325_ (.A1(_07579_),
    .A2(_07947_),
    .A3(_08158_),
    .Z(_08159_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _12326_ (.A1(_08000_),
    .A2(net2022),
    .A3(net2019),
    .A4(_07833_),
    .Z(_08160_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12327_ (.A1(\id_stage_i.controller_i.instr_i[29] ),
    .A2(\id_stage_i.controller_i.instr_i[28] ),
    .A3(\id_stage_i.controller_i.instr_i[31] ),
    .Z(_08161_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12328_ (.A1(net1896),
    .A2(net1897),
    .Z(_08162_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12329_ (.A1(_08161_),
    .A2(_08162_),
    .ZN(_08163_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12330_ (.A1(_08157_),
    .A2(_08159_),
    .A3(_08160_),
    .B(_08163_),
    .ZN(_08164_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12331_ (.A1(_07579_),
    .A2(net1892),
    .A3(_08158_),
    .Z(_08165_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12332_ (.A1(net2020),
    .A2(net1845),
    .A3(_08143_),
    .Z(_08166_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12333_ (.A1(_08109_),
    .A2(_08110_),
    .Z(_08167_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12334_ (.A1(_08165_),
    .A2(_08166_),
    .B(_08167_),
    .ZN(_08168_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12335_ (.A1(_08156_),
    .A2(_08164_),
    .A3(_08168_),
    .Z(_08169_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12336_ (.A1(_08155_),
    .A2(_08148_),
    .A3(_08140_),
    .A4(_08169_),
    .Z(_08170_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12337_ (.A1(net2019),
    .A2(_08105_),
    .A3(_08145_),
    .Z(_08171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12338_ (.A1(_07860_),
    .A2(_08171_),
    .B(_08108_),
    .ZN(_08172_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12339_ (.A1(_08157_),
    .A2(_08159_),
    .A3(_08160_),
    .Z(_08173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12340_ (.I0(_07579_),
    .I1(_08047_),
    .S(net2021),
    .Z(_08174_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12341_ (.A1(net2020),
    .A2(_07947_),
    .A3(_08143_),
    .ZN(_08175_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12342_ (.A1(_07579_),
    .A2(net1892),
    .A3(_08158_),
    .ZN(_08176_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12343_ (.A1(net1892),
    .A2(_08174_),
    .B(_08175_),
    .C(_08176_),
    .ZN(_08177_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12344_ (.A1(_08163_),
    .A2(_08173_),
    .B1(_08177_),
    .B2(_08167_),
    .C(_08108_),
    .ZN(_08178_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12345_ (.A1(_07711_),
    .A2(_08114_),
    .Z(_08179_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12346_ (.A1(\id_stage_i.controller_i.instr_i[27] ),
    .A2(\id_stage_i.controller_i.instr_i[26] ),
    .A3(\id_stage_i.controller_i.instr_i[30] ),
    .Z(_08180_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12347_ (.A1(_07833_),
    .A2(_08161_),
    .A3(_08180_),
    .ZN(_08181_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _12348_ (.A1(_07616_),
    .A2(_08107_),
    .A3(_08181_),
    .Z(_08182_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12349_ (.A1(_08179_),
    .A2(_08135_),
    .A3(_08139_),
    .A4(_08182_),
    .Z(_08183_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _12350_ (.A1(_08183_),
    .A2(_08178_),
    .A3(_08172_),
    .ZN(_08184_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12351_ (.A1(_08170_),
    .A2(_08129_),
    .B(_08184_),
    .ZN(_08185_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1646 (.I(_09807_),
    .Z(net1645));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12353_ (.I(net2111),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12354_ (.A1(_08156_),
    .A2(net1825),
    .ZN(_08187_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1652 (.I(_09794_),
    .Z(net1651));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1639 (.I(net1637),
    .Z(net1638));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1638 (.I(net1636),
    .Z(net1637));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12358_ (.I(net2092),
    .ZN(_08191_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12359_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .ZN(_08192_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1637 (.I(_09827_),
    .Z(net1636));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12361_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .ZN(_08194_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1636 (.I(_09832_),
    .Z(net1635));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12363_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .ZN(_08196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12364_ (.A1(_08194_),
    .A2(_08196_),
    .Z(_08197_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1654 (.I(_09792_),
    .Z(net1653));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12366_ (.A1(_08194_),
    .A2(_08196_),
    .ZN(_08199_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12367_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A3(_08199_),
    .Z(_08200_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12368_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .B2(_08197_),
    .C1(_08200_),
    .C2(net1798),
    .ZN(_08201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12369_ (.A1(net2028),
    .A2(net1737),
    .B(_08201_),
    .ZN(_08202_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12370_ (.A1(_08187_),
    .A2(_08202_),
    .Z(_08203_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12371_ (.A1(_07595_),
    .A2(_07579_),
    .A3(net1892),
    .Z(_08204_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12372_ (.A1(net2022),
    .A2(net2019),
    .A3(net1845),
    .Z(_08205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12373_ (.A1(_08204_),
    .A2(_08205_),
    .B(net2020),
    .ZN(_08206_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12374_ (.A1(net1892),
    .A2(_08105_),
    .ZN(_08207_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12375_ (.A1(_08206_),
    .A2(_08207_),
    .B(_08156_),
    .C(_08167_),
    .ZN(_08208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12376_ (.A1(_07607_),
    .A2(_07711_),
    .Z(_08209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12377_ (.A1(net2019),
    .A2(net1845),
    .ZN(_08210_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12378_ (.A1(_08152_),
    .A2(_08210_),
    .A3(_08124_),
    .B(_08105_),
    .ZN(_08211_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12379_ (.A1(net2020),
    .A2(_08113_),
    .ZN(_08212_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12380_ (.A1(_08209_),
    .A2(_08211_),
    .B1(_08212_),
    .B2(_08179_),
    .ZN(_08213_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12381_ (.A1(_08121_),
    .A2(_08126_),
    .Z(_08214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12382_ (.A1(_08208_),
    .A2(_08213_),
    .B(_08127_),
    .C(_08214_),
    .ZN(_08215_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12383_ (.A1(_08155_),
    .A2(_08148_),
    .A3(_08140_),
    .A4(_08169_),
    .ZN(_08216_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _12384_ (.A1(_08179_),
    .A2(_08140_),
    .A3(_08172_),
    .A4(_08178_),
    .Z(_08217_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12385_ (.A1(_08216_),
    .A2(_08215_),
    .B(_08217_),
    .ZN(_08218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12386_ (.I0(net1693),
    .I1(net1694),
    .S(_07695_),
    .Z(_08219_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12387_ (.A1(_08203_),
    .A2(_08219_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12388_ (.I(_00008_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12389_ (.A1(_01139_),
    .A2(_08187_),
    .Z(_08220_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1635 (.I(_09835_),
    .Z(net1634));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1632 (.I(_09841_),
    .Z(net1631));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1633 (.I(net1631),
    .Z(net1632));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12393_ (.A1(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .A2(net1814),
    .A3(net1823),
    .Z(_08224_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12394_ (.A1(_08220_),
    .A2(_08224_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12395_ (.I(_00814_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12396_ (.A1(_00010_),
    .A2(net2071),
    .ZN(\alu_adder_result_ex[1] ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12397_ (.I(\alu_adder_result_ex[1] ),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1631 (.I(_09844_),
    .Z(net1630));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1634 (.I(net1632),
    .Z(net1633));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12400_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .ZN(_08227_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12401_ (.A1(_08227_),
    .A2(_08192_),
    .A3(_08197_),
    .Z(_08228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1630 (.I(_09846_),
    .Z(net1629));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1657 (.I(_09787_),
    .Z(net1656));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1628 (.I(_09849_),
    .Z(net1627));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1626 (.I(_09853_),
    .Z(net1625));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12406_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08233_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12407_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1627 (.I(net1625),
    .Z(net1626));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1625 (.I(_09859_),
    .Z(net1624));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12410_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12411_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net1999),
    .Z(_08238_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1629 (.I(net1627),
    .Z(net1628));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12413_ (.A1(net1999),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .Z(_08240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12414_ (.I0(_08238_),
    .I1(_08240_),
    .S(net1872),
    .Z(_08241_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1623 (.I(_09871_),
    .Z(net1622));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12416_ (.I0(_08233_),
    .I1(_08234_),
    .I2(_08237_),
    .I3(_08241_),
    .S0(_07518_),
    .S1(net1867),
    .Z(_08243_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1624 (.I(_09871_),
    .Z(net1623));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1621 (.I(_09880_),
    .Z(net1620));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12419_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08246_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12420_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08247_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12421_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08248_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12422_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S0(net1999),
    .S1(net1964),
    .Z(_08249_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12423_ (.I0(_08246_),
    .I1(_08247_),
    .I2(_08248_),
    .I3(_08249_),
    .S0(_07518_),
    .S1(net1867),
    .Z(_08250_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12424_ (.A1(net1842),
    .A2(_08250_),
    .Z(_08251_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12425_ (.A1(net1958),
    .A2(_08243_),
    .B(_08251_),
    .ZN(_08252_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1622 (.I(net1620),
    .Z(net1621));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1620 (.I(_09891_),
    .Z(net1619));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1619 (.I(_09955_),
    .Z(net1618));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _12429_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .B2(net1824),
    .ZN(_08256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12430_ (.A1(_07765_),
    .A2(_08228_),
    .B1(net1781),
    .B2(net2028),
    .C(_08256_),
    .ZN(_08257_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1618 (.I(_03879_),
    .Z(net1617));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12432_ (.I0(_08218_),
    .I1(net1694),
    .S(_07772_),
    .Z(_08259_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12433_ (.A1(_08187_),
    .A2(_08257_),
    .B(_08259_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12434_ (.I(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .ZN(_08260_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1617 (.I(_04583_),
    .Z(net1616));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1614 (.I(_05837_),
    .Z(net1613));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12437_ (.A1(net1962),
    .A2(_08043_),
    .Z(_08263_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12438_ (.A1(_07613_),
    .A2(_07619_),
    .B(_08263_),
    .C(net1816),
    .ZN(_08264_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12439_ (.A1(_08260_),
    .A2(_08041_),
    .B(_08264_),
    .C(_08049_),
    .ZN(_08265_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12440_ (.A1(_07613_),
    .A2(_07619_),
    .B(\cs_registers_i.pc_id_i[2] ),
    .C(net1816),
    .ZN(_08266_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12441_ (.A1(_08041_),
    .A2(net1781),
    .B(_08266_),
    .C(net2063),
    .ZN(_08267_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12442_ (.A1(_08265_),
    .A2(_08267_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12443_ (.I(_01151_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12444_ (.I(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .ZN(_08268_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1613 (.I(_07695_),
    .Z(net1612));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12446_ (.A1(net1960),
    .A2(_08043_),
    .Z(_08270_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12447_ (.A1(_07613_),
    .A2(_07619_),
    .B(_08270_),
    .C(net1816),
    .ZN(_08271_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12448_ (.A1(_08268_),
    .A2(_08041_),
    .B(_08271_),
    .C(_08049_),
    .ZN(_08272_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12449_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net1994),
    .S1(net1973),
    .Z(_08273_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12450_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S0(net1994),
    .S1(net1973),
    .Z(_08274_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1612 (.I(_07772_),
    .Z(net1611));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1611 (.I(_07997_),
    .Z(net1610));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12453_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S0(net1995),
    .S1(net1973),
    .Z(_08277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12454_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net1994),
    .Z(_08278_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12455_ (.A1(net1994),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .Z(_08279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12456_ (.I0(_08278_),
    .I1(_08279_),
    .S(net1874),
    .Z(_08280_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1615 (.I(_04672_),
    .Z(net1614));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12458_ (.I0(_08273_),
    .I1(_08274_),
    .I2(_08277_),
    .I3(_08280_),
    .S0(net1877),
    .S1(net1866),
    .Z(_08282_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12459_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net1995),
    .S1(net1973),
    .Z(_08283_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12460_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S0(net1995),
    .S1(net1973),
    .Z(_08284_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1616 (.I(_04636_),
    .Z(net1615));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1665 (.I(net1663),
    .Z(net1664));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12463_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net1994),
    .S1(net1973),
    .Z(_08287_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12464_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S0(net1994),
    .S1(net1973),
    .Z(_08288_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12465_ (.I0(_08283_),
    .I1(_08284_),
    .I2(_08287_),
    .I3(_08288_),
    .S0(net1877),
    .S1(net1866),
    .Z(_08289_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12466_ (.A1(net1843),
    .A2(_08289_),
    .Z(_08290_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12467_ (.A1(net1958),
    .A2(_08282_),
    .B(_08290_),
    .ZN(_08291_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12468_ (.A1(_07613_),
    .A2(_07619_),
    .B(\cs_registers_i.pc_id_i[3] ),
    .C(net1816),
    .ZN(_08292_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12469_ (.A1(_08041_),
    .A2(net1780),
    .B(_08292_),
    .C(net2063),
    .ZN(_08293_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12470_ (.A1(_08272_),
    .A2(_08293_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12471_ (.I(net2103),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12472_ (.I(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .ZN(_08294_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12473_ (.A1(net1958),
    .A2(net1816),
    .A3(_08043_),
    .Z(_08295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12474_ (.A1(_07613_),
    .A2(_07619_),
    .B(_08295_),
    .ZN(_08296_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12475_ (.A1(_08294_),
    .A2(_08041_),
    .B(_08296_),
    .C(_08049_),
    .ZN(_08297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12476_ (.A1(net2193),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B(_08003_),
    .ZN(_08298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1666 (.I(_09772_),
    .Z(net1665));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12478_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08300_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1609 (.I(_09595_),
    .Z(net1608));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12480_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08302_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12481_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08303_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12482_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08304_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1668 (.I(net1666),
    .Z(net1667));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12484_ (.I0(_08300_),
    .I1(_08302_),
    .I2(_08303_),
    .I3(_08304_),
    .S0(net1883),
    .S1(net1959),
    .Z(_08306_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12485_ (.A1(net1842),
    .A2(_08306_),
    .ZN(_08307_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12486_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S0(net2000),
    .S1(net1973),
    .Z(_08308_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12487_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S0(net2003),
    .S1(net1973),
    .Z(_08309_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12488_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12489_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net1989),
    .Z(_08311_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12490_ (.A1(net1870),
    .A2(_08311_),
    .Z(_08312_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12491_ (.I0(_08308_),
    .I1(_08309_),
    .I2(_08310_),
    .I3(_08312_),
    .S0(net1883),
    .S1(net1867),
    .Z(_08313_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12492_ (.A1(net1958),
    .A2(_08313_),
    .ZN(_08314_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12493_ (.A1(_08298_),
    .A2(_08307_),
    .A3(_08314_),
    .Z(_08315_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12494_ (.A1(_07613_),
    .A2(_07619_),
    .B(\cs_registers_i.pc_id_i[4] ),
    .C(net1816),
    .ZN(_08316_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12495_ (.A1(_08041_),
    .A2(_08315_),
    .B(_08316_),
    .C(net2063),
    .ZN(_08317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12496_ (.A1(_08297_),
    .A2(_08317_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12497_ (.I(_01165_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1610 (.I(net1608),
    .Z(net1609));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1607 (.I(_09764_),
    .Z(net1606));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1603 (.I(_09796_),
    .Z(net1602));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12501_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net2134),
    .S1(net1973),
    .Z(_08321_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12502_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S0(net2134),
    .S1(net1973),
    .Z(_08322_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1601 (.I(_09819_),
    .Z(net1600));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12504_ (.I0(_08321_),
    .I1(_08322_),
    .S(net1881),
    .Z(_08324_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1602 (.I(_09801_),
    .Z(net1601));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12506_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net2005),
    .S1(net1962),
    .Z(_08326_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12507_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .S0(net2005),
    .S1(net1962),
    .Z(_08327_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1598 (.I(net2495),
    .Z(net1597));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12509_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S0(net2005),
    .S1(net1962),
    .Z(_08329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12510_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .S(net2005),
    .Z(_08330_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12511_ (.A1(net2005),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .Z(_08331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12512_ (.I0(_08330_),
    .I1(_08331_),
    .S(_07518_),
    .Z(_08332_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1590 (.I(_09950_),
    .Z(net1589));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12514_ (.I0(_08326_),
    .I1(_08327_),
    .I2(_08329_),
    .I3(_08332_),
    .S0(net1870),
    .S1(net1864),
    .Z(_08334_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12515_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net2134),
    .S1(net1973),
    .Z(_08335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12516_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S0(net2134),
    .S1(net1973),
    .Z(_08336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12517_ (.I0(_08335_),
    .I1(_08336_),
    .S(net1881),
    .Z(_08337_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12518_ (.A1(_07547_),
    .A2(_08337_),
    .Z(_08338_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12519_ (.A1(_07523_),
    .A2(_08324_),
    .B1(_08334_),
    .B2(net1958),
    .C(_08338_),
    .ZN(_08339_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1589 (.I(_03987_),
    .Z(net1588));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12521_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(net2063),
    .ZN(_08341_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1588 (.I(_04669_),
    .Z(net1587));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1587 (.I(_07742_),
    .Z(net1586));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12524_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(net1818),
    .ZN(_08344_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12525_ (.A1(net2126),
    .A2(net1778),
    .B1(_08341_),
    .B2(net1741),
    .C(_08344_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12526_ (.I(net1692),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1600 (.I(net1598),
    .Z(net1599));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12528_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net2137),
    .S1(net1967),
    .Z(_08346_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12529_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S0(net2003),
    .S1(net1968),
    .Z(_08347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12530_ (.I0(_08346_),
    .I1(_08347_),
    .S(net1882),
    .Z(_08348_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12531_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net2137),
    .S1(net1967),
    .Z(_08349_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1604 (.I(_09783_),
    .Z(net1603));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12533_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S0(net2137),
    .S1(net1967),
    .Z(_08351_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12534_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S0(net2005),
    .S1(net1964),
    .Z(_08352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12535_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net2005),
    .Z(_08353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12536_ (.A1(net2005),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .Z(_08354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12537_ (.I0(_08353_),
    .I1(_08354_),
    .S(net1869),
    .Z(_08355_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12538_ (.I0(_08349_),
    .I1(_08351_),
    .I2(_08352_),
    .I3(_08355_),
    .S0(net1882),
    .S1(net1864),
    .Z(_08356_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12539_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S0(net2005),
    .S1(net1964),
    .Z(_08357_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12540_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S0(net2005),
    .S1(net1964),
    .Z(_08358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12541_ (.I0(_08357_),
    .I1(_08358_),
    .S(net1882),
    .Z(_08359_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12542_ (.A1(_07547_),
    .A2(_08359_),
    .Z(_08360_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12543_ (.A1(_07523_),
    .A2(_08348_),
    .B1(_08356_),
    .B2(net1958),
    .C(_08360_),
    .ZN(_08361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12544_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(net2063),
    .ZN(_08362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12545_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net1818),
    .ZN(_08363_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12546_ (.A1(net2126),
    .A2(net1777),
    .B1(_08362_),
    .B2(net1741),
    .C(_08363_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12547_ (.I(net1691),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12548_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net2009),
    .S1(net1975),
    .Z(_08364_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12549_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S0(net2009),
    .S1(net1975),
    .Z(_08365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12550_ (.I0(_08364_),
    .I1(_08365_),
    .S(net1878),
    .Z(_08366_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12551_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net2008),
    .S1(net1975),
    .Z(_08367_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12552_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S0(net2008),
    .S1(net1975),
    .Z(_08368_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12553_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S0(net2008),
    .S1(net1975),
    .Z(_08369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12554_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net2008),
    .Z(_08370_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12555_ (.A1(net2193),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .Z(_08371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12556_ (.I0(_08370_),
    .I1(_08371_),
    .S(net1868),
    .Z(_08372_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12557_ (.I0(_08367_),
    .I1(_08368_),
    .I2(_08369_),
    .I3(_08372_),
    .S0(net1878),
    .S1(net1866),
    .Z(_08373_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12558_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S0(net2193),
    .S1(net1975),
    .Z(_08374_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12559_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S0(net2193),
    .S1(net1975),
    .Z(_08375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12560_ (.I0(_08374_),
    .I1(_08375_),
    .S(net1878),
    .Z(_08376_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12561_ (.A1(net1832),
    .A2(_08376_),
    .Z(_08377_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12562_ (.A1(net1876),
    .A2(_08366_),
    .B1(net1958),
    .B2(_08373_),
    .C(_08377_),
    .ZN(_08378_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12563_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(net2063),
    .ZN(_08379_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12564_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net1818),
    .ZN(_08380_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12565_ (.A1(net2126),
    .A2(net1776),
    .B1(_08379_),
    .B2(net2052),
    .C(_08380_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12566_ (.I(net2116),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12567_ (.I(_00841_),
    .ZN(_08381_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12568_ (.A1(_00833_),
    .A2(_00832_),
    .Z(_08382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12569_ (.A1(_08382_),
    .A2(_00837_),
    .B(_00836_),
    .ZN(_08383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12570_ (.I(_00821_),
    .ZN(_08384_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12571_ (.I(_00820_),
    .ZN(_08385_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12572_ (.A1(_08384_),
    .A2(_00010_),
    .B(_08385_),
    .ZN(_08386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12573_ (.A1(_00825_),
    .A2(_00829_),
    .Z(_08387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12574_ (.A1(_00824_),
    .A2(_00829_),
    .B(_00828_),
    .ZN(_08388_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12575_ (.A1(_00832_),
    .A2(_00836_),
    .ZN(_08389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12576_ (.A1(_08388_),
    .A2(_08389_),
    .ZN(_08390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12577_ (.A1(_08387_),
    .A2(_08386_),
    .B(_08390_),
    .ZN(_08391_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12578_ (.I(_00840_),
    .ZN(_08392_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12579_ (.A1(_08381_),
    .A2(net2178),
    .A3(net2125),
    .B(_08392_),
    .ZN(_08393_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12580_ (.A1(net2082),
    .A2(_08393_),
    .Z(net183));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12581_ (.A1(_00833_),
    .A2(_00837_),
    .A3(_08387_),
    .Z(_08394_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12582_ (.A1(_00817_),
    .A2(net2071),
    .Z(_08395_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12583_ (.A1(_00841_),
    .A2(_08394_),
    .A3(_08395_),
    .Z(_08396_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12584_ (.A1(net2290),
    .A2(_00837_),
    .ZN(_08397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12585_ (.A1(_00837_),
    .A2(_00832_),
    .B(_00836_),
    .ZN(_08398_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12586_ (.A1(_08397_),
    .A2(net2300),
    .B(_08398_),
    .ZN(_08399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12587_ (.A1(_00821_),
    .A2(_00816_),
    .Z(_08400_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12588_ (.A1(_00820_),
    .A2(_08400_),
    .Z(_08401_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12589_ (.A1(_00841_),
    .A2(net2291),
    .A3(_08401_),
    .Z(_08402_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12590_ (.A1(_08172_),
    .A2(_08178_),
    .A3(_08183_),
    .Z(_08403_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12591_ (.A1(_08215_),
    .A2(net2121),
    .B(_08402_),
    .C(_08403_),
    .ZN(_08404_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12592_ (.A1(_00841_),
    .A2(net2291),
    .A3(_08394_),
    .Z(_08405_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12593_ (.A1(_00841_),
    .A2(net2291),
    .A3(_08401_),
    .A4(_08395_),
    .Z(_08406_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12594_ (.A1(_08394_),
    .A2(_08401_),
    .Z(_08407_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12595_ (.A1(net2291),
    .A2(_08407_),
    .B(_00841_),
    .ZN(_08408_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _12596_ (.A1(_08405_),
    .A2(_08406_),
    .A3(_08408_),
    .ZN(_08409_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12597_ (.A1(net2111),
    .A2(_08396_),
    .B(_08404_),
    .C(_08409_),
    .ZN(net182));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1605 (.I(net1603),
    .Z(net1604));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1606 (.I(net1603),
    .Z(net1605));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1608 (.I(_09764_),
    .Z(net1607));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12601_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net2010),
    .S1(net1977),
    .Z(_08413_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12602_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S0(net2010),
    .S1(net1977),
    .Z(_08414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12603_ (.I0(_08413_),
    .I1(_08414_),
    .S(net1878),
    .Z(_08415_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12604_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S0(net2013),
    .S1(net1984),
    .Z(_08416_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12605_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S0(net2013),
    .S1(net1984),
    .Z(_08417_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12606_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net2193),
    .S1(net1975),
    .Z(_08418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12607_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net2008),
    .Z(_08419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12608_ (.A1(net2193),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .Z(_08420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12609_ (.I0(_08419_),
    .I1(_08420_),
    .S(net1868),
    .Z(_08421_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12610_ (.I0(_08416_),
    .I1(_08417_),
    .I2(_08418_),
    .I3(_08421_),
    .S0(net1878),
    .S1(net1866),
    .Z(_08422_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12611_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S0(net2010),
    .S1(net1977),
    .Z(_08423_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12612_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S0(net2010),
    .S1(net1977),
    .Z(_08424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12613_ (.I0(_08423_),
    .I1(_08424_),
    .S(net1878),
    .Z(_08425_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12614_ (.A1(net1832),
    .A2(_08425_),
    .Z(_08426_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12615_ (.A1(net1876),
    .A2(_08415_),
    .B1(_08422_),
    .B2(net1958),
    .C(_08426_),
    .ZN(_08427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12616_ (.A1(\cs_registers_i.pc_id_i[8] ),
    .A2(net2063),
    .ZN(_08428_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1670 (.I(net1668),
    .Z(net1669));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12618_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(net2483),
    .ZN(_08430_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12619_ (.A1(net1775),
    .A2(net2127),
    .B1(_08428_),
    .B2(net2053),
    .C(_08430_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12620_ (.I(net2072),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1586 (.I(_09779_),
    .Z(net1585));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload12 (.I(clknet_leaf_7_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload13 (.I(clknet_leaf_16_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12624_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08434_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1584 (.I(_09839_),
    .Z(net1583));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12626_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08436_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12627_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08437_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12628_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08438_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12629_ (.I0(_08434_),
    .I1(_08436_),
    .I2(_08437_),
    .I3(_08438_),
    .S0(net1884),
    .S1(net1867),
    .Z(_08439_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12630_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S0(net2000),
    .S1(net1962),
    .Z(_08440_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12631_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .S0(net2000),
    .S1(net1962),
    .Z(_08441_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12632_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net2000),
    .S1(net1962),
    .Z(_08442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12633_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .S(net2000),
    .Z(_08443_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12634_ (.A1(net2000),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .Z(_08444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12635_ (.I0(_08443_),
    .I1(_08444_),
    .S(net1881),
    .Z(_08445_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12636_ (.I0(_08440_),
    .I1(_08441_),
    .I2(_08442_),
    .I3(_08445_),
    .S0(net1873),
    .S1(net1867),
    .Z(_08446_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12637_ (.A1(net1958),
    .A2(_08446_),
    .Z(_08447_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12638_ (.A1(net1842),
    .A2(_08439_),
    .B(_08447_),
    .ZN(_08448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12639_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(net2063),
    .ZN(_08449_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12640_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(net2483),
    .ZN(_08450_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12641_ (.A1(net2127),
    .A2(net1736),
    .B1(_08449_),
    .B2(net2053),
    .C(_08450_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12642_ (.I(net2097),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12643_ (.A1(_00841_),
    .A2(net2082),
    .ZN(_08451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12644_ (.A1(_00845_),
    .A2(_00840_),
    .B(_00844_),
    .ZN(_08452_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12645_ (.A1(net2178),
    .A2(net2125),
    .A3(_08451_),
    .B(_08452_),
    .ZN(_08453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12646_ (.A1(net2073),
    .A2(_08453_),
    .B(_00848_),
    .ZN(_08454_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _12647_ (.A1(_00853_),
    .A2(_08454_),
    .Z(_08455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12648_ (.I(_08455_),
    .ZN(net185));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12649_ (.I(net2109),
    .ZN(_08456_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12650_ (.A1(_00820_),
    .A2(_08400_),
    .ZN(_08457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12651_ (.I(_00824_),
    .ZN(_08458_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12652_ (.A1(_08456_),
    .A2(_08457_),
    .B(_08458_),
    .ZN(_08459_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12653_ (.A1(_00829_),
    .A2(_08459_),
    .B(_00828_),
    .ZN(_08460_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12654_ (.A1(_08397_),
    .A2(_08451_),
    .ZN(_08461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12655_ (.I(_08461_),
    .ZN(_08462_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12656_ (.A1(_08381_),
    .A2(_08398_),
    .B(_08392_),
    .ZN(_08463_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12657_ (.A1(net2082),
    .A2(_08463_),
    .B(_00844_),
    .ZN(_08464_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12658_ (.A1(_08460_),
    .A2(_08462_),
    .B(_08464_),
    .ZN(_08465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12659_ (.A1(_08387_),
    .A2(_08395_),
    .Z(_08466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12660_ (.I(_08466_),
    .ZN(_08467_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12661_ (.A1(_08466_),
    .A2(_08461_),
    .Z(_08468_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12662_ (.A1(_08112_),
    .A2(_08120_),
    .B(_08128_),
    .C(_08468_),
    .ZN(_08469_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_4 _12663_ (.A1(_08184_),
    .A2(_08467_),
    .A3(_08462_),
    .B1(_08170_),
    .B2(_08469_),
    .ZN(_08470_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12664_ (.A1(_08465_),
    .A2(_08470_),
    .B(net2073),
    .ZN(_08471_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12665_ (.A1(net2073),
    .A2(_08465_),
    .A3(_08470_),
    .Z(_08472_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12666_ (.A1(_08471_),
    .A2(_08472_),
    .Z(net184));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12667_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net1990),
    .S1(net1974),
    .Z(_08473_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12668_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S0(net1990),
    .S1(net1974),
    .Z(_08474_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12669_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S0(net2000),
    .S1(net1974),
    .Z(_08475_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12670_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S0(net2000),
    .S1(net1974),
    .Z(_08476_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12671_ (.I0(_08473_),
    .I1(_08474_),
    .I2(_08475_),
    .I3(_08476_),
    .S0(net1881),
    .S1(net1867),
    .Z(_08477_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12672_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S0(net1989),
    .S1(net1974),
    .Z(_08478_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12673_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S0(net1989),
    .S1(net1974),
    .Z(_08479_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12674_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net1989),
    .S1(net1974),
    .Z(_08480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12675_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net1994),
    .Z(_08481_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12676_ (.A1(net2134),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .Z(_08482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12677_ (.I0(_08481_),
    .I1(_08482_),
    .S(net1874),
    .Z(_08483_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12678_ (.I0(_08478_),
    .I1(_08479_),
    .I2(_08480_),
    .I3(_08483_),
    .S0(net1881),
    .S1(net1867),
    .Z(_08484_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _12679_ (.A1(net1958),
    .A2(_08484_),
    .Z(_08485_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12680_ (.A1(net1842),
    .A2(_08477_),
    .B(_08485_),
    .ZN(_08486_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12681_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(net2064),
    .ZN(_08487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12682_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net2483),
    .ZN(_08488_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12683_ (.A1(net2127),
    .A2(net1735),
    .B1(_08487_),
    .B2(net2053),
    .C(_08488_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12684_ (.I(net2102),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12685_ (.I(_00856_),
    .ZN(_08489_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12686_ (.A1(_00849_),
    .A2(_00853_),
    .ZN(_08490_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _12687_ (.A1(_08391_),
    .A2(_08383_),
    .A3(_08451_),
    .A4(_08490_),
    .ZN(_08491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12688_ (.A1(_00853_),
    .A2(_00848_),
    .B(_00852_),
    .ZN(_08492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12689_ (.A1(_08452_),
    .A2(_08490_),
    .B(_08492_),
    .ZN(_08493_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12690_ (.A1(_08491_),
    .A2(_08493_),
    .B(net2173),
    .ZN(_08494_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12691_ (.I(net2062),
    .ZN(_08495_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12692_ (.A1(_08489_),
    .A2(_08494_),
    .B(_08495_),
    .ZN(_08496_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12693_ (.A1(_08495_),
    .A2(_08489_),
    .A3(_08494_),
    .Z(_08497_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12694_ (.A1(_08496_),
    .A2(_08497_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12695_ (.A1(_00841_),
    .A2(net2082),
    .Z(_08498_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12696_ (.A1(_08401_),
    .A2(_08395_),
    .B(_08394_),
    .ZN(_08499_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12697_ (.A1(net2300),
    .A2(_08397_),
    .B(_08499_),
    .C(_08398_),
    .ZN(_08500_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12698_ (.A1(_08498_),
    .A2(_08500_),
    .ZN(_08501_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _12699_ (.A1(_08401_),
    .A2(_08399_),
    .ZN(_08502_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12700_ (.I(_08502_),
    .ZN(_08503_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _12701_ (.A1(_08215_),
    .A2(net2121),
    .B(_08403_),
    .C(_08503_),
    .ZN(_08504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12702_ (.A1(_08452_),
    .A2(_08490_),
    .ZN(_08505_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12703_ (.A1(_00853_),
    .A2(_00848_),
    .Z(_08506_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _12704_ (.A1(_00852_),
    .A2(_08505_),
    .A3(_08506_),
    .ZN(_08507_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12705_ (.A1(_08490_),
    .A2(_08501_),
    .A3(net2094),
    .B(_08507_),
    .ZN(_08508_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _12706_ (.A1(net2173),
    .A2(_08508_),
    .ZN(_08509_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _12707_ (.I(_08509_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1585 (.I(net1583),
    .Z(net1584));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1583 (.I(_09894_),
    .Z(net1582));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1582 (.I(_10012_),
    .Z(net1581));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1581 (.I(_03989_),
    .Z(net1580));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1580 (.I(_04152_),
    .Z(net1579));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1579 (.I(_04676_),
    .Z(net1578));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload14 (.I(clknet_leaf_17_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12716_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08518_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload15 (.I(clknet_leaf_18_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload16 (.I(clknet_leaf_20_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12719_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08521_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload17 (.I(clknet_leaf_21_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload18 (.I(clknet_leaf_22_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload19 (.I(clknet_leaf_23_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12723_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08525_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12724_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08526_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload20 (.I(clknet_leaf_24_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload21 (.I(clknet_leaf_26_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1576 (.I(_00293_),
    .Z(net1575));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1577 (.I(net1575),
    .Z(net1576));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12729_ (.I0(_08518_),
    .I1(_08521_),
    .I2(_08525_),
    .I3(_08526_),
    .S0(net1849),
    .S1(net1901),
    .Z(_08531_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1578 (.I(net1576),
    .Z(net1577));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1569 (.I(_00486_),
    .Z(net1568));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12732_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12733_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net2089),
    .Z(_08535_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1568 (.I(_00589_),
    .Z(net1567));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1567 (.I(_00680_),
    .Z(net1566));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12736_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A2(_07745_),
    .B1(_08535_),
    .B2(net1946),
    .ZN(_08538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12737_ (.I(_08538_),
    .ZN(_08539_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12738_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08540_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12739_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S0(net1946),
    .S1(net1910),
    .Z(_08541_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12740_ (.I0(_08534_),
    .I1(_08539_),
    .I2(_08540_),
    .I3(_08541_),
    .S0(net1849),
    .S1(net1901),
    .Z(_08542_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1570 (.I(_00412_),
    .Z(net1569));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12742_ (.I0(_08531_),
    .I1(_08542_),
    .S(net1862),
    .Z(_08544_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1571 (.I(_00336_),
    .Z(net1570));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12744_ (.I(net1891),
    .ZN(_08546_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12745_ (.A1(net1800),
    .A2(_07767_),
    .Z(_08547_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _12746_ (.A1(_08547_),
    .A2(_07699_),
    .A3(_08546_),
    .Z(_08548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12747_ (.A1(_07767_),
    .A2(net1800),
    .ZN(_08549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12748_ (.A1(net1800),
    .A2(net1799),
    .A3(_07767_),
    .Z(_08550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12749_ (.A1(_08549_),
    .A2(_08550_),
    .ZN(_08551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12750_ (.A1(net2022),
    .A2(_08551_),
    .ZN(_08552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12751_ (.A1(net2060),
    .A2(_08552_),
    .ZN(_08553_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1565 (.I(_10149_),
    .Z(net1564));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1566 (.I(_10149_),
    .Z(net1565));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12754_ (.I0(net1687),
    .I1(_08553_),
    .S(net1795),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1572 (.I(net1570),
    .Z(net1571));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1564 (.I(_10183_),
    .Z(net1563));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1563 (.I(_10247_),
    .Z(net1562));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1573 (.I(net1570),
    .Z(net1572));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12759_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .B2(_08197_),
    .C1(_08200_),
    .C2(net1687),
    .ZN(_08560_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12760_ (.A1(net2028),
    .A2(net1803),
    .B(_08560_),
    .ZN(_08561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12761_ (.I0(net1693),
    .I1(net2111),
    .S(_01225_),
    .Z(_08562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12762_ (.A1(_08187_),
    .A2(_08561_),
    .B(_08562_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1574 (.I(net1572),
    .Z(net1573));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1575 (.I(net1573),
    .Z(net1574));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload22 (.I(clknet_leaf_5_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08566_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload23 (.I(clknet_leaf_6_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12768_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08568_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload24 (.I(clknet_leaf_8_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12770_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08570_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload25 (.I(clknet_leaf_9_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload26 (.I(clknet_leaf_11_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12774_ (.I0(_08566_),
    .I1(_08568_),
    .I2(_08570_),
    .I3(_08571_),
    .S0(net1852),
    .S1(net1902),
    .Z(_08574_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12775_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12776_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net1918),
    .Z(_08576_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1562 (.I(_10159_),
    .Z(net1561));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12778_ (.A1(net1918),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .Z(_08578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1561 (.I(_10162_),
    .Z(net1560));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12781_ (.I0(_08576_),
    .I1(_08578_),
    .S(net1853),
    .Z(_08581_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12782_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S0(net1954),
    .S1(net1920),
    .Z(_08582_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12783_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S0(net1954),
    .S1(net1918),
    .Z(_08583_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12784_ (.I0(_08575_),
    .I1(_08581_),
    .I2(_08582_),
    .I3(_08583_),
    .S0(net1852),
    .S1(net1902),
    .Z(_08584_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1560 (.I(_10188_),
    .Z(net1559));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12786_ (.I0(_08574_),
    .I1(_08584_),
    .S(net1863),
    .Z(_08586_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12787_ (.A1(net2020),
    .A2(_08551_),
    .ZN(_08587_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12788_ (.A1(_08548_),
    .A2(_08587_),
    .ZN(_08588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12789_ (.I0(net1774),
    .I1(_08588_),
    .S(net1795),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12790_ (.A1(net1958),
    .A2(net1959),
    .Z(_08589_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12791_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net1997),
    .S1(net1962),
    .Z(_08590_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12792_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .S0(net1997),
    .S1(net1962),
    .Z(_08591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12793_ (.I0(_08590_),
    .I1(_08591_),
    .S(net1874),
    .Z(_08592_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12794_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08593_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12795_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12796_ (.I0(_08593_),
    .I1(_08594_),
    .S(net1879),
    .Z(_08595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12797_ (.A1(net1958),
    .A2(net1866),
    .Z(_08596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12798_ (.A1(_08589_),
    .A2(_08592_),
    .B1(_08595_),
    .B2(net1822),
    .ZN(_08597_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12799_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12800_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net1997),
    .Z(_08599_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12801_ (.A1(net1997),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .Z(_08600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12802_ (.I0(_08599_),
    .I1(_08600_),
    .S(net1874),
    .Z(_08601_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12803_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08602_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12804_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08603_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12805_ (.I0(_08598_),
    .I1(_08601_),
    .I2(_08602_),
    .I3(_08603_),
    .S0(net1880),
    .S1(net1959),
    .Z(_08604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _12806_ (.A1(net1842),
    .A2(_08604_),
    .ZN(_08605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12807_ (.A1(net1813),
    .A2(_08605_),
    .Z(_08606_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12808_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1774),
    .ZN(_08607_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12809_ (.A1(net2028),
    .A2(net1734),
    .B(_08607_),
    .ZN(_08608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12810_ (.I0(net1693),
    .I1(net1694),
    .S(_01229_),
    .Z(_08609_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12811_ (.A1(_08187_),
    .A2(_08608_),
    .B(_08609_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12812_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(net1801),
    .ZN(_08610_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1559 (.I(_10197_),
    .Z(net1558));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12814_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net1818),
    .ZN(_08612_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _12815_ (.A1(net2127),
    .A2(net1734),
    .B1(_08610_),
    .B2(net1741),
    .C(_08612_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12816_ (.I(net2070),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _12817_ (.A1(net2178),
    .A2(net2124),
    .A3(_08451_),
    .A4(_08490_),
    .Z(_08613_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12818_ (.I(net2173),
    .ZN(_08614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12819_ (.A1(_08613_),
    .A2(_08507_),
    .B(_08614_),
    .ZN(_08615_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12820_ (.A1(_00856_),
    .A2(_08615_),
    .B(net2088),
    .C(net2062),
    .ZN(_08616_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _12821_ (.A1(_00865_),
    .A2(_00860_),
    .B(_00864_),
    .ZN(_08617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12822_ (.A1(_08616_),
    .A2(_08617_),
    .Z(_08618_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12823_ (.A1(net2083),
    .A2(_08618_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12824_ (.A1(_00857_),
    .A2(_00861_),
    .Z(_08619_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _12825_ (.A1(net2073),
    .A2(_00853_),
    .A3(_08619_),
    .Z(_08620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12826_ (.A1(net2484),
    .A2(_08620_),
    .Z(_08621_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12827_ (.A1(net2088),
    .A2(_08620_),
    .ZN(_08622_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12828_ (.A1(_08614_),
    .A2(_08492_),
    .B(_08489_),
    .ZN(_08623_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12829_ (.A1(net2062),
    .A2(_08623_),
    .B(_00860_),
    .ZN(_08624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12830_ (.I0(net2088),
    .I1(_08622_),
    .S(_08624_),
    .Z(_08625_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12831_ (.I(net2088),
    .ZN(_08626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12832_ (.A1(_08626_),
    .A2(_08624_),
    .ZN(_08627_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12833_ (.A1(_08465_),
    .A2(_08627_),
    .ZN(_08628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12834_ (.I0(_08628_),
    .I1(_08621_),
    .S(_08470_),
    .Z(_08629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _12835_ (.A1(_08465_),
    .A2(_08621_),
    .B(_08625_),
    .C(_08629_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1558 (.I(_10197_),
    .Z(net1557));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1557 (.I(_10203_),
    .Z(net1556));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12838_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S0(net1950),
    .S1(net1911),
    .Z(_08632_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12839_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S0(net1950),
    .S1(net1911),
    .Z(_08633_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload27 (.I(clknet_leaf_12_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1556 (.I(_10211_),
    .Z(net1555));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12842_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net2114),
    .S1(net1911),
    .Z(_08636_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net1950),
    .S1(net1911),
    .Z(_08637_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload28 (.I(clknet_leaf_13_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1555 (.I(_10216_),
    .Z(net1554));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12846_ (.I0(_08632_),
    .I1(_08633_),
    .I2(_08636_),
    .I3(_08637_),
    .S0(net1850),
    .S1(net1901),
    .Z(_08640_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12847_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net1949),
    .S1(net1919),
    .Z(_08641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12848_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net2089),
    .Z(_08642_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12849_ (.A1(net2089),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .Z(_08643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12850_ (.I0(_08642_),
    .I1(_08643_),
    .S(net1853),
    .Z(_08644_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1554 (.I(_10219_),
    .Z(net1553));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12852_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08646_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12853_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08647_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12854_ (.I0(_08641_),
    .I1(_08644_),
    .I2(_08646_),
    .I3(_08647_),
    .S0(net1850),
    .S1(net1901),
    .Z(_08648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12855_ (.I0(_08640_),
    .I1(_08648_),
    .S(net1863),
    .Z(_08649_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12856_ (.A1(net2019),
    .A2(_08551_),
    .ZN(_08650_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12857_ (.A1(net2060),
    .A2(_08650_),
    .ZN(_08651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12858_ (.I0(net1773),
    .I1(_08651_),
    .S(net1795),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12859_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net1993),
    .S1(net1969),
    .Z(_08652_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12860_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net1993),
    .S1(net1969),
    .Z(_08653_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12861_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S0(net1993),
    .S1(net1969),
    .Z(_08654_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12862_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S0(net1993),
    .S1(net1969),
    .Z(_08655_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_4 _12863_ (.I0(_08652_),
    .I1(_08653_),
    .I2(_08654_),
    .I3(_08655_),
    .S0(net1881),
    .S1(net1866),
    .Z(_08656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12864_ (.A1(net1871),
    .A2(net1989),
    .Z(_08657_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1553 (.I(_10239_),
    .Z(net1552));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12866_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net1991),
    .Z(_08659_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _12867_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .A2(net1820),
    .B1(_08659_),
    .B2(net1970),
    .C(net1962),
    .ZN(_08660_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload30 (.I(clknet_leaf_15_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12869_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_08662_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12870_ (.A1(net1881),
    .A2(_08662_),
    .B(net1866),
    .ZN(_08663_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12871_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_08664_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_08665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12873_ (.I0(_08664_),
    .I1(_08665_),
    .S(net1881),
    .Z(_08666_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12874_ (.A1(net1961),
    .A2(_08666_),
    .ZN(_08667_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12875_ (.A1(_08660_),
    .A2(_08663_),
    .B(_08667_),
    .C(net1842),
    .ZN(_08668_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _12876_ (.A1(net1842),
    .A2(_08656_),
    .B(_08668_),
    .ZN(_08669_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12877_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .B2(_08197_),
    .C1(_08200_),
    .C2(net1773),
    .ZN(_08670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12878_ (.A1(net2028),
    .A2(net1733),
    .B(_08670_),
    .ZN(_08671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12879_ (.I0(net1693),
    .I1(net2111),
    .S(_01236_),
    .Z(_08672_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12880_ (.A1(_08187_),
    .A2(_08671_),
    .B(_08672_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12881_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(net1801),
    .ZN(_08673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12882_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net1818),
    .ZN(_08674_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12883_ (.A1(net1742),
    .A2(net1733),
    .B1(_08673_),
    .B2(net1741),
    .C(_08674_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12884_ (.I(net1685),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload29 (.I(clknet_leaf_14_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1552 (.I(_04596_),
    .Z(net1551));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net2188),
    .S1(net1921),
    .Z(_08677_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S0(net2188),
    .S1(net1921),
    .Z(_08678_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12889_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net2188),
    .S1(net1921),
    .Z(_08679_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net2188),
    .S1(net1921),
    .Z(_08681_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12892_ (.I0(_08677_),
    .I1(_08678_),
    .I2(_08679_),
    .I3(_08681_),
    .S0(net1852),
    .S1(net1902),
    .Z(_08682_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net2188),
    .S1(net1919),
    .Z(_08683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12894_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net1919),
    .Z(_08684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12895_ (.A1(net1919),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .Z(_08685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12896_ (.I0(_08684_),
    .I1(_08685_),
    .S(net1853),
    .Z(_08686_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12897_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net2188),
    .S1(net1918),
    .Z(_08687_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12898_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S0(net2188),
    .S1(net1918),
    .Z(_08688_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12899_ (.I0(_08683_),
    .I1(_08686_),
    .I2(_08687_),
    .I3(_08688_),
    .S0(net1852),
    .S1(net1902),
    .Z(_08689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12900_ (.I0(_08682_),
    .I1(_08689_),
    .S(net1863),
    .Z(_08690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12901_ (.A1(net2009),
    .A2(_08551_),
    .ZN(_08691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12902_ (.A1(net2060),
    .A2(_08691_),
    .ZN(_08692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12903_ (.I0(net1772),
    .I1(_08692_),
    .S(net1795),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12904_ (.A1(net1842),
    .A2(net1866),
    .Z(_08693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12905_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net1991),
    .Z(_08694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12906_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S(net1991),
    .Z(_08695_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12907_ (.A1(net1991),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .Z(_08696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12908_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .S(net1991),
    .Z(_08697_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12910_ (.I0(_08694_),
    .I1(_08695_),
    .I2(_08696_),
    .I3(_08697_),
    .S0(net1962),
    .S1(net1874),
    .Z(_08699_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12911_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S0(net2162),
    .S1(net1968),
    .Z(_08700_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12912_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S0(net2162),
    .S1(net1968),
    .Z(_08701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12913_ (.I0(_08700_),
    .I1(_08701_),
    .S(net1880),
    .Z(_08702_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12914_ (.A1(net1842),
    .A2(net1959),
    .Z(_08703_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12915_ (.A1(_08693_),
    .A2(_08699_),
    .B1(_08702_),
    .B2(_08703_),
    .ZN(_08704_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12916_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08705_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12917_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12918_ (.I0(_08705_),
    .I1(_08706_),
    .S(net1880),
    .Z(_08707_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08708_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12920_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S0(net1997),
    .S1(net1971),
    .Z(_08709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12921_ (.I0(_08708_),
    .I1(_08709_),
    .S(net1880),
    .Z(_08710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12922_ (.A1(_08589_),
    .A2(_08707_),
    .B1(_08710_),
    .B2(net1822),
    .ZN(_08711_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12923_ (.A1(net1812),
    .A2(net1811),
    .Z(_08712_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12924_ (.A1(net2028),
    .A2(_08712_),
    .Z(_08713_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12925_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .B2(_08197_),
    .C1(_08200_),
    .C2(net1772),
    .ZN(_08714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1551 (.I(net2492),
    .Z(net1550));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12927_ (.A1(_08713_),
    .A2(_08714_),
    .B(net1814),
    .ZN(_08716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12928_ (.I0(net1693),
    .I1(net2111),
    .S(_01243_),
    .Z(_08717_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12929_ (.A1(_08716_),
    .A2(_08717_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12930_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(net1801),
    .ZN(_08718_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12931_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net1818),
    .ZN(_08719_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12932_ (.A1(net2126),
    .A2(_08712_),
    .B1(_08718_),
    .B2(net1741),
    .C(_08719_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12933_ (.I(net1684),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12934_ (.I(_08617_),
    .ZN(_08720_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12935_ (.A1(net2083),
    .A2(_08720_),
    .Z(_08721_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _12936_ (.A1(net2095),
    .A2(_08721_),
    .ZN(_08722_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12937_ (.A1(_00869_),
    .A2(_00868_),
    .Z(_08723_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _12938_ (.A1(_00865_),
    .A2(net2062),
    .A3(_08723_),
    .ZN(_08724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12939_ (.A1(_08489_),
    .A2(_08722_),
    .Z(_08725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12940_ (.A1(_08722_),
    .A2(_08724_),
    .B1(_08725_),
    .B2(_08494_),
    .ZN(_08726_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12941_ (.I(_00872_),
    .ZN(_08727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12942_ (.A1(net2077),
    .A2(_08727_),
    .ZN(_08728_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12943_ (.I(net2079),
    .ZN(_08729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12944_ (.A1(_08729_),
    .A2(net2077),
    .ZN(_08730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12945_ (.I0(net2077),
    .I1(_08730_),
    .S(_08727_),
    .Z(_08731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12946_ (.A1(_08489_),
    .A2(_08722_),
    .ZN(_08732_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _12947_ (.I(net2076),
    .ZN(_08733_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12948_ (.A1(net2079),
    .A2(_08733_),
    .Z(_08734_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12949_ (.A1(_08722_),
    .A2(_08724_),
    .ZN(_08735_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12950_ (.A1(_08615_),
    .A2(_08732_),
    .B(_08734_),
    .C(_08735_),
    .ZN(_08736_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _12951_ (.A1(_08726_),
    .A2(_08728_),
    .B(_08731_),
    .C(_08736_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12952_ (.A1(net2083),
    .A2(_08621_),
    .ZN(_08737_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _12953_ (.A1(_00860_),
    .A2(_00864_),
    .A3(_00868_),
    .Z(_08738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _12954_ (.A1(net2062),
    .A2(_00856_),
    .B1(_08493_),
    .B2(_08619_),
    .C(_08738_),
    .ZN(_08739_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12955_ (.A1(_00865_),
    .A2(_00864_),
    .A3(_00868_),
    .B(_08723_),
    .ZN(_08740_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _12956_ (.A1(_08740_),
    .A2(_08739_),
    .Z(_08741_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _12957_ (.A1(_08501_),
    .A2(net2094),
    .A3(_08737_),
    .B(net2074),
    .ZN(_08742_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _12958_ (.A1(_08729_),
    .A2(_08742_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12959_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S0(net1956),
    .S1(net1930),
    .Z(_08743_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12960_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S0(net1956),
    .S1(net1930),
    .Z(_08744_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net1956),
    .S1(net1930),
    .Z(_08745_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12962_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net1956),
    .S1(net1930),
    .Z(_08746_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12963_ (.I0(_08743_),
    .I1(_08744_),
    .I2(_08745_),
    .I3(_08746_),
    .S0(net1847),
    .S1(net1902),
    .Z(_08747_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12964_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S0(net1954),
    .S1(net1918),
    .Z(_08748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12965_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net1918),
    .Z(_08749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12966_ (.A1(net1918),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .Z(_08750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12967_ (.I0(_08749_),
    .I1(_08750_),
    .S(net1853),
    .Z(_08751_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12968_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net1954),
    .S1(net1918),
    .Z(_08752_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12969_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net2188),
    .S1(net1918),
    .Z(_08753_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12970_ (.I0(_08748_),
    .I1(_08751_),
    .I2(_08752_),
    .I3(_08753_),
    .S0(net1852),
    .S1(net1902),
    .Z(_08754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _12971_ (.I0(_08747_),
    .I1(_08754_),
    .S(net1863),
    .Z(_08755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12972_ (.A1(net1965),
    .A2(_08551_),
    .ZN(_08756_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12973_ (.A1(net2059),
    .A2(_08756_),
    .ZN(_08757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12974_ (.I0(net1771),
    .I1(_08757_),
    .S(net1795),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12975_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .S(net2164),
    .Z(_08758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12976_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(net2163),
    .Z(_08759_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _12977_ (.A1(net2163),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .Z(_08760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12978_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net2163),
    .Z(_08761_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12980_ (.I0(_08758_),
    .I1(_08759_),
    .I2(_08760_),
    .I3(_08761_),
    .S0(net1968),
    .S1(net1880),
    .Z(_08763_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S0(net2162),
    .S1(net1962),
    .Z(_08764_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12982_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .S0(net2162),
    .S1(net1962),
    .Z(_08765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12983_ (.I0(_08764_),
    .I1(_08765_),
    .S(net1874),
    .Z(_08766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12984_ (.A1(_08693_),
    .A2(_08763_),
    .B1(_08766_),
    .B2(_08703_),
    .ZN(_08767_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12985_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S0(net2164),
    .S1(net1985),
    .Z(_08768_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12986_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S0(net2164),
    .S1(net1985),
    .Z(_08769_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12987_ (.I0(_08768_),
    .I1(_08769_),
    .S(net1879),
    .Z(_08770_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12988_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S0(net2164),
    .S1(net1968),
    .Z(_08771_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _12989_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S0(net2164),
    .S1(net1968),
    .Z(_08772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12990_ (.I0(_08771_),
    .I1(_08772_),
    .S(net1879),
    .Z(_08773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _12991_ (.A1(_08589_),
    .A2(_08770_),
    .B1(_08773_),
    .B2(_08596_),
    .ZN(_08774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _12992_ (.A1(_08767_),
    .A2(_08774_),
    .Z(_08775_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _12993_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1771),
    .ZN(_08776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _12994_ (.A1(net2028),
    .A2(net1770),
    .B(_08776_),
    .ZN(_08777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _12995_ (.I0(net1693),
    .I1(net2111),
    .S(_01250_),
    .Z(_08778_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _12996_ (.A1(_08187_),
    .A2(_08777_),
    .B(_08778_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12997_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(net1801),
    .ZN(_08779_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _12998_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net2483),
    .ZN(_08780_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _12999_ (.A1(net2127),
    .A2(net1770),
    .B1(_08779_),
    .B2(net2053),
    .C(_08780_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13000_ (.I(net1683),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13001_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08781_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13002_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08782_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13003_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08783_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13004_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08784_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13005_ (.I0(_08781_),
    .I1(_08782_),
    .I2(_08783_),
    .I3(_08784_),
    .S0(net1847),
    .S1(net1901),
    .Z(_08785_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13006_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13007_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net1911),
    .Z(_08787_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13008_ (.A1(net1911),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .Z(_08788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13009_ (.I0(_08787_),
    .I1(_08788_),
    .S(net1853),
    .Z(_08789_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13010_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08790_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13011_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net1947),
    .S1(net1911),
    .Z(_08791_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13012_ (.I0(_08786_),
    .I1(_08789_),
    .I2(_08790_),
    .I3(_08791_),
    .S0(net1849),
    .S1(net1901),
    .Z(_08792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13013_ (.I0(_08785_),
    .I1(_08792_),
    .S(net1862),
    .Z(_08793_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13014_ (.A1(net1962),
    .A2(_08551_),
    .ZN(_08794_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13015_ (.A1(net2060),
    .A2(_08794_),
    .ZN(_08795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13016_ (.I0(net1769),
    .I1(_08795_),
    .S(net1795),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13017_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08796_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13018_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08797_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13019_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08798_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13020_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08799_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13021_ (.I0(_08796_),
    .I1(_08797_),
    .I2(_08798_),
    .I3(_08799_),
    .S0(net1884),
    .S1(net1867),
    .Z(_08800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13022_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net1990),
    .Z(_08801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13023_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A2(_08657_),
    .B1(_08801_),
    .B2(net1970),
    .C(net1962),
    .ZN(_08802_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13024_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08803_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13025_ (.A1(net1884),
    .A2(_08803_),
    .B(net1867),
    .ZN(_08804_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13026_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08805_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13027_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net2001),
    .S1(net1968),
    .Z(_08806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13028_ (.I0(_08805_),
    .I1(_08806_),
    .S(net1884),
    .Z(_08807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13029_ (.A1(net1961),
    .A2(_08807_),
    .ZN(_08808_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13030_ (.A1(_08802_),
    .A2(_08804_),
    .B(_08808_),
    .C(net1842),
    .ZN(_08809_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13031_ (.A1(net1842),
    .A2(_08800_),
    .B(_08809_),
    .ZN(_08810_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13032_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1769),
    .ZN(_08811_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13033_ (.A1(net2028),
    .A2(net1732),
    .B(_08811_),
    .ZN(_08812_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13035_ (.I0(net2175),
    .I1(net1694),
    .S(_01257_),
    .Z(_08814_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13036_ (.A1(_08187_),
    .A2(_08812_),
    .B(_08814_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13037_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(net1801),
    .ZN(_08815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13038_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net1818),
    .ZN(_08816_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _13039_ (.A1(net1742),
    .A2(net1732),
    .B1(_08815_),
    .B2(net1741),
    .C(_08816_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13040_ (.I(_01256_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13041_ (.A1(_00881_),
    .A2(_00877_),
    .A3(_00873_),
    .Z(_08817_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13042_ (.A1(net2484),
    .A2(_08619_),
    .A3(_08723_),
    .A4(_08817_),
    .Z(_08818_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13043_ (.A1(_08506_),
    .A2(_08505_),
    .A3(_08491_),
    .B(_08818_),
    .ZN(_08819_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13044_ (.I(_00880_),
    .ZN(_08820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13045_ (.A1(net2079),
    .A2(net2095),
    .B(_00872_),
    .ZN(_08821_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13046_ (.I(_00876_),
    .ZN(_08822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13047_ (.A1(_08733_),
    .A2(_08821_),
    .B(_08822_),
    .ZN(_08823_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13048_ (.A1(_00881_),
    .A2(_08823_),
    .ZN(_08824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13049_ (.A1(net2173),
    .A2(_00852_),
    .ZN(_08825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13050_ (.A1(_08489_),
    .A2(_08825_),
    .B(_08724_),
    .ZN(_08826_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13051_ (.A1(_08721_),
    .A2(_08826_),
    .B(_08817_),
    .ZN(_08827_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13052_ (.A1(_08827_),
    .A2(_08824_),
    .A3(_08820_),
    .Z(_08828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13053_ (.A1(net2287),
    .A2(_08828_),
    .Z(_08829_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13054_ (.A1(_00885_),
    .A2(_08829_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13055_ (.I(_00864_),
    .ZN(_08830_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13056_ (.A1(_08626_),
    .A2(_08624_),
    .B(_08830_),
    .ZN(_08831_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13057_ (.A1(net2083),
    .A2(net2079),
    .A3(net2077),
    .A4(_08831_),
    .Z(_08832_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13058_ (.A1(_08823_),
    .A2(_08832_),
    .ZN(_08833_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13059_ (.A1(net2083),
    .A2(_08621_),
    .Z(_08834_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13060_ (.A1(net2079),
    .A2(net2077),
    .A3(_08834_),
    .Z(_08835_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13061_ (.A1(_08465_),
    .A2(_08470_),
    .B(_08835_),
    .ZN(_08836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13062_ (.I(_00881_),
    .ZN(_08837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13063_ (.A1(_08833_),
    .A2(_08836_),
    .B(_08837_),
    .ZN(_08838_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _13064_ (.A1(_08837_),
    .A2(_08833_),
    .A3(_08836_),
    .Z(_08839_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13065_ (.A1(net1455),
    .A2(_08839_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13066_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_08840_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13067_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_08841_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13068_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_08842_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13069_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_08843_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13070_ (.I0(_08840_),
    .I1(_08841_),
    .I2(_08842_),
    .I3(_08843_),
    .S0(net1847),
    .S1(net1900),
    .Z(_08844_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13071_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S0(net1940),
    .S1(net1927),
    .Z(_08845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13072_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net1927),
    .Z(_08846_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13073_ (.A1(net1927),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .Z(_08847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13074_ (.I0(_08846_),
    .I1(_08847_),
    .S(net1853),
    .Z(_08848_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13075_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net1940),
    .S1(net1927),
    .Z(_08849_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13076_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net1940),
    .S1(net1927),
    .Z(_08850_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13077_ (.I0(_08845_),
    .I1(_08848_),
    .I2(_08849_),
    .I3(_08850_),
    .S0(net1847),
    .S1(net1902),
    .Z(_08851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13078_ (.I0(_08844_),
    .I1(_08851_),
    .S(net1863),
    .Z(_08852_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13080_ (.A1(net1960),
    .A2(_08551_),
    .ZN(_08854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13081_ (.A1(net2059),
    .A2(_08854_),
    .ZN(_08855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13082_ (.I0(net1768),
    .I1(_08855_),
    .S(net1795),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13083_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net2015),
    .S1(net1983),
    .Z(_08856_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13084_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net2015),
    .S1(net1983),
    .Z(_08857_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13085_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S0(net2015),
    .S1(net1983),
    .Z(_08858_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13086_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S0(net2015),
    .S1(net1983),
    .Z(_08859_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13087_ (.I0(_08856_),
    .I1(_08857_),
    .I2(_08858_),
    .I3(_08859_),
    .S0(net1877),
    .S1(net1866),
    .Z(_08860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13088_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net2134),
    .Z(_08861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13089_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .A2(_08657_),
    .B1(_08861_),
    .B2(net1986),
    .C(net1962),
    .ZN(_08862_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13090_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S0(net2134),
    .S1(net1985),
    .Z(_08863_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13091_ (.A1(net1877),
    .A2(_08863_),
    .B(net1866),
    .ZN(_08864_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13092_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net1989),
    .S1(net1983),
    .Z(_08865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13093_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net2134),
    .S1(net1983),
    .Z(_08866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13094_ (.I0(_08865_),
    .I1(_08866_),
    .S(net1877),
    .Z(_08867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13095_ (.A1(net1959),
    .A2(_08867_),
    .ZN(_08868_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13096_ (.A1(_08862_),
    .A2(_08864_),
    .B(_08868_),
    .C(net1842),
    .ZN(_08869_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13097_ (.A1(net1842),
    .A2(_08860_),
    .B(_08869_),
    .ZN(_08870_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13098_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1768),
    .ZN(_08871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13099_ (.A1(net2028),
    .A2(net1731),
    .B(_08871_),
    .ZN(_08872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13100_ (.I0(net2175),
    .I1(net2111),
    .S(_01264_),
    .Z(_08873_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13101_ (.A1(_08187_),
    .A2(_08872_),
    .B(_08873_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13102_ (.A1(\cs_registers_i.pc_id_i[18] ),
    .A2(net1801),
    .ZN(_08874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13103_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net1818),
    .ZN(_08875_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13104_ (.A1(net1742),
    .A2(net1731),
    .B1(_08874_),
    .B2(net1741),
    .C(_08875_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13105_ (.I(net1682),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13107_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net2182),
    .S1(net1924),
    .Z(_08877_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13108_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08878_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13109_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net2182),
    .S1(net1924),
    .Z(_08879_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13110_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net2182),
    .S1(net1924),
    .Z(_08880_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13111_ (.I0(_08877_),
    .I1(_08878_),
    .I2(_08879_),
    .I3(_08880_),
    .S0(net1851),
    .S1(net1900),
    .Z(_08881_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13112_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net1938),
    .S1(net1922),
    .Z(_08882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13113_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net1922),
    .Z(_08883_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13114_ (.A1(net1922),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .Z(_08884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13115_ (.I0(_08883_),
    .I1(_08884_),
    .S(net1854),
    .Z(_08885_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13116_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net1938),
    .S1(net1922),
    .Z(_08886_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13117_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net1938),
    .S1(net1922),
    .Z(_08887_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13118_ (.I0(_08882_),
    .I1(_08885_),
    .I2(_08886_),
    .I3(_08887_),
    .S0(net1851),
    .S1(net1900),
    .Z(_08888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13119_ (.I0(_08881_),
    .I1(_08888_),
    .S(net1860),
    .Z(_08889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13120_ (.A1(net1958),
    .A2(_08551_),
    .ZN(_08890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13121_ (.A1(net2060),
    .A2(_08890_),
    .ZN(_08891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13122_ (.I0(net1767),
    .I1(_08891_),
    .S(net1795),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13123_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S0(net2011),
    .S1(net1980),
    .Z(_08892_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13124_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S0(net2011),
    .S1(net1980),
    .Z(_08893_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13125_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net2011),
    .S1(net1980),
    .Z(_08894_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13126_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S0(net2011),
    .S1(net1980),
    .Z(_08895_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13127_ (.I0(_08892_),
    .I1(_08893_),
    .I2(_08894_),
    .I3(_08895_),
    .S0(net1878),
    .S1(net1866),
    .Z(_08896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13128_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net2193),
    .Z(_08897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13129_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A2(net1821),
    .B1(_08897_),
    .B2(net1982),
    .C(net1963),
    .ZN(_08898_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13130_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net2193),
    .S1(net1982),
    .Z(_08899_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13131_ (.A1(net1878),
    .A2(_08899_),
    .B(net1866),
    .ZN(_08900_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13132_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S0(net2008),
    .S1(net1976),
    .Z(_08901_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13133_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S0(net2008),
    .S1(net1976),
    .Z(_08902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13134_ (.I0(_08901_),
    .I1(_08902_),
    .S(net1878),
    .Z(_08903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13135_ (.A1(net1959),
    .A2(_08903_),
    .ZN(_08904_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13136_ (.A1(_08898_),
    .A2(_08900_),
    .B(_08904_),
    .C(net1843),
    .ZN(_08905_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13137_ (.A1(net1843),
    .A2(_08896_),
    .B(_08905_),
    .ZN(_08906_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13138_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1767),
    .ZN(_08907_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13139_ (.A1(net2028),
    .A2(net1730),
    .B(_08907_),
    .ZN(_08908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13140_ (.I0(net1693),
    .I1(net2111),
    .S(_01271_),
    .Z(_08909_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13141_ (.A1(_08187_),
    .A2(_08908_),
    .B(_08909_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13142_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(net1801),
    .ZN(_08910_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13143_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net1818),
    .ZN(_08911_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13144_ (.A1(net1742),
    .A2(net1730),
    .B1(_08910_),
    .B2(net1741),
    .C(_08911_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13145_ (.I(net1681),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13146_ (.I(_00893_),
    .ZN(_08912_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13147_ (.A1(_00889_),
    .A2(_00884_),
    .Z(_08913_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13148_ (.A1(_00888_),
    .A2(_08913_),
    .Z(_08914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13149_ (.A1(_00885_),
    .A2(net2108),
    .ZN(_08915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13150_ (.A1(net2287),
    .A2(_08828_),
    .B(_08915_),
    .ZN(_08916_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13151_ (.A1(_08914_),
    .A2(_08916_),
    .Z(_08917_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13152_ (.A1(_08912_),
    .A2(_08917_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13153_ (.A1(_08129_),
    .A2(_08170_),
    .B(_08502_),
    .C(_08184_),
    .ZN(_08918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13154_ (.A1(_08498_),
    .A2(_08500_),
    .Z(_08919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _13155_ (.A1(_00885_),
    .A2(net2194),
    .ZN(_08920_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _13156_ (.A1(_08920_),
    .A2(_08737_),
    .ZN(_08921_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13157_ (.A1(_08919_),
    .A2(_08921_),
    .Z(_08922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13158_ (.A1(net2076),
    .A2(_00872_),
    .B(_00876_),
    .ZN(_08923_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13159_ (.A1(_08923_),
    .A2(_08837_),
    .B(_08820_),
    .ZN(_08924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13160_ (.A1(_00885_),
    .A2(_08924_),
    .B(_00884_),
    .ZN(_08925_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13161_ (.A1(_08920_),
    .A2(_08740_),
    .A3(_08739_),
    .B(_08925_),
    .ZN(_08926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13162_ (.A1(_08918_),
    .A2(_08922_),
    .B(_08926_),
    .ZN(_08927_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13163_ (.A1(_08927_),
    .A2(net2107),
    .Z(_08928_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13164_ (.I(_08928_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13165_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08929_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13166_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08930_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13167_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08931_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13168_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08932_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13169_ (.I0(_08929_),
    .I1(_08930_),
    .I2(_08931_),
    .I3(_08932_),
    .S0(net1851),
    .S1(net1900),
    .Z(_08933_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13170_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net1938),
    .S1(net1924),
    .Z(_08934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13171_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net1922),
    .Z(_08935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13172_ (.A1(net1922),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .Z(_08936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13173_ (.I0(_08935_),
    .I1(_08936_),
    .S(net1854),
    .Z(_08937_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13174_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net1938),
    .S1(net1922),
    .Z(_08938_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13175_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net1938),
    .S1(net1922),
    .Z(_08939_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13176_ (.I0(_08934_),
    .I1(_08937_),
    .I2(_08938_),
    .I3(_08939_),
    .S0(net1851),
    .S1(net1900),
    .Z(_08940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13177_ (.I0(_08933_),
    .I1(_08940_),
    .S(net1860),
    .Z(_08941_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13178_ (.A1(_08546_),
    .A2(_07861_),
    .Z(_08942_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13180_ (.A1(net1855),
    .A2(net2054),
    .B(_08942_),
    .ZN(_08944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13181_ (.I0(net1766),
    .I1(_08944_),
    .S(net1795),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13182_ (.I(_08941_),
    .ZN(_08945_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13183_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net2008),
    .S1(net1976),
    .Z(_08946_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13184_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net2008),
    .S1(net1976),
    .Z(_08947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13185_ (.I0(_08946_),
    .I1(_08947_),
    .S(net1878),
    .Z(_08948_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13186_ (.A1(net1959),
    .A2(_08948_),
    .Z(_08949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13187_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net2193),
    .Z(_08950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13188_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .A2(net1821),
    .B1(_08950_),
    .B2(net1976),
    .ZN(_08951_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13189_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net2193),
    .S1(net1979),
    .Z(_08952_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13190_ (.A1(net1878),
    .A2(_08952_),
    .B(net1866),
    .ZN(_08953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13191_ (.A1(net1878),
    .A2(_08951_),
    .B(_08953_),
    .ZN(_08954_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13192_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net2010),
    .S1(net1979),
    .Z(_08955_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13193_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net2010),
    .S1(net1979),
    .Z(_08956_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13194_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S0(net2010),
    .S1(net1979),
    .Z(_08957_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13195_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S0(net2193),
    .S1(net1979),
    .Z(_08958_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13196_ (.I0(_08955_),
    .I1(_08956_),
    .I2(_08957_),
    .I3(_08958_),
    .S0(net1878),
    .S1(net1866),
    .Z(_08959_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13197_ (.A1(net1843),
    .A2(_08959_),
    .ZN(_08960_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13198_ (.I(_08960_),
    .ZN(_08961_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13199_ (.A1(net1958),
    .A2(net1810),
    .A3(net1765),
    .B(net1764),
    .ZN(_08962_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13200_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .B2(net1824),
    .ZN(_08963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13201_ (.A1(_08228_),
    .A2(net1729),
    .B1(net1728),
    .B2(net2028),
    .C(_08963_),
    .ZN(_08964_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1550 (.I(_09687_),
    .Z(net1549));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13203_ (.I0(net1693),
    .I1(net1694),
    .S(_01278_),
    .Z(_08966_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13204_ (.A1(_08187_),
    .A2(_08964_),
    .B(_08966_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13205_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(net1801),
    .ZN(_08967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13206_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net1818),
    .ZN(_08968_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _13207_ (.A1(net2160),
    .A2(net1742),
    .B1(_08967_),
    .B2(net1741),
    .C(_08968_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13208_ (.I(net2135),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13209_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08969_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13210_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08970_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13211_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08971_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13212_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08972_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13213_ (.I0(_08969_),
    .I1(_08970_),
    .I2(_08971_),
    .I3(_08972_),
    .S0(net1850),
    .S1(net1901),
    .Z(_08973_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13214_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net1949),
    .S1(net2089),
    .Z(_08974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13215_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net2089),
    .Z(_08975_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13216_ (.A1(net2089),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .Z(_08976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13217_ (.I0(_08975_),
    .I1(_08976_),
    .S(net1853),
    .Z(_08977_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13218_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08978_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13219_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net1949),
    .S1(net1911),
    .Z(_08979_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13220_ (.I0(_08974_),
    .I1(_08977_),
    .I2(_08978_),
    .I3(_08979_),
    .S0(net1850),
    .S1(net1901),
    .Z(_08980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13221_ (.I0(_08973_),
    .I1(_08980_),
    .S(net1863),
    .Z(_08981_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1548 (.I(_00452_),
    .Z(net1547));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13223_ (.A1(net1908),
    .A2(_08547_),
    .ZN(_08983_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13224_ (.A1(net2057),
    .A2(_08983_),
    .ZN(_08984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13225_ (.I0(net1763),
    .I1(_08984_),
    .S(net1795),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13226_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net1990),
    .S1(net1962),
    .Z(_08985_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13227_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .S0(net1990),
    .S1(net1962),
    .Z(_08986_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13228_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net1990),
    .S1(net1962),
    .Z(_08987_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13229_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .S0(net1990),
    .S1(net1962),
    .Z(_08988_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13230_ (.I0(_08985_),
    .I1(_08986_),
    .I2(_08987_),
    .I3(_08988_),
    .S0(net1874),
    .S1(net1866),
    .Z(_08989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13231_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net1990),
    .Z(_08990_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13232_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A2(net1820),
    .B1(_08990_),
    .B2(net1970),
    .C(net1962),
    .ZN(_08991_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13233_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net1990),
    .S1(net1970),
    .Z(_08992_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13234_ (.A1(net1881),
    .A2(_08992_),
    .B(net1866),
    .ZN(_08993_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13235_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_08994_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13236_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_08995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13237_ (.I0(_08994_),
    .I1(_08995_),
    .S(net1881),
    .Z(_08996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13238_ (.A1(net1961),
    .A2(_08996_),
    .ZN(_08997_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13239_ (.A1(_08991_),
    .A2(_08993_),
    .B(_08997_),
    .C(net1842),
    .ZN(_08998_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13240_ (.A1(net1842),
    .A2(_08989_),
    .B(_08998_),
    .ZN(_08999_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1547 (.I(_00659_),
    .Z(net1546));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13242_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1763),
    .ZN(_09001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13243_ (.A1(net2028),
    .A2(net1727),
    .B(_09001_),
    .ZN(_09002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13244_ (.I0(net2175),
    .I1(net1694),
    .S(_01285_),
    .Z(_09003_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13245_ (.A1(net1783),
    .A2(_09002_),
    .B(_09003_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13246_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(net1801),
    .ZN(_09004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13247_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net1818),
    .ZN(_09005_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13248_ (.A1(net1742),
    .A2(net1727),
    .B1(_09004_),
    .B2(net1741),
    .C(_09005_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13249_ (.I(net1680),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13250_ (.A1(_00885_),
    .A2(net2172),
    .Z(_09006_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13251_ (.A1(_00897_),
    .A2(_00901_),
    .Z(_09007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13252_ (.A1(_00893_),
    .A2(_09007_),
    .Z(_09008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13253_ (.A1(_09006_),
    .A2(_09008_),
    .ZN(_09009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13254_ (.A1(_08819_),
    .A2(_08828_),
    .B(_09009_),
    .ZN(_09010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13255_ (.A1(_08914_),
    .A2(_09008_),
    .Z(_09011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13256_ (.A1(_00897_),
    .A2(_00892_),
    .Z(_09012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13257_ (.A1(_00896_),
    .A2(_09012_),
    .Z(_09013_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13258_ (.A1(_00901_),
    .A2(_09013_),
    .Z(_09014_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13259_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09014_),
    .Z(_09015_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13260_ (.A1(_00893_),
    .A2(_00897_),
    .Z(_09016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13261_ (.A1(_08917_),
    .A2(_09016_),
    .B(_09013_),
    .C(_00901_),
    .ZN(_09017_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13262_ (.A1(_09015_),
    .A2(net1434),
    .ZN(net167));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13263_ (.A1(_08919_),
    .A2(_08834_),
    .A3(_08817_),
    .A4(_09006_),
    .ZN(_09018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13264_ (.A1(net2107),
    .A2(_08926_),
    .B(_00892_),
    .C(_00888_),
    .ZN(_09019_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13265_ (.A1(_00897_),
    .A2(_09019_),
    .Z(_09020_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13266_ (.A1(net2123),
    .A2(_09018_),
    .B(_09020_),
    .ZN(_09021_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13267_ (.A1(_08912_),
    .A2(_00897_),
    .Z(_09022_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13268_ (.A1(net2123),
    .A2(_09018_),
    .A3(_09022_),
    .Z(_09023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13269_ (.A1(net2108),
    .A2(_08926_),
    .B(_00888_),
    .ZN(_09024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13270_ (.I(_00892_),
    .ZN(_09025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13271_ (.A1(_08912_),
    .A2(_09025_),
    .ZN(_09026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13272_ (.I0(_09025_),
    .I1(_09026_),
    .S(_00897_),
    .Z(_09027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13273_ (.A1(_09024_),
    .A2(_09022_),
    .B(_09027_),
    .ZN(_09028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13274_ (.I(_09028_),
    .ZN(_09029_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13275_ (.A1(_09021_),
    .A2(_09023_),
    .A3(_09029_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13276_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net1952),
    .S1(net1918),
    .Z(_09030_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13277_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S0(net1952),
    .S1(net1918),
    .Z(_09031_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13278_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net2114),
    .S1(net1918),
    .Z(_09032_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13279_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net1952),
    .S1(net1918),
    .Z(_09033_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13280_ (.I0(_09030_),
    .I1(_09031_),
    .I2(_09032_),
    .I3(_09033_),
    .S0(net1847),
    .S1(net1902),
    .Z(_09034_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13281_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net1953),
    .S1(net1918),
    .Z(_09035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13282_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net1918),
    .Z(_09036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13283_ (.A1(net1918),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .Z(_09037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13284_ (.I0(_09036_),
    .I1(_09037_),
    .S(net1853),
    .Z(_09038_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13285_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net1951),
    .S1(net1918),
    .Z(_09039_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13286_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net1951),
    .S1(net1918),
    .Z(_09040_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13287_ (.I0(_09035_),
    .I1(_09038_),
    .I2(_09039_),
    .I3(_09040_),
    .S0(net1847),
    .S1(net1902),
    .Z(_09041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13288_ (.I0(_09034_),
    .I1(_09041_),
    .S(net1863),
    .Z(_09042_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13289_ (.A1(net1848),
    .A2(net2054),
    .B(_08942_),
    .ZN(_09043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13290_ (.I0(net1762),
    .I1(_09043_),
    .S(net1795),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1546 (.I(_00490_),
    .Z(net1545));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13292_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net2166),
    .S1(net1963),
    .Z(_09045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13293_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .S0(net2166),
    .S1(net1963),
    .Z(_09046_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13294_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net2134),
    .S1(net1963),
    .Z(_09047_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13295_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .S0(net2134),
    .S1(net1963),
    .Z(_09048_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13296_ (.I0(_09045_),
    .I1(_09046_),
    .I2(_09047_),
    .I3(_09048_),
    .S0(net1874),
    .S1(net1866),
    .Z(_09049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13297_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net2166),
    .Z(_09050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13298_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A2(_08657_),
    .B1(_09050_),
    .B2(net1973),
    .C(net1962),
    .ZN(_09051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13299_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net2166),
    .S1(net1973),
    .Z(_09052_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13300_ (.A1(net1881),
    .A2(_09052_),
    .B(net1866),
    .ZN(_09053_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13301_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net1990),
    .S1(net1973),
    .Z(_09054_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13302_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net1990),
    .S1(net1973),
    .Z(_09055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13303_ (.I0(_09054_),
    .I1(_09055_),
    .S(net1881),
    .Z(_09056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13304_ (.A1(net1961),
    .A2(_09056_),
    .ZN(_09057_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13305_ (.A1(_09051_),
    .A2(_09053_),
    .B(_09057_),
    .C(net1842),
    .ZN(_09058_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13306_ (.A1(net1843),
    .A2(_09049_),
    .B(_09058_),
    .ZN(_09059_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1545 (.I(_00684_),
    .Z(net1544));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1549 (.I(_09702_),
    .Z(net1548));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13309_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1762),
    .ZN(_09062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13310_ (.A1(net2028),
    .A2(net1726),
    .B(_09062_),
    .ZN(_09063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13311_ (.I0(net1693),
    .I1(net1694),
    .S(_01292_),
    .Z(_09064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13312_ (.A1(net1783),
    .A2(_09063_),
    .B(_09064_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13313_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(net1801),
    .ZN(_09065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13314_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net1818),
    .ZN(_09066_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13315_ (.A1(net1742),
    .A2(net1726),
    .B1(_09065_),
    .B2(net1741),
    .C(_09066_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13316_ (.I(net1679),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13317_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net2114),
    .S1(net1930),
    .Z(_09067_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13318_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net2114),
    .S1(net1930),
    .Z(_09068_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13319_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net2114),
    .S1(net1930),
    .Z(_09069_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13320_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net2114),
    .S1(net1930),
    .Z(_09070_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13321_ (.I0(_09067_),
    .I1(_09068_),
    .I2(_09069_),
    .I3(_09070_),
    .S0(net1847),
    .S1(net1902),
    .Z(_09071_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13322_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net1955),
    .S1(net1930),
    .Z(_09072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13323_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net1927),
    .Z(_09073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13324_ (.A1(net1927),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .Z(_09074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13325_ (.I0(_09073_),
    .I1(_09074_),
    .S(net1853),
    .Z(_09075_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13326_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net2114),
    .S1(net1930),
    .Z(_09076_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13327_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net1955),
    .S1(net1930),
    .Z(_09077_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13328_ (.I0(_09072_),
    .I1(_09075_),
    .I2(_09076_),
    .I3(_09077_),
    .S0(net1847),
    .S1(net1902),
    .Z(_09078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13329_ (.I0(_09071_),
    .I1(_09078_),
    .S(net1863),
    .Z(_09079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13330_ (.A1(net1858),
    .A2(net2054),
    .B(_08942_),
    .ZN(_09080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13331_ (.I0(net1761),
    .I1(_09080_),
    .S(net1795),
    .Z(_01299_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13332_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net1998),
    .S1(net1988),
    .Z(_09081_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13333_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net1998),
    .S1(net1988),
    .Z(_09082_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13334_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net1998),
    .S1(net1988),
    .Z(_09083_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13335_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net1998),
    .S1(net1988),
    .Z(_09084_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13336_ (.I0(_09081_),
    .I1(_09082_),
    .I2(_09083_),
    .I3(_09084_),
    .S0(net1877),
    .S1(net1866),
    .Z(_09085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13337_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net1998),
    .Z(_09086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13338_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .A2(net1821),
    .B1(_09086_),
    .B2(net1986),
    .C(net1962),
    .ZN(_09087_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13339_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net1998),
    .S1(net1985),
    .Z(_09088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13340_ (.A1(net1879),
    .A2(_09088_),
    .B(net1866),
    .ZN(_09089_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13341_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net2165),
    .S1(net1986),
    .Z(_09090_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13342_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net2165),
    .S1(net1986),
    .Z(_09091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13343_ (.I0(_09090_),
    .I1(_09091_),
    .S(net1879),
    .Z(_09092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13344_ (.A1(net1959),
    .A2(_09092_),
    .ZN(_09093_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13345_ (.A1(_09087_),
    .A2(_09089_),
    .B(_09093_),
    .C(net1842),
    .ZN(_09094_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13346_ (.A1(net1842),
    .A2(_09085_),
    .B(_09094_),
    .ZN(_09095_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13347_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1761),
    .ZN(_09096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13348_ (.A1(net2028),
    .A2(net1725),
    .B(_09096_),
    .ZN(_09097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13349_ (.I0(net1693),
    .I1(net2111),
    .S(_01299_),
    .Z(_09098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13350_ (.A1(net1783),
    .A2(_09097_),
    .B(_09098_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13351_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(net1801),
    .ZN(_09099_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13352_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net1818),
    .ZN(_09100_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13353_ (.A1(net1742),
    .A2(net1725),
    .B1(_09099_),
    .B2(net1741),
    .C(_09100_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13354_ (.I(net1678),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13355_ (.I(_00904_),
    .ZN(_09101_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13356_ (.A1(_00900_),
    .A2(_09014_),
    .Z(_09102_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13357_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09102_),
    .B(net2186),
    .ZN(_09103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _13358_ (.I(_00909_),
    .ZN(_09104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13359_ (.A1(_09101_),
    .A2(_09103_),
    .B(_09104_),
    .ZN(_09105_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13360_ (.A1(_09104_),
    .A2(_09101_),
    .A3(_09103_),
    .Z(_09106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13361_ (.A1(_09105_),
    .A2(_09106_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13362_ (.A1(net2107),
    .A2(_09008_),
    .Z(_09107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13363_ (.A1(_08919_),
    .A2(_08921_),
    .A3(_09107_),
    .Z(_09108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13364_ (.A1(_08924_),
    .A2(_09006_),
    .B(_08914_),
    .ZN(_09109_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13365_ (.A1(_08912_),
    .A2(_09109_),
    .B(_09025_),
    .ZN(_09110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13366_ (.A1(_00901_),
    .A2(_00896_),
    .Z(_09111_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13367_ (.A1(_00900_),
    .A2(_09111_),
    .Z(_09112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13368_ (.A1(_09007_),
    .A2(_09110_),
    .B(_09112_),
    .ZN(_09113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13369_ (.A1(net2107),
    .A2(_09008_),
    .ZN(_09114_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13370_ (.A1(_08741_),
    .A2(_08920_),
    .A3(_09114_),
    .Z(_09115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13371_ (.A1(_09113_),
    .A2(_09115_),
    .ZN(_09116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _13372_ (.A1(_08918_),
    .A2(_09108_),
    .B(_09116_),
    .ZN(_09117_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13373_ (.A1(net2186),
    .A2(_09117_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13374_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net1948),
    .S1(net1911),
    .Z(_09118_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1544 (.I(_04411_),
    .Z(net1543));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13376_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S0(net1948),
    .S1(net1911),
    .Z(_09120_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13377_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net1948),
    .S1(net1911),
    .Z(_09121_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13378_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .S0(net1948),
    .S1(net1911),
    .Z(_09122_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13379_ (.I0(_09118_),
    .I1(_09120_),
    .I2(_09121_),
    .I3(_09122_),
    .S0(net1847),
    .S1(net1901),
    .Z(_09123_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13380_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S0(net1953),
    .S1(net2089),
    .Z(_09124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13381_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net2089),
    .Z(_09125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13382_ (.A1(net2089),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .Z(_09126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13383_ (.I0(_09125_),
    .I1(_09126_),
    .S(net1853),
    .Z(_09127_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13384_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net1953),
    .S1(net2089),
    .Z(_09128_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13385_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net1953),
    .S1(net2089),
    .Z(_09129_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13386_ (.I0(_09124_),
    .I1(_09127_),
    .I2(_09128_),
    .I3(_09129_),
    .S0(net1847),
    .S1(net1901),
    .Z(_09130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13387_ (.I0(_09123_),
    .I1(_09130_),
    .S(net1862),
    .Z(_09131_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13388_ (.A1(net1860),
    .A2(net2054),
    .B(_08942_),
    .ZN(_09132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13389_ (.I0(net1760),
    .I1(_09132_),
    .S(net1795),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13391_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net1992),
    .S1(net1962),
    .Z(_09134_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13392_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .S0(net1992),
    .S1(net1962),
    .Z(_09135_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13393_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net1992),
    .S1(net1962),
    .Z(_09136_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13394_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .S0(net1992),
    .S1(net1962),
    .Z(_09137_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13395_ (.I0(_09134_),
    .I1(_09135_),
    .I2(_09136_),
    .I3(_09137_),
    .S0(net1873),
    .S1(net1866),
    .Z(_09138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13396_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net1990),
    .Z(_09139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13397_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A2(net1820),
    .B1(_09139_),
    .B2(net1970),
    .C(net1962),
    .ZN(_09140_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13398_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S0(net1990),
    .S1(net1970),
    .Z(_09141_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13399_ (.A1(net1881),
    .A2(_09141_),
    .B(net1866),
    .ZN(_09142_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13400_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net1990),
    .S1(net1970),
    .Z(_09143_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13401_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net1990),
    .S1(net1968),
    .Z(_09144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13402_ (.I0(_09143_),
    .I1(_09144_),
    .S(net1881),
    .Z(_09145_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13403_ (.A1(net1961),
    .A2(_09145_),
    .ZN(_09146_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13404_ (.A1(_09140_),
    .A2(_09142_),
    .B(_09146_),
    .C(net1842),
    .ZN(_09147_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13405_ (.A1(net1842),
    .A2(_09138_),
    .B(_09147_),
    .ZN(_09148_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13406_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1760),
    .ZN(_09149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13407_ (.A1(net2028),
    .A2(net1723),
    .B(_09149_),
    .ZN(_09150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13408_ (.I0(net1693),
    .I1(net2111),
    .S(_01306_),
    .Z(_09151_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13409_ (.A1(net1783),
    .A2(_09150_),
    .B(_09151_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13410_ (.A1(\cs_registers_i.pc_id_i[24] ),
    .A2(net1801),
    .ZN(_09152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13411_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net1818),
    .ZN(_09153_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13412_ (.A1(net1742),
    .A2(net1723),
    .B1(_09152_),
    .B2(net1741),
    .C(_09153_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13413_ (.I(net1677),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13414_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09154_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13415_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09155_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13416_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09156_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13417_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09157_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13418_ (.I0(_09154_),
    .I1(_09155_),
    .I2(_09156_),
    .I3(_09157_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09158_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13419_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13420_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net1927),
    .Z(_09160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13421_ (.A1(net1927),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .Z(_09161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13422_ (.I0(_09160_),
    .I1(_09161_),
    .S(net1854),
    .Z(_09162_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13423_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09163_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13424_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09164_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13425_ (.I0(_09159_),
    .I1(_09162_),
    .I2(_09163_),
    .I3(_09164_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13426_ (.I0(_09158_),
    .I1(_09165_),
    .S(net1860),
    .Z(_09166_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13427_ (.A1(_07833_),
    .A2(net2054),
    .B(_08942_),
    .ZN(_09167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13428_ (.I0(net1759),
    .I1(_09167_),
    .S(net1795),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13429_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S0(net2014),
    .S1(net1963),
    .Z(_09168_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13430_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .S0(net2014),
    .S1(net1963),
    .Z(_09169_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13431_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S0(net2014),
    .S1(net1963),
    .Z(_09170_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13432_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .S0(net2014),
    .S1(net1963),
    .Z(_09171_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13433_ (.I0(_09168_),
    .I1(_09169_),
    .I2(_09170_),
    .I3(_09171_),
    .S0(net1875),
    .S1(net1866),
    .Z(_09172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13434_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net2014),
    .Z(_09173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13435_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A2(net1821),
    .B1(_09173_),
    .B2(net1984),
    .C(net1963),
    .ZN(_09174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13436_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net2014),
    .S1(net1984),
    .Z(_09175_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13437_ (.A1(net1877),
    .A2(_09175_),
    .B(net1866),
    .ZN(_09176_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13438_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S0(net2013),
    .S1(net1984),
    .Z(_09177_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13439_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S0(net2014),
    .S1(net1984),
    .Z(_09178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13440_ (.I0(_09177_),
    .I1(_09178_),
    .S(net1877),
    .Z(_09179_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13441_ (.A1(net1959),
    .A2(_09179_),
    .ZN(_09180_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13442_ (.A1(_09174_),
    .A2(_09176_),
    .B(_09180_),
    .C(net1843),
    .ZN(_09181_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13443_ (.A1(net1843),
    .A2(_09172_),
    .B(_09181_),
    .ZN(_09182_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13444_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .B2(_08197_),
    .C1(_08200_),
    .C2(net1759),
    .ZN(_09183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13445_ (.A1(net2028),
    .A2(net1722),
    .B(_09183_),
    .ZN(_09184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13446_ (.I0(net2175),
    .I1(net2111),
    .S(_01313_),
    .Z(_09185_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13447_ (.A1(net1783),
    .A2(_09184_),
    .B(_09185_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13448_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(net1801),
    .ZN(_09186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13449_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net1818),
    .ZN(_09187_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _13450_ (.A1(net1742),
    .A2(net1722),
    .B1(_09186_),
    .B2(net1741),
    .C(_09187_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13451_ (.I(_01312_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13452_ (.A1(_00905_),
    .A2(_00900_),
    .B(_00904_),
    .ZN(_09188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13453_ (.I(_00908_),
    .ZN(_09189_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13454_ (.A1(_09104_),
    .A2(_09188_),
    .B(_09189_),
    .ZN(_09190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13455_ (.A1(_09190_),
    .A2(_00913_),
    .B(_00912_),
    .ZN(_09191_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13456_ (.A1(_00905_),
    .A2(_00909_),
    .A3(_00913_),
    .Z(_09192_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13457_ (.A1(_00917_),
    .A2(_09192_),
    .ZN(_09193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13458_ (.I(_00917_),
    .ZN(_09194_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13459_ (.A1(_09194_),
    .A2(_09191_),
    .ZN(_09195_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13460_ (.A1(net2129),
    .A2(_09193_),
    .B(_09195_),
    .ZN(_09196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _13461_ (.A1(_00917_),
    .A2(_09192_),
    .Z(_09197_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13462_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09014_),
    .B(_09197_),
    .ZN(_09198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13463_ (.A1(_09194_),
    .A2(net2129),
    .ZN(_09199_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13464_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09014_),
    .A4(_09199_),
    .Z(_09200_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13465_ (.A1(_09196_),
    .A2(_09198_),
    .A3(_09200_),
    .Z(net171));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13466_ (.A1(net2123),
    .A2(_09018_),
    .B(_09019_),
    .ZN(_09201_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13467_ (.A1(net2186),
    .A2(_09007_),
    .A3(_09026_),
    .Z(_09202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13468_ (.A1(net2186),
    .A2(_09112_),
    .B(_00904_),
    .ZN(_09203_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13469_ (.A1(_00913_),
    .A2(_09189_),
    .A3(_09203_),
    .ZN(_09204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13470_ (.A1(_09201_),
    .A2(_09202_),
    .B(_09204_),
    .ZN(_09205_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13471_ (.I(_00913_),
    .ZN(_09206_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13472_ (.A1(_00909_),
    .A2(_09206_),
    .A3(_09201_),
    .A4(_09202_),
    .Z(_09207_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13473_ (.A1(_09104_),
    .A2(_00913_),
    .A3(_09203_),
    .ZN(_09208_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13474_ (.A1(_09104_),
    .A2(_00913_),
    .Z(_09209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13475_ (.I0(_09206_),
    .I1(_09209_),
    .S(_09189_),
    .Z(_09210_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13476_ (.A1(_09207_),
    .A2(_09205_),
    .A3(_09208_),
    .A4(_09210_),
    .Z(net170));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13477_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S0(net2182),
    .S1(net1925),
    .Z(_09211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13478_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S0(net2182),
    .S1(net1925),
    .Z(_09212_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13479_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net2182),
    .S1(net1924),
    .Z(_09213_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13480_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net2182),
    .S1(net1924),
    .Z(_09214_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13481_ (.I0(_09211_),
    .I1(_09212_),
    .I2(_09213_),
    .I3(_09214_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09215_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13482_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net2182),
    .S1(net1925),
    .Z(_09216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13483_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net1922),
    .Z(_09217_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13484_ (.A1(net1922),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .Z(_09218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13485_ (.I0(_09217_),
    .I1(_09218_),
    .S(net1854),
    .Z(_09219_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13486_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S0(net2182),
    .S1(net1925),
    .Z(_09220_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13487_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S0(net1942),
    .S1(net1925),
    .Z(_09221_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13488_ (.I0(_09216_),
    .I1(_09219_),
    .I2(_09220_),
    .I3(_09221_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13489_ (.I0(_09215_),
    .I1(_09222_),
    .S(net1860),
    .Z(_09223_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13490_ (.A1(_07860_),
    .A2(net2054),
    .B(net2056),
    .ZN(_09224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13491_ (.I0(net1758),
    .I1(_09224_),
    .S(net1795),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13492_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net2012),
    .S1(net1981),
    .Z(_09225_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13493_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net2012),
    .S1(net1981),
    .Z(_09226_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13494_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S0(net2012),
    .S1(net1981),
    .Z(_09227_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13495_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S0(net2012),
    .S1(net1981),
    .Z(_09228_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13496_ (.I0(_09225_),
    .I1(_09226_),
    .I2(_09227_),
    .I3(_09228_),
    .S0(net1878),
    .S1(net1866),
    .Z(_09229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13497_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net2012),
    .Z(_09230_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13498_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .A2(net1821),
    .B1(_09230_),
    .B2(net1982),
    .C(net1963),
    .ZN(_09231_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13499_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net2012),
    .S1(net1981),
    .Z(_09232_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13500_ (.A1(net1878),
    .A2(_09232_),
    .B(net1866),
    .ZN(_09233_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13501_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S0(net2012),
    .S1(net1980),
    .Z(_09234_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13502_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S0(net2012),
    .S1(net1982),
    .Z(_09235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13503_ (.I0(_09234_),
    .I1(_09235_),
    .S(net1878),
    .Z(_09236_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13504_ (.A1(net1959),
    .A2(_09236_),
    .ZN(_09237_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13505_ (.A1(_09231_),
    .A2(_09233_),
    .B(_09237_),
    .C(net1843),
    .ZN(_09238_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13506_ (.A1(net1843),
    .A2(_09229_),
    .B(_09238_),
    .ZN(_09239_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13507_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1758),
    .ZN(_09240_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13508_ (.A1(net2028),
    .A2(net1721),
    .B(_09240_),
    .ZN(_09241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13509_ (.I0(net2175),
    .I1(net2111),
    .S(_01320_),
    .Z(_09242_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13510_ (.A1(_08187_),
    .A2(_09241_),
    .B(_09242_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13511_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(net1801),
    .ZN(_09243_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13512_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net1818),
    .ZN(_09244_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _13513_ (.A1(net1742),
    .A2(net1721),
    .B1(_09243_),
    .B2(net1741),
    .C(_09244_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13514_ (.I(_01319_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13515_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09245_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13516_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09246_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13518_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09248_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13519_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net2112),
    .S1(net1927),
    .Z(_09249_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13520_ (.I0(_09245_),
    .I1(_09246_),
    .I2(_09248_),
    .I3(_09249_),
    .S0(net1847),
    .S1(net1900),
    .Z(_09250_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13521_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net1942),
    .S1(net1927),
    .Z(_09251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13522_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net1927),
    .Z(_09252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13523_ (.A1(net1927),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .Z(_09253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13524_ (.I0(_09252_),
    .I1(_09253_),
    .S(net1853),
    .Z(_09254_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13525_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net1941),
    .S1(net1927),
    .Z(_09255_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13526_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net1941),
    .S1(net1927),
    .Z(_09256_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13527_ (.I0(_09251_),
    .I1(_09254_),
    .I2(_09255_),
    .I3(_09256_),
    .S0(net1847),
    .S1(net1900),
    .Z(_09257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13528_ (.I0(_09250_),
    .I1(_09257_),
    .S(net1863),
    .Z(_09258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13529_ (.A1(net1896),
    .A2(_08547_),
    .ZN(_09259_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13530_ (.A1(net2057),
    .A2(_09259_),
    .ZN(_09260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13531_ (.I0(net1757),
    .I1(_09260_),
    .S(net1795),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13532_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net2014),
    .S1(net1985),
    .Z(_09261_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13533_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net2014),
    .S1(net1985),
    .Z(_09262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13534_ (.I0(_09261_),
    .I1(_09262_),
    .S(net1879),
    .Z(_09263_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13535_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net2014),
    .S1(net1962),
    .Z(_09264_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13536_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .S0(net2014),
    .S1(net1962),
    .Z(_09265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13537_ (.I0(_09264_),
    .I1(_09265_),
    .S(net1875),
    .Z(_09266_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13538_ (.A1(net1822),
    .A2(_09263_),
    .B1(_09266_),
    .B2(_08589_),
    .ZN(_09267_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13539_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net2014),
    .S1(net1987),
    .Z(_09268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13540_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net2014),
    .Z(_09269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13541_ (.A1(net2014),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .Z(_09270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13542_ (.I0(_09269_),
    .I1(_09270_),
    .S(net1875),
    .Z(_09271_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13543_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net2014),
    .S1(net1984),
    .Z(_09272_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13544_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net2014),
    .S1(net1985),
    .Z(_09273_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13545_ (.I0(_09268_),
    .I1(_09271_),
    .I2(_09272_),
    .I3(_09273_),
    .S0(net1877),
    .S1(net1959),
    .Z(_09274_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13546_ (.A1(net1842),
    .A2(_09274_),
    .ZN(_09275_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13547_ (.A1(_09267_),
    .A2(_09275_),
    .Z(_09276_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13548_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1757),
    .ZN(_09277_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13549_ (.A1(net2028),
    .A2(net1720),
    .B(_09277_),
    .ZN(_09278_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1543 (.I(_06192_),
    .Z(net1542));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13551_ (.I0(net2175),
    .I1(net2111),
    .S(_01327_),
    .Z(_09280_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13552_ (.A1(_08187_),
    .A2(_09278_),
    .B(_09280_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13553_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(net1801),
    .ZN(_09281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13554_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net1818),
    .ZN(_09282_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_4 _13555_ (.A1(net1742),
    .A2(net1720),
    .B1(_09281_),
    .B2(net1741),
    .C(_09282_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13556_ (.I(_01326_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13557_ (.A1(_00916_),
    .A2(_00920_),
    .A3(_09014_),
    .A4(_09195_),
    .Z(_09283_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13558_ (.A1(_00916_),
    .A2(_00920_),
    .A3(_09195_),
    .A4(_09197_),
    .Z(_09284_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13559_ (.I(_00921_),
    .ZN(_09285_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13560_ (.I(_00920_),
    .ZN(_09286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13561_ (.A1(_09285_),
    .A2(_09286_),
    .ZN(_09287_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13562_ (.A1(_09284_),
    .A2(_09287_),
    .Z(_09288_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13563_ (.A1(_09010_),
    .A2(_09011_),
    .A3(_09283_),
    .B(_09288_),
    .ZN(_09289_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _13564_ (.A1(_00925_),
    .A2(_09289_),
    .ZN(net173));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13565_ (.A1(net2074),
    .A2(_08920_),
    .ZN(_09290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13566_ (.A1(_08919_),
    .A2(_08921_),
    .B(_09290_),
    .ZN(_09291_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _13567_ (.A1(net2074),
    .A2(_08920_),
    .B(_08502_),
    .ZN(_09292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13568_ (.A1(_08215_),
    .A2(net2121),
    .B(_09292_),
    .C(_08403_),
    .ZN(_09293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13569_ (.A1(_00909_),
    .A2(_00904_),
    .B(_00908_),
    .ZN(_09294_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13570_ (.I(_00912_),
    .ZN(_09295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13571_ (.A1(_09206_),
    .A2(_09294_),
    .B(_09295_),
    .ZN(_09296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13572_ (.A1(_00917_),
    .A2(_09296_),
    .B(_00916_),
    .ZN(_09297_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13573_ (.A1(_09285_),
    .A2(_09113_),
    .A3(_09297_),
    .Z(_09298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13574_ (.A1(_09291_),
    .A2(_09293_),
    .B(_09298_),
    .ZN(_09299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13575_ (.A1(_09107_),
    .A2(_09197_),
    .ZN(_09300_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _13576_ (.A1(_09285_),
    .A2(_09291_),
    .A3(_09293_),
    .A4(_09300_),
    .Z(_09301_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13577_ (.A1(_00917_),
    .A2(_09192_),
    .ZN(_09302_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13578_ (.A1(_09285_),
    .A2(_09302_),
    .Z(_09303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13579_ (.I0(_00921_),
    .I1(_09303_),
    .S(_09297_),
    .Z(_09304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13580_ (.A1(_00921_),
    .A2(_09197_),
    .Z(_09305_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13581_ (.A1(_09285_),
    .A2(_09114_),
    .A3(_09297_),
    .Z(_09306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13582_ (.I0(_09305_),
    .I1(_09306_),
    .S(net2085),
    .Z(_09307_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13583_ (.A1(_09304_),
    .A2(_09307_),
    .ZN(_09308_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _13584_ (.A1(_09299_),
    .A2(_09308_),
    .A3(_09301_),
    .ZN(_09309_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13585_ (.I(_09309_),
    .ZN(net172));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13586_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net1937),
    .S1(net1923),
    .Z(_09310_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13587_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S0(net1937),
    .S1(net1923),
    .Z(_09311_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13588_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net1937),
    .S1(net1923),
    .Z(_09312_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13589_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net1937),
    .S1(net1923),
    .Z(_09313_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13590_ (.I0(_09310_),
    .I1(_09311_),
    .I2(_09312_),
    .I3(_09313_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09314_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13591_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net1937),
    .S1(net1922),
    .Z(_09315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13592_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net1922),
    .Z(_09316_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13593_ (.A1(net1922),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .Z(_09317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13594_ (.I0(_09316_),
    .I1(_09317_),
    .S(net1854),
    .Z(_09318_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13595_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net1937),
    .S1(net1923),
    .Z(_09319_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13596_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S0(net2112),
    .S1(net1922),
    .Z(_09320_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13597_ (.I0(_09315_),
    .I1(_09318_),
    .I2(_09319_),
    .I3(_09320_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _13598_ (.I0(_09314_),
    .I1(_09321_),
    .S(net1860),
    .Z(_09322_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13599_ (.A1(_07905_),
    .A2(net2054),
    .B(net2057),
    .ZN(_09323_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13600_ (.I0(net1756),
    .I1(_09323_),
    .S(net1795),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13601_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09324_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13602_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S0(net2193),
    .S1(net1978),
    .Z(_09325_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13603_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13604_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net2193),
    .Z(_09327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13605_ (.A1(net2010),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .Z(_09328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13606_ (.I0(_09327_),
    .I1(_09328_),
    .S(net1868),
    .Z(_09329_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13607_ (.I0(_09324_),
    .I1(_09325_),
    .I2(_09326_),
    .I3(_09329_),
    .S0(net1878),
    .S1(net1866),
    .Z(_09330_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13608_ (.A1(net1958),
    .A2(_09330_),
    .ZN(_09331_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13609_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09332_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13610_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13611_ (.I0(_09332_),
    .I1(_09333_),
    .S(net1878),
    .Z(_09334_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13612_ (.A1(net1876),
    .A2(_09334_),
    .ZN(_09335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13613_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09336_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13614_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S0(net2010),
    .S1(net1978),
    .Z(_09337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13615_ (.I0(_09336_),
    .I1(_09337_),
    .S(net1878),
    .Z(_09338_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13616_ (.A1(net1832),
    .A2(_09338_),
    .ZN(_09339_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13617_ (.A1(_09331_),
    .A2(_09335_),
    .A3(_09339_),
    .Z(_09340_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _13618_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1756),
    .ZN(_09341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13619_ (.A1(net2028),
    .A2(_09340_),
    .B(_09341_),
    .ZN(_09342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13620_ (.I0(net2175),
    .I1(net2111),
    .S(_01334_),
    .Z(_09343_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13621_ (.A1(_08187_),
    .A2(_09342_),
    .B(_09343_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13622_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(net1801),
    .ZN(_09344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13623_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net1818),
    .ZN(_09345_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13624_ (.A1(net1742),
    .A2(_09340_),
    .B1(_09344_),
    .B2(net1741),
    .C(_09345_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13625_ (.I(net1676),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13626_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S0(net1943),
    .S1(net1926),
    .Z(_09346_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13627_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S0(net1943),
    .S1(net1926),
    .Z(_09347_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13628_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net2182),
    .S1(net1926),
    .Z(_09348_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13629_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net1943),
    .S1(net1926),
    .Z(_09349_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13630_ (.I0(_09346_),
    .I1(_09347_),
    .I2(_09348_),
    .I3(_09349_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09350_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13631_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net1943),
    .S1(net1925),
    .Z(_09351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13632_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net1925),
    .Z(_09352_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13633_ (.A1(net1925),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .Z(_09353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13634_ (.I0(_09352_),
    .I1(_09353_),
    .S(net1853),
    .Z(_09354_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13635_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net2182),
    .S1(net1926),
    .Z(_09355_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13636_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S0(net1943),
    .S1(net1925),
    .Z(_09356_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13637_ (.I0(_09351_),
    .I1(_09354_),
    .I2(_09355_),
    .I3(_09356_),
    .S0(net1851),
    .S1(net1900),
    .Z(_09357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13638_ (.I0(_09350_),
    .I1(_09357_),
    .S(net1860),
    .Z(_09358_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1542 (.I(_06893_),
    .Z(net1541));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13640_ (.A1(_07926_),
    .A2(net2054),
    .B(net2057),
    .ZN(_09360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13641_ (.I0(net1755),
    .I1(_09360_),
    .S(net1795),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13642_ (.I(_01341_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13643_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09361_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13644_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09362_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13645_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13646_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net2016),
    .Z(_09364_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13647_ (.A1(net2016),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .Z(_09365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13648_ (.I0(_09364_),
    .I1(_09365_),
    .S(net1875),
    .Z(_09366_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13649_ (.I0(_09361_),
    .I1(_09362_),
    .I2(_09363_),
    .I3(_09366_),
    .S0(net1878),
    .S1(net1866),
    .Z(_09367_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13650_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09368_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13651_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09369_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13652_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09370_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13653_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S0(net2016),
    .S1(net1981),
    .Z(_09371_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13654_ (.I0(_09368_),
    .I1(_09369_),
    .I2(_09370_),
    .I3(_09371_),
    .S0(net1878),
    .S1(net1866),
    .Z(_09372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13655_ (.A1(net1843),
    .A2(_09372_),
    .Z(_09373_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13656_ (.A1(net1958),
    .A2(_09367_),
    .B(_09373_),
    .ZN(_09374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13657_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(net1801),
    .ZN(_09375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13658_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net1818),
    .ZN(_09376_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13659_ (.A1(net1742),
    .A2(net1754),
    .B1(_09375_),
    .B2(net1741),
    .C(_09376_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13660_ (.I(net1675),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13661_ (.I(_00925_),
    .ZN(_09377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13662_ (.I(_00929_),
    .ZN(_09378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13663_ (.A1(_00929_),
    .A2(_00924_),
    .B(_00928_),
    .ZN(_09379_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13664_ (.A1(_09377_),
    .A2(_09378_),
    .A3(_09289_),
    .B(_09379_),
    .ZN(_09380_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_4 _13665_ (.A1(_00933_),
    .A2(_09380_),
    .Z(net175));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13666_ (.A1(_08919_),
    .A2(_08921_),
    .A3(_09107_),
    .ZN(_09381_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13667_ (.A1(_09115_),
    .A2(_09113_),
    .Z(_09382_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13668_ (.A1(net2123),
    .A2(_09381_),
    .B(_09382_),
    .ZN(_09383_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13669_ (.I(_09297_),
    .ZN(_09384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13670_ (.A1(_09197_),
    .A2(_09383_),
    .B(_09384_),
    .ZN(_09385_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13671_ (.A1(_09285_),
    .A2(_09377_),
    .A3(_00929_),
    .Z(_09386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13672_ (.A1(_00925_),
    .A2(_09287_),
    .Z(_09387_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13673_ (.A1(_00924_),
    .A2(_09387_),
    .Z(_09388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13674_ (.A1(_00925_),
    .A2(_00920_),
    .B(_00924_),
    .ZN(_09389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13675_ (.I0(_09388_),
    .I1(_09389_),
    .S(_09378_),
    .Z(_09390_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13676_ (.A1(_09378_),
    .A2(_00920_),
    .A3(_00924_),
    .ZN(_09391_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13677_ (.A1(_09302_),
    .A2(_09117_),
    .B(_09297_),
    .C(_09391_),
    .ZN(_09392_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13678_ (.A1(_09386_),
    .A2(_09385_),
    .B(_09390_),
    .C(_09392_),
    .ZN(net174));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13679_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_09393_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13680_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_09394_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13681_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_09395_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13682_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net1943),
    .S1(net1928),
    .Z(_09396_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13683_ (.I0(_09393_),
    .I1(_09394_),
    .I2(_09395_),
    .I3(_09396_),
    .S0(net1847),
    .S1(net1900),
    .Z(_09397_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13684_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net1943),
    .S1(net1929),
    .Z(_09398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13685_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net1929),
    .Z(_09399_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13686_ (.A1(net1929),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .Z(_09400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13687_ (.I0(_09399_),
    .I1(_09400_),
    .S(net1853),
    .Z(_09401_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13688_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net1942),
    .S1(net1929),
    .Z(_09402_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13689_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net1943),
    .S1(net1929),
    .Z(_09403_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13690_ (.I0(_09398_),
    .I1(_09401_),
    .I2(_09402_),
    .I3(_09403_),
    .S0(net1847),
    .S1(net1900),
    .Z(_09404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13691_ (.I0(_09397_),
    .I1(_09404_),
    .S(net1860),
    .Z(_09405_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1541 (.I(_00011_),
    .Z(net1540));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13693_ (.A1(net1845),
    .A2(net2054),
    .B(net2056),
    .ZN(_09407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13694_ (.I0(net1753),
    .I1(_09407_),
    .S(net1795),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13695_ (.I(_01348_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13696_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09408_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13697_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09409_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13698_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13699_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net2016),
    .Z(_09411_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13700_ (.A1(net2016),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .Z(_09412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13701_ (.I0(_09411_),
    .I1(_09412_),
    .S(net1875),
    .Z(_09413_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13702_ (.I0(_09408_),
    .I1(_09409_),
    .I2(_09410_),
    .I3(_09413_),
    .S0(net1877),
    .S1(net1866),
    .Z(_09414_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13703_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09415_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13704_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09416_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13705_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09417_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13706_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S0(net2016),
    .S1(net1987),
    .Z(_09418_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13707_ (.I0(_09415_),
    .I1(_09416_),
    .I2(_09417_),
    .I3(_09418_),
    .S0(net1877),
    .S1(net1866),
    .Z(_09419_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13708_ (.A1(net1842),
    .A2(_09419_),
    .Z(_09420_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13709_ (.A1(net1958),
    .A2(_09414_),
    .B(_09420_),
    .ZN(_09421_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13710_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(net1801),
    .ZN(_09422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13711_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net1818),
    .ZN(_09423_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13712_ (.A1(net1742),
    .A2(net1752),
    .B1(_09422_),
    .B2(net1741),
    .C(_09423_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13713_ (.I(_01347_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13714_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net2140),
    .S1(net1914),
    .Z(_09424_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13715_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net2139),
    .S1(net1914),
    .Z(_09425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13716_ (.I0(_09424_),
    .I1(_09425_),
    .S(net1847),
    .Z(_09426_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13717_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_09427_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13718_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .S0(net1914),
    .S1(net1904),
    .Z(_09428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13719_ (.I0(_09427_),
    .I1(_09428_),
    .S(net1857),
    .Z(_09429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13720_ (.I0(_09426_),
    .I1(_09429_),
    .S(net1859),
    .Z(_09430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13721_ (.A1(net1899),
    .A2(_09430_),
    .ZN(_09431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13722_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net1914),
    .Z(_09432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13723_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(net1828),
    .B1(_09432_),
    .B2(net1936),
    .C(net1904),
    .ZN(_09433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13724_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .S(net1914),
    .Z(_09434_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13725_ (.A1(net1936),
    .A2(net1848),
    .A3(_09434_),
    .ZN(_09435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13726_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S(net1914),
    .Z(_09436_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13727_ (.A1(_07840_),
    .A2(_09436_),
    .ZN(_09437_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13728_ (.A1(_07684_),
    .A2(_09433_),
    .A3(_09435_),
    .A4(_09437_),
    .Z(_09438_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13729_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S0(net1935),
    .S1(net1914),
    .Z(_09439_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13730_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S0(net1935),
    .S1(net1914),
    .Z(_09440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13731_ (.I0(_09439_),
    .I1(_09440_),
    .S(net1848),
    .Z(_09441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13732_ (.A1(_07846_),
    .A2(_09441_),
    .ZN(_09442_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13733_ (.A1(_09431_),
    .A2(_09438_),
    .A3(_09442_),
    .ZN(_09443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13734_ (.A1(_07706_),
    .A2(_07714_),
    .B(net2061),
    .ZN(_09444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13735_ (.A1(net1891),
    .A2(net1795),
    .ZN(_09445_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13736_ (.A1(_09444_),
    .A2(_09445_),
    .ZN(_09446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13737_ (.A1(net1797),
    .A2(net1719),
    .B(_09446_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13738_ (.I(_00943_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13739_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S0(net2006),
    .S1(net1975),
    .Z(_09447_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13740_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S0(net2006),
    .S1(net1975),
    .Z(_09448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13741_ (.I0(_09447_),
    .I1(_09448_),
    .S(net1881),
    .Z(_09449_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13742_ (.A1(net1832),
    .A2(_09449_),
    .ZN(_09450_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13743_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net2006),
    .S1(net1975),
    .Z(_09451_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13744_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net2006),
    .S1(net1975),
    .Z(_09452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13745_ (.I0(_09451_),
    .I1(_09452_),
    .S(net1881),
    .Z(_09453_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13746_ (.A1(_07523_),
    .A2(_09453_),
    .ZN(_09454_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13747_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S0(net2005),
    .S1(net1962),
    .Z(_09455_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13748_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net2008),
    .S1(net1962),
    .Z(_09456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13749_ (.I0(_09455_),
    .I1(_09456_),
    .S(net1866),
    .Z(_09457_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13750_ (.A1(net1958),
    .A2(net1868),
    .A3(_09457_),
    .ZN(_09458_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13751_ (.A1(net1975),
    .A2(_09455_),
    .Z(_09459_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _13752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .I2(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .I3(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .S0(net2007),
    .S1(net1962),
    .Z(_09460_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13753_ (.A1(net1958),
    .A2(net1866),
    .A3(_09459_),
    .A4(_09460_),
    .Z(_09461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13754_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .S(net2005),
    .Z(_09462_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13755_ (.A1(net2008),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .Z(_09463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13756_ (.I0(_09462_),
    .I1(_09463_),
    .S(net1877),
    .Z(_09464_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13757_ (.A1(net1958),
    .A2(net1959),
    .A3(net1975),
    .A4(_09464_),
    .Z(_09465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13758_ (.A1(_09461_),
    .A2(_09465_),
    .ZN(_09466_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13759_ (.A1(_09450_),
    .A2(_09454_),
    .A3(_09458_),
    .A4(_09466_),
    .Z(_09467_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13760_ (.A1(\cs_registers_i.pc_id_i[31] ),
    .A2(net1801),
    .Z(_09468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13761_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net1818),
    .B1(net2100),
    .B2(_09468_),
    .ZN(_09469_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13762_ (.A1(net2127),
    .A2(_09467_),
    .B(_09469_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13763_ (.I(_00938_),
    .ZN(_09470_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13765_ (.A1(_09431_),
    .A2(_09438_),
    .A3(_09442_),
    .Z(_09471_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13766_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .B2(net1824),
    .ZN(_09472_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13767_ (.A1(_08228_),
    .A2(_09471_),
    .B1(_09467_),
    .B2(net2028),
    .C(_09472_),
    .ZN(_09473_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13768_ (.A1(net2175),
    .A2(_00939_),
    .B(_09473_),
    .ZN(_09474_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13769_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net1823),
    .Z(_09475_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13770_ (.A1(_09474_),
    .A2(_09475_),
    .Z(_09476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13771_ (.I(_09379_),
    .ZN(_09477_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13772_ (.A1(_00933_),
    .A2(_09477_),
    .Z(_09478_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13773_ (.A1(_00932_),
    .A2(_09478_),
    .Z(_09479_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13774_ (.A1(_00937_),
    .A2(_09479_),
    .B(_00936_),
    .ZN(_09480_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13775_ (.A1(_00925_),
    .A2(_00929_),
    .A3(_00933_),
    .A4(_00937_),
    .ZN(_09481_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13776_ (.A1(_09289_),
    .A2(_09481_),
    .Z(_09482_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _13777_ (.A1(net2175),
    .A2(_00939_),
    .A3(_09470_),
    .ZN(_09483_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13778_ (.A1(net1815),
    .A2(_09483_),
    .ZN(_09484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _13779_ (.A1(net1815),
    .A2(_09476_),
    .B1(_09482_),
    .B2(_09480_),
    .C(_09484_),
    .ZN(_09485_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _13780_ (.A1(_09474_),
    .A2(_09475_),
    .ZN(_09486_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13781_ (.A1(_09481_),
    .A2(_09289_),
    .B(_09480_),
    .ZN(_09487_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13782_ (.A1(net1783),
    .A2(_09483_),
    .Z(_09488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13783_ (.A1(net1815),
    .A2(_09486_),
    .B(_09488_),
    .C(_09487_),
    .ZN(_09489_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _13784_ (.A1(_09485_),
    .A2(_09489_),
    .Z(net178));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13785_ (.A1(_00921_),
    .A2(_00925_),
    .A3(_00929_),
    .A4(_00933_),
    .ZN(_09490_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13786_ (.A1(_09285_),
    .A2(_09297_),
    .B(_09286_),
    .ZN(_09491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13787_ (.A1(_00925_),
    .A2(_09491_),
    .B(_00924_),
    .ZN(_09492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13788_ (.I(_00928_),
    .ZN(_09493_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13789_ (.A1(_09378_),
    .A2(_09492_),
    .B(_09493_),
    .ZN(_09494_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13790_ (.A1(_00933_),
    .A2(_09494_),
    .B(_00932_),
    .ZN(_09495_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13791_ (.A1(_09302_),
    .A2(_09117_),
    .A3(_09490_),
    .B(_09495_),
    .ZN(_09496_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _13792_ (.A1(_09496_),
    .A2(_00937_),
    .Z(net177));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13793_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_09497_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13794_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .ZN(_09498_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13795_ (.A1(_09497_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A3(_09498_),
    .A4(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_09499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13796_ (.I(_09499_),
    .ZN(_09500_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13797_ (.A1(_08143_),
    .A2(_08145_),
    .Z(_09501_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13798_ (.A1(_08156_),
    .A2(_08164_),
    .A3(_08168_),
    .A4(_09501_),
    .Z(_09502_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13799_ (.A1(_08121_),
    .A2(_08209_),
    .A3(_08123_),
    .Z(_09503_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13800_ (.A1(net2147),
    .A2(\id_stage_i.controller_i.instr_i[13] ),
    .A3(_07579_),
    .Z(_09504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13801_ (.A1(_07566_),
    .A2(\id_stage_i.controller_i.instr_i[14] ),
    .Z(_09505_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13802_ (.A1(_09504_),
    .A2(_09505_),
    .B(\id_stage_i.controller_i.instr_i[5] ),
    .ZN(_09506_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13803_ (.A1(net2147),
    .A2(_08000_),
    .A3(_08150_),
    .Z(_09507_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13804_ (.A1(_07586_),
    .A2(_07615_),
    .ZN(_09508_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13805_ (.A1(_09506_),
    .A2(_09507_),
    .B(net1889),
    .C(_09508_),
    .ZN(_09509_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13806_ (.A1(_07568_),
    .A2(_08122_),
    .B(net2132),
    .ZN(_09510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _13807_ (.A1(_07560_),
    .A2(_07590_),
    .B1(_08047_),
    .B2(_07588_),
    .ZN(_09511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13808_ (.A1(_07559_),
    .A2(net1831),
    .ZN(_09512_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13809_ (.A1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .A2(_07582_),
    .ZN(_09513_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13810_ (.A1(_07565_),
    .A2(_09510_),
    .B1(_09511_),
    .B2(_09512_),
    .C(_09513_),
    .ZN(_09514_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _13811_ (.A1(_09502_),
    .A2(_09503_),
    .A3(_09509_),
    .A4(_09514_),
    .ZN(_09515_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13812_ (.A1(_08158_),
    .A2(net1826),
    .Z(_09516_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13813_ (.A1(\id_stage_i.controller_i.instr_i[14] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .Z(_09517_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13814_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Z(_09518_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13815_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .ZN(_09519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13816_ (.A1(_07968_),
    .A2(_09519_),
    .ZN(_09520_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13817_ (.A1(_08004_),
    .A2(_09517_),
    .A3(_09518_),
    .A4(_09520_),
    .Z(_09521_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13818_ (.A1(_09516_),
    .A2(_09521_),
    .Z(_09522_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13819_ (.A1(net1908),
    .A2(net1903),
    .A3(net1892),
    .ZN(_09523_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13820_ (.A1(net1827),
    .A2(_08167_),
    .A3(_09523_),
    .ZN(_09524_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13821_ (.A1(net1899),
    .A2(net1898),
    .A3(net1891),
    .Z(_09525_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13822_ (.A1(net1908),
    .A2(_08180_),
    .A3(_09525_),
    .Z(_09526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13823_ (.A1(net1858),
    .A2(net1895),
    .ZN(_09527_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13824_ (.A1(net1894),
    .A2(_07840_),
    .A3(_09526_),
    .A4(_09527_),
    .Z(_09528_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13825_ (.A1(_07860_),
    .A2(_08546_),
    .ZN(_09529_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13826_ (.A1(net1899),
    .A2(net1898),
    .A3(net1896),
    .A4(net1892),
    .Z(_09530_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _13827_ (.A1(net1899),
    .A2(net1898),
    .A3(net1896),
    .A4(net1892),
    .ZN(_09531_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13828_ (.A1(_09530_),
    .A2(_09531_),
    .ZN(_09532_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13829_ (.A1(net1900),
    .A2(_07926_),
    .A3(_07905_),
    .Z(_09533_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13830_ (.A1(net1855),
    .A2(net1908),
    .A3(net1848),
    .ZN(_09534_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13831_ (.A1(_09529_),
    .A2(_09532_),
    .A3(_09533_),
    .A4(_09534_),
    .Z(_09535_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13832_ (.A1(_09516_),
    .A2(_09524_),
    .A3(_09528_),
    .A4(_09535_),
    .Z(_09536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13833_ (.A1(_09522_),
    .A2(_09536_),
    .ZN(_09537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13834_ (.A1(_09515_),
    .A2(_09537_),
    .Z(_09538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13835_ (.I(_09538_),
    .ZN(_09539_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13836_ (.A1(_08043_),
    .A2(_09539_),
    .B(\id_stage_i.controller_i.instr_valid_i ),
    .ZN(_09540_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13837_ (.A1(_08043_),
    .A2(_09515_),
    .A3(_09537_),
    .Z(_09541_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13839_ (.A1(net1699),
    .A2(net1698),
    .A3(net1697),
    .A4(_09541_),
    .Z(_09543_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13840_ (.A1(_07708_),
    .A2(_07716_),
    .A3(_07741_),
    .A4(net1701),
    .Z(_09544_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13841_ (.A1(net2068),
    .A2(net1610),
    .ZN(_09545_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13842_ (.A1(_07859_),
    .A2(_01180_),
    .A3(_09541_),
    .Z(_09546_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13843_ (.A1(_09543_),
    .A2(_09544_),
    .A3(_09545_),
    .A4(_09546_),
    .Z(_09547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13844_ (.A1(net1896),
    .A2(_07860_),
    .ZN(_09548_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13845_ (.A1(_07893_),
    .A2(_07897_),
    .A3(_07903_),
    .ZN(_09549_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13846_ (.A1(net1795),
    .A2(net1790),
    .A3(_09549_),
    .Z(_09550_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13847_ (.A1(net1797),
    .A2(_07861_),
    .A3(_09548_),
    .B(_09550_),
    .ZN(_09551_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13848_ (.A1(net1700),
    .A2(_09551_),
    .Z(_09552_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13849_ (.A1(net1699),
    .A2(net1698),
    .A3(_01212_),
    .Z(_09553_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13850_ (.A1(net1701),
    .A2(net1696),
    .A3(_09541_),
    .Z(_09554_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13851_ (.A1(_09541_),
    .A2(_09552_),
    .A3(_09553_),
    .A4(_09554_),
    .Z(_09555_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13852_ (.A1(_07710_),
    .A2(_07768_),
    .A3(_07769_),
    .ZN(_09556_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13853_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(net2061),
    .A3(net2067),
    .Z(_09557_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13854_ (.A1(_09556_),
    .A2(_09557_),
    .A3(_01159_),
    .B(_09541_),
    .ZN(_09558_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13855_ (.A1(_09547_),
    .A2(_09555_),
    .B(_09558_),
    .ZN(_09559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13856_ (.A1(\id_stage_i.controller_i.instr_is_compressed_i ),
    .A2(_07697_),
    .A3(_07699_),
    .ZN(_09560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13857_ (.A1(net1908),
    .A2(_07706_),
    .ZN(_09561_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13858_ (.A1(_09560_),
    .A2(_09561_),
    .B(_07775_),
    .ZN(_09562_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _13859_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A2(net2061),
    .A3(_07710_),
    .A4(net2067),
    .Z(_09563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13860_ (.I0(net1855),
    .I1(_07968_),
    .S(net2069),
    .Z(_09564_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13861_ (.A1(net2061),
    .A2(_07655_),
    .ZN(_09565_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13862_ (.A1(net1798),
    .A2(net2185),
    .B(net1797),
    .ZN(_09566_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13863_ (.A1(_09564_),
    .A2(_09565_),
    .B(_09566_),
    .ZN(_09567_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13864_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09567_),
    .ZN(_09568_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13865_ (.A1(net1612),
    .A2(_07708_),
    .A3(_07716_),
    .A4(_07741_),
    .Z(_09569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13866_ (.I0(_09568_),
    .I1(_09569_),
    .S(_07859_),
    .Z(_09570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13867_ (.A1(net1699),
    .A2(_09541_),
    .Z(_09571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13868_ (.I(_08162_),
    .ZN(_09572_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13869_ (.A1(net1797),
    .A2(_07861_),
    .A3(_09572_),
    .Z(_09573_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13870_ (.A1(net1790),
    .A2(net1788),
    .B(net1797),
    .ZN(_09574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13871_ (.A1(_09573_),
    .A2(_09574_),
    .Z(_09575_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13872_ (.A1(net1698),
    .A2(_01212_),
    .Z(_09576_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13873_ (.A1(net1696),
    .A2(_09571_),
    .A3(_09575_),
    .A4(_09576_),
    .Z(_09577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13874_ (.A1(net1702),
    .A2(_09541_),
    .Z(_09578_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13875_ (.A1(_07773_),
    .A2(_09578_),
    .Z(_09579_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13876_ (.A1(net1701),
    .A2(_09570_),
    .A3(_09577_),
    .A4(_09579_),
    .ZN(_09580_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13877_ (.A1(net1611),
    .A2(_09568_),
    .A3(_09578_),
    .Z(_09581_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13878_ (.A1(net2068),
    .A2(_09553_),
    .A3(_09546_),
    .A4(_09554_),
    .Z(_09582_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13879_ (.A1(_09558_),
    .A2(_09581_),
    .B(_09582_),
    .ZN(_09583_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13880_ (.A1(_09559_),
    .A2(_09580_),
    .A3(_09583_),
    .Z(_09584_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13881_ (.A1(net1831),
    .A2(net1826),
    .ZN(_09585_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13882_ (.A1(_09502_),
    .A2(_09503_),
    .A3(_09509_),
    .A4(_09514_),
    .Z(_09586_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13883_ (.A1(_09522_),
    .A2(_09536_),
    .Z(_09587_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13884_ (.A1(_09585_),
    .A2(_09586_),
    .A3(_09587_),
    .Z(_09588_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13885_ (.A1(net1797),
    .A2(net2185),
    .Z(_09589_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13886_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09589_),
    .B(net1612),
    .ZN(_09590_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13887_ (.A1(net1702),
    .A2(net1701),
    .Z(_09591_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13888_ (.A1(_07773_),
    .A2(_09590_),
    .A3(_09591_),
    .Z(_09592_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13889_ (.A1(net1702),
    .A2(net1701),
    .A3(_07859_),
    .Z(_09593_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13890_ (.A1(_09588_),
    .A2(_09593_),
    .ZN(_09594_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13891_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09567_),
    .B(_09541_),
    .ZN(_09595_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13892_ (.A1(net1611),
    .A2(_09569_),
    .B(net1608),
    .ZN(_09596_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _13893_ (.A1(_07859_),
    .A2(_09588_),
    .A3(_09592_),
    .B1(_09594_),
    .B2(_09596_),
    .ZN(_09597_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _13894_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09567_),
    .Z(_09598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13895_ (.A1(net1702),
    .A2(_09541_),
    .ZN(_09599_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13896_ (.A1(_07773_),
    .A2(_09598_),
    .A3(_09599_),
    .Z(_09600_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13897_ (.A1(net1701),
    .A2(_09588_),
    .ZN(_09601_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _13898_ (.A1(net1797),
    .A2(_07861_),
    .A3(_09572_),
    .B(_09574_),
    .ZN(_09602_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13899_ (.A1(net1700),
    .A2(_09602_),
    .ZN(_09603_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13900_ (.A1(net1610),
    .A2(_09601_),
    .A3(_09603_),
    .ZN(_09604_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13901_ (.A1(net1698),
    .A2(net1697),
    .A3(_09571_),
    .ZN(_09605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13902_ (.A1(_07770_),
    .A2(_07771_),
    .Z(_09606_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _13903_ (.A1(_09606_),
    .A2(net1702),
    .B(_01212_),
    .C(_09588_),
    .ZN(_09607_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13904_ (.A1(net1698),
    .A2(_09571_),
    .ZN(_09608_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13905_ (.A1(net1696),
    .A2(_09552_),
    .A3(_09601_),
    .ZN(_09609_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_4 _13906_ (.A1(_09600_),
    .A2(_09604_),
    .A3(_09605_),
    .B1(_09607_),
    .B2(_09608_),
    .B3(_09609_),
    .ZN(_09610_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13907_ (.A1(net1797),
    .A2(_07861_),
    .A3(_09548_),
    .Z(_09611_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13908_ (.A1(_09550_),
    .A2(_09611_),
    .Z(_09612_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13909_ (.A1(_07773_),
    .A2(_09598_),
    .A3(_09544_),
    .A4(_09578_),
    .Z(_09613_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _13910_ (.A1(_07859_),
    .A2(net1610),
    .A3(_09541_),
    .A4(_09553_),
    .ZN(_09614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13911_ (.A1(_09612_),
    .A2(_09602_),
    .B(_09613_),
    .C(_09614_),
    .ZN(_09615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13912_ (.A1(_09577_),
    .A2(_09597_),
    .B(_09610_),
    .C(_09615_),
    .ZN(_09616_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13913_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .ZN(_09617_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13914_ (.A1(_09498_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_09618_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13915_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09617_),
    .A3(_09618_),
    .Z(_09619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13916_ (.A1(_07642_),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .ZN(_09620_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13917_ (.A1(_09619_),
    .A2(_09620_),
    .ZN(_09621_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13918_ (.A1(_00952_),
    .A2(_09621_),
    .Z(_09622_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _13919_ (.A1(_01212_),
    .A2(net1696),
    .A3(_09585_),
    .A4(_09622_),
    .Z(_09623_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13920_ (.A1(_09538_),
    .A2(_09623_),
    .ZN(_09624_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13921_ (.A1(_09585_),
    .A2(_09586_),
    .A3(_09587_),
    .Z(_09625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13922_ (.A1(_07773_),
    .A2(net1702),
    .B(_09625_),
    .ZN(_09626_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13923_ (.A1(_08043_),
    .A2(_09515_),
    .A3(_09537_),
    .Z(_09627_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _13924_ (.A1(net1699),
    .A2(net1698),
    .A3(net1697),
    .A4(_09627_),
    .Z(_09628_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13925_ (.A1(net1700),
    .A2(_09627_),
    .A3(_09551_),
    .Z(_09629_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13926_ (.A1(net1701),
    .A2(net1610),
    .ZN(_09630_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13927_ (.A1(_09628_),
    .A2(_09629_),
    .A3(_09630_),
    .ZN(_09631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13928_ (.I(_00958_),
    .ZN(_09632_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13929_ (.A1(_00956_),
    .A2(_09632_),
    .B(_00955_),
    .ZN(_09633_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13930_ (.A1(_00956_),
    .A2(_00959_),
    .Z(_09634_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13931_ (.A1(_09633_),
    .A2(_09634_),
    .Z(_09635_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _13932_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09626_),
    .A3(_09631_),
    .B(_09635_),
    .ZN(_09636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13933_ (.A1(_09584_),
    .A2(_09616_),
    .B(_09624_),
    .C(_09636_),
    .ZN(_09637_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _13934_ (.A1(_07860_),
    .A2(_08546_),
    .A3(_09530_),
    .ZN(_09638_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13935_ (.A1(_09533_),
    .A2(_09534_),
    .A3(_09638_),
    .Z(_09639_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13936_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(\cs_registers_i.priv_mode_id_o[0] ),
    .Z(_09640_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13937_ (.I(_09528_),
    .ZN(_09641_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _13938_ (.A1(_08180_),
    .A2(_09525_),
    .A3(_09533_),
    .A4(_09534_),
    .ZN(_09642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13939_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_09641_),
    .B(_09642_),
    .ZN(_09643_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _13940_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09639_),
    .B1(_09640_),
    .B2(_09643_),
    .ZN(_09644_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13941_ (.A1(_07595_),
    .A2(_07574_),
    .Z(_09645_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13942_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_09645_),
    .A3(net1826),
    .Z(_09646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13943_ (.A1(_09644_),
    .A2(_09646_),
    .ZN(_09647_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13944_ (.A1(_09540_),
    .A2(_09637_),
    .B(_09647_),
    .ZN(_09648_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13945_ (.A1(_09500_),
    .A2(_09648_),
    .Z(\id_stage_i.controller_i.illegal_insn_d ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13946_ (.A1(net1827),
    .A2(_08167_),
    .A3(_09523_),
    .Z(_09649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13947_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Z(_09650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _13948_ (.A1(_09649_),
    .A2(_09646_),
    .B(net1840),
    .ZN(_09651_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _13949_ (.A1(_09540_),
    .A2(_09637_),
    .B(_09647_),
    .C(_09651_),
    .ZN(_09652_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13950_ (.A1(_09500_),
    .A2(_09652_),
    .Z(\id_stage_i.controller_i.exc_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13951_ (.A1(_07553_),
    .A2(_07550_),
    .Z(_09653_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13952_ (.A1(net64),
    .A2(_09653_),
    .ZN(_09654_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13953_ (.I(net30),
    .ZN(_09655_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13954_ (.I(\load_store_unit_i.lsu_err_q ),
    .ZN(_09656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13955_ (.A1(_09655_),
    .A2(_09656_),
    .Z(_09657_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13956_ (.A1(_09654_),
    .A2(_09657_),
    .ZN(_09658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13957_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_09658_),
    .Z(\id_stage_i.controller_i.store_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _13958_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_09654_),
    .A3(_09657_),
    .ZN(\id_stage_i.controller_i.load_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13960_ (.A1(net1831),
    .A2(_08182_),
    .Z(_09660_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13962_ (.I(net1751),
    .ZN(_09662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13963_ (.A1(net2032),
    .A2(_09662_),
    .Z(_09663_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13964_ (.A1(net2030),
    .A2(_09663_),
    .Z(_09664_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13965_ (.A1(_07579_),
    .A2(net1897),
    .A3(net1783),
    .Z(_09665_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13968_ (.A1(net2019),
    .A2(_07860_),
    .A3(net1815),
    .Z(_09668_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _13970_ (.A1(net2031),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(net1823),
    .Z(_09670_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _13971_ (.A1(_09450_),
    .A2(_09454_),
    .A3(_09458_),
    .A4(_09466_),
    .ZN(_09671_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13972_ (.A1(net2021),
    .A2(_08047_),
    .ZN(_09672_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13973_ (.A1(_07596_),
    .A2(_08182_),
    .A3(_09672_),
    .Z(_09673_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13974_ (.A1(net1717),
    .A2(_09673_),
    .ZN(_09674_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13975_ (.A1(_07579_),
    .A2(net1825),
    .ZN(_09675_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13976_ (.A1(net2020),
    .A2(_07860_),
    .B(_09675_),
    .ZN(_09676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _13977_ (.A1(net2020),
    .A2(net1825),
    .B1(_09676_),
    .B2(net2022),
    .C(_08108_),
    .ZN(_09677_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13978_ (.A1(net2019),
    .A2(net1825),
    .A3(_09677_),
    .Z(_09678_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _13980_ (.A1(net1674),
    .A2(net1673),
    .ZN(_09680_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13981_ (.A1(net2022),
    .A2(_07579_),
    .B(_07640_),
    .ZN(_09681_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13982_ (.A1(_08182_),
    .A2(_09681_),
    .A3(_09443_),
    .Z(_09682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13983_ (.I0(net1674),
    .I1(_09680_),
    .S(net1672),
    .Z(_09683_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _13984_ (.A1(net1674),
    .A2(net1673),
    .B1(_09683_),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .C(net2031),
    .ZN(_09684_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _13985_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_09670_),
    .B(_09684_),
    .ZN(_09685_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _13986_ (.A1(_09539_),
    .A2(_09621_),
    .Z(_09686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _13987_ (.A1(net1750),
    .A2(_09685_),
    .B(_08187_),
    .C(_09686_),
    .ZN(_09687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13988_ (.A1(net1718),
    .A2(net1549),
    .Z(_09688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13989_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .I1(_09664_),
    .S(_09688_),
    .Z(_00000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _13990_ (.A1(net2032),
    .A2(net1751),
    .Z(_09689_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _13992_ (.I0(net2030),
    .I1(net1716),
    .S(_09688_),
    .Z(_00001_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1540 (.I(\alu_adder_result_ex[1] ),
    .Z(net1539));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _13997_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .ZN(_09695_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _13998_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .ZN(_09696_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _13999_ (.A1(_09695_),
    .A2(_00968_),
    .A3(_09696_),
    .Z(_09697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14000_ (.A1(net2027),
    .A2(_09697_),
    .Z(_09698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14001_ (.I(_09686_),
    .ZN(_09699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14002_ (.A1(_09699_),
    .A2(net1750),
    .Z(_09700_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14004_ (.I0(net2029),
    .I1(_09698_),
    .S(_09700_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14005_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A2(_09700_),
    .Z(_09702_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14007_ (.A1(_09700_),
    .A2(_09697_),
    .B(_08194_),
    .ZN(_09704_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14008_ (.A1(net1548),
    .A2(_09704_),
    .Z(_00005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14009_ (.A1(net2111),
    .A2(_08395_),
    .B(_08401_),
    .ZN(_09705_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14010_ (.A1(net2109),
    .A2(_09705_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14011_ (.I(_01366_),
    .ZN(_09706_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14012_ (.A1(net2080),
    .A2(_08387_),
    .ZN(_09707_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14013_ (.A1(_09707_),
    .A2(net2300),
    .ZN(_09708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14014_ (.A1(_00833_),
    .A2(_09708_),
    .B(_00832_),
    .ZN(_09709_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14015_ (.A1(_00837_),
    .A2(_09709_),
    .ZN(net181));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14016_ (.A1(net2109),
    .A2(net2080),
    .B(_00824_),
    .ZN(_09710_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14017_ (.A1(_00829_),
    .A2(_09710_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14018_ (.A1(_09706_),
    .A2(net183),
    .A3(net181),
    .A4(net179),
    .Z(_09711_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14019_ (.A1(net185),
    .A2(net157),
    .A3(net163),
    .A4(_09711_),
    .Z(_09712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14020_ (.A1(_08460_),
    .A2(_08467_),
    .ZN(_09713_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14021_ (.A1(_08129_),
    .A2(_08170_),
    .B(_08460_),
    .C(_08184_),
    .ZN(_09714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14022_ (.A1(_09713_),
    .A2(_09714_),
    .ZN(_09715_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _14023_ (.A1(net2290),
    .A2(_09715_),
    .ZN(net180));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14024_ (.A1(net182),
    .A2(net165),
    .A3(net180),
    .Z(_09716_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14025_ (.A1(net156),
    .A2(net160),
    .A3(net164),
    .Z(_09717_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14026_ (.A1(net176),
    .A2(_09712_),
    .A3(_09716_),
    .A4(_09717_),
    .Z(_09718_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14027_ (.A1(net167),
    .A2(net168),
    .A3(net171),
    .A4(net172),
    .Z(_09719_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14028_ (.A1(net184),
    .A2(net159),
    .A3(net158),
    .A4(net161),
    .Z(_09720_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14029_ (.A1(net162),
    .A2(net166),
    .A3(net177),
    .A4(_09720_),
    .Z(_09721_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _14030_ (.A1(net169),
    .A2(_09718_),
    .A3(_09719_),
    .A4(_09721_),
    .ZN(_09722_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14031_ (.A1(_00925_),
    .A2(_09480_),
    .ZN(_09723_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14032_ (.A1(_09289_),
    .A2(_09723_),
    .Z(_09724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14033_ (.A1(net1783),
    .A2(_09483_),
    .ZN(_09725_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14034_ (.A1(net1783),
    .A2(_09476_),
    .B(_09724_),
    .C(_09725_),
    .ZN(_09726_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14035_ (.A1(net1815),
    .A2(_09483_),
    .Z(_09727_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14036_ (.A1(_09377_),
    .A2(_09289_),
    .A3(_09480_),
    .Z(_09728_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14037_ (.A1(net1783),
    .A2(_09486_),
    .B(_09727_),
    .C(_09728_),
    .ZN(_09729_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14038_ (.A1(_09726_),
    .A2(_09729_),
    .Z(_09730_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14039_ (.A1(_09480_),
    .A2(_09481_),
    .ZN(_09731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14040_ (.A1(_00925_),
    .A2(_09731_),
    .ZN(_09732_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14041_ (.A1(_09289_),
    .A2(_09732_),
    .Z(_09733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14042_ (.A1(net1815),
    .A2(_09486_),
    .B(_09733_),
    .C(_09488_),
    .ZN(_09734_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14043_ (.A1(_09377_),
    .A2(_09289_),
    .A3(_09731_),
    .Z(_09735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14044_ (.A1(net1815),
    .A2(_09476_),
    .B(_09484_),
    .C(_09735_),
    .ZN(_09736_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14045_ (.A1(_09734_),
    .A2(_09736_),
    .ZN(_09737_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14046_ (.A1(net2065),
    .A2(net2169),
    .A3(net174),
    .Z(_09738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14047_ (.A1(_09730_),
    .A2(_09737_),
    .B(_09738_),
    .ZN(_09739_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14048_ (.A1(_09722_),
    .A2(_09739_),
    .Z(_09740_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14049_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_09700_),
    .ZN(_09741_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14050_ (.A1(_08227_),
    .A2(_09700_),
    .B1(_09740_),
    .B2(_09741_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14051_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_09740_),
    .ZN(_09742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14052_ (.A1(_08192_),
    .A2(_09742_),
    .ZN(_09743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14053_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .I1(_09743_),
    .S(_09700_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14054_ (.I(\cs_registers_i.pc_if_i[2] ),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14055_ (.I(net1540),
    .ZN(\alu_adder_result_ex[0] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14056_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .S(net1751),
    .Z(_09744_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14057_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .Z(_09745_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_24_clk (.I(clknet_2_3_0_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14060_ (.A1(net2032),
    .A2(_09744_),
    .B1(net1839),
    .B2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .ZN(_09748_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14061_ (.I(_09748_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14062_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .ZN(_09749_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14063_ (.A1(_08755_),
    .A2(_09745_),
    .Z(_09750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14064_ (.A1(_07691_),
    .A2(net1838),
    .B(_09750_),
    .ZN(_09751_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_25_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14066_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(_09753_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_26_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14068_ (.I0(_08191_),
    .I1(_08775_),
    .S(net1836),
    .Z(_09755_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14069_ (.A1(net1671),
    .A2(_09755_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_27_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1539 (.I(_11434_),
    .Z(net1538));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14072_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .S(net1751),
    .Z(_09758_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1538 (.I(_00584_),
    .Z(net1537));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14074_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(net1839),
    .B1(_09758_),
    .B2(net2032),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14075_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .S(net1751),
    .Z(_09760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14076_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(net1839),
    .B1(_09760_),
    .B2(net2032),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_28_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_29_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14079_ (.A1(net1739),
    .A2(_09749_),
    .Z(_09763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14080_ (.A1(_08852_),
    .A2(_09745_),
    .B(_09763_),
    .ZN(_09764_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14081_ (.A1(_09755_),
    .A2(net1606),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14082_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .S(net1751),
    .Z(_09765_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14083_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(net1839),
    .B1(_09765_),
    .B2(net2032),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14084_ (.I0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .S(net1751),
    .Z(_09766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14085_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(net1839),
    .B1(_09766_),
    .B2(net2032),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_30_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14087_ (.I0(net2272),
    .I1(_08870_),
    .S(_09753_),
    .Z(_09768_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_31_clk (.I(clknet_2_2_0_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14089_ (.A1(net1606),
    .A2(net1666),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _14090_ (.A1(_07787_),
    .A2(_07793_),
    .A3(_07799_),
    .A4(_07803_),
    .ZN(_09770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14091_ (.A1(_08889_),
    .A2(_09745_),
    .Z(_09771_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14092_ (.A1(_09770_),
    .A2(_09749_),
    .B(_09771_),
    .ZN(_09772_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_32_clk (.I(clknet_2_1_0_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14094_ (.I0(net1785),
    .I1(_08810_),
    .S(_09753_),
    .Z(_09774_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_33_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14096_ (.A1(net1664),
    .A2(net1660),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14097_ (.I0(net1793),
    .I1(_08945_),
    .S(_09745_),
    .Z(_09776_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14098_ (.A1(_09755_),
    .A2(net1659),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14099_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .S(net1751),
    .Z(_09777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14100_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(net1839),
    .B1(_09777_),
    .B2(net2032),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14101_ (.I0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .S(net1751),
    .Z(_09778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14102_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(net1839),
    .B1(_09778_),
    .B2(net2032),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14103_ (.I(_09764_),
    .ZN(_09779_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _14104_ (.A1(_08298_),
    .A2(_08307_),
    .A3(_08314_),
    .ZN(_09780_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14105_ (.A1(net1958),
    .A2(_08949_),
    .A3(_08954_),
    .Z(_09781_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14106_ (.A1(_08961_),
    .A2(_09781_),
    .Z(_09782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14107_ (.I0(net1714),
    .I1(_09782_),
    .S(net1836),
    .Z(_09783_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14108_ (.A1(_09779_),
    .A2(net1603),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14109_ (.I0(net1779),
    .I1(_08906_),
    .S(_09753_),
    .Z(_09784_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_35_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14111_ (.A1(net1663),
    .A2(_09784_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14112_ (.A1(net1666),
    .A2(_09776_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14113_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .S(net1751),
    .Z(_09786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14114_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(net1839),
    .B1(_09786_),
    .B2(net2032),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14115_ (.I0(_08339_),
    .I1(_08999_),
    .S(_09753_),
    .Z(_09787_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_34_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14117_ (.A1(net1607),
    .A2(_09787_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14118_ (.I(_09772_),
    .ZN(_09789_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14119_ (.A1(_09789_),
    .A2(net1603),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_36_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14121_ (.A1(_09776_),
    .A2(_09784_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14122_ (.A1(net1791),
    .A2(net1838),
    .Z(_09791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14123_ (.A1(_08981_),
    .A2(_09745_),
    .B(_09791_),
    .ZN(_09792_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14124_ (.A1(net1666),
    .A2(_09792_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14125_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .S(net1751),
    .Z(_09793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14126_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(net1839),
    .B1(_09793_),
    .B2(net2032),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14127_ (.I0(_08361_),
    .I1(_09059_),
    .S(_09753_),
    .Z(_09794_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_37_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14129_ (.A1(net1607),
    .A2(net1649),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14130_ (.A1(net1663),
    .A2(_09787_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14131_ (.I(_09776_),
    .ZN(_09796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14132_ (.A1(_09796_),
    .A2(net1604),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14133_ (.A1(_09784_),
    .A2(_09792_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14134_ (.I0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .S(net1751),
    .Z(_09797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14135_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net1839),
    .B1(_09797_),
    .B2(net2032),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14136_ (.I0(_08378_),
    .I1(net1724),
    .S(net1837),
    .Z(_09798_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_38_clk (.I(clknet_2_0_0_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14138_ (.A1(net1606),
    .A2(_09798_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14139_ (.A1(net1662),
    .A2(net1651),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14140_ (.A1(_09776_),
    .A2(net1656),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14142_ (.I(net1653),
    .ZN(_09801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14143_ (.A1(net1603),
    .A2(_09801_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14144_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .S(net1751),
    .Z(_09802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14145_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net1839),
    .B1(_09802_),
    .B2(net2032),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14146_ (.I0(_08427_),
    .I1(_09148_),
    .S(net1837),
    .Z(_09803_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14148_ (.A1(net1607),
    .A2(_09803_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14149_ (.A1(net1662),
    .A2(_09798_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14150_ (.A1(_09776_),
    .A2(net1651),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14151_ (.A1(_09787_),
    .A2(net1653),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14152_ (.A1(_07914_),
    .A2(_07918_),
    .A3(_07923_),
    .Z(_09805_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14153_ (.A1(_09131_),
    .A2(_09745_),
    .Z(_09806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14154_ (.A1(_09805_),
    .A2(_09749_),
    .B(_09806_),
    .ZN(_09807_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_1_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14156_ (.A1(net1666),
    .A2(net1644),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14157_ (.I0(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .S(net1751),
    .Z(_09809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14158_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net1839),
    .B1(_09809_),
    .B2(net2032),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14159_ (.I0(net2167),
    .I1(_09182_),
    .S(net1837),
    .Z(_09810_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14161_ (.A1(net1607),
    .A2(net1642),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14162_ (.A1(net1662),
    .A2(_09803_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14163_ (.A1(_09776_),
    .A2(_09798_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_2_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_2_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14165_ (.A1(net1653),
    .A2(net1651),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14166_ (.A1(_09784_),
    .A2(_09807_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14167_ (.A1(_09258_),
    .A2(_09745_),
    .Z(_09813_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14168_ (.A1(net2075),
    .A2(net1838),
    .B(_09813_),
    .ZN(_09814_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload31 (.I(clknet_2_0_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14170_ (.A1(net1668),
    .A2(_09814_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14171_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .S(net1751),
    .Z(_09816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14172_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net1839),
    .B1(_09816_),
    .B2(net2032),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14173_ (.I0(_08486_),
    .I1(_09239_),
    .S(net1837),
    .Z(_09817_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1537 (.I(_00585_),
    .Z(net1536));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14175_ (.A1(net1607),
    .A2(_09817_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14176_ (.A1(net1663),
    .A2(net1642),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14177_ (.A1(_09776_),
    .A2(_09803_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14178_ (.A1(net1653),
    .A2(_09798_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14179_ (.I(_09807_),
    .ZN(_09819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14180_ (.A1(net1603),
    .A2(_09819_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14181_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .S(net1751),
    .Z(_09820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14182_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net1839),
    .B1(_09820_),
    .B2(net2032),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14183_ (.I0(net1738),
    .I1(_09276_),
    .S(net1837),
    .Z(_09821_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1536 (.I(_10228_),
    .Z(net1535));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14185_ (.A1(net1607),
    .A2(_09821_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14186_ (.A1(net1665),
    .A2(_09817_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14187_ (.A1(_09776_),
    .A2(net1642),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14188_ (.A1(net1653),
    .A2(net1646),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14189_ (.A1(_09787_),
    .A2(_09807_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14190_ (.A1(net1666),
    .A2(_09814_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14191_ (.A1(_09322_),
    .A2(_09745_),
    .Z(_09823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14192_ (.A1(net2105),
    .A2(net1838),
    .B(_09823_),
    .ZN(_09824_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1535 (.I(_01360_),
    .Z(net1534));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14194_ (.A1(net1661),
    .A2(net1598),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14195_ (.A1(_08586_),
    .A2(net1838),
    .Z(_09826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14196_ (.A1(_09358_),
    .A2(_09745_),
    .B(_09826_),
    .ZN(_09827_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1534 (.I(_01362_),
    .Z(net1533));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14198_ (.A1(net1668),
    .A2(_09827_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14199_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .S(net1751),
    .Z(_09829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14200_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net1839),
    .B1(_09829_),
    .B2(net2032),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14201_ (.I(net1802),
    .ZN(_09830_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _14202_ (.A1(_09331_),
    .A2(_09335_),
    .A3(_09339_),
    .ZN(_09831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14203_ (.I0(_09830_),
    .I1(_09831_),
    .S(net1836),
    .Z(_09832_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload32 (.I(clknet_2_2_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14205_ (.A1(net1585),
    .A2(_09832_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14206_ (.A1(net1653),
    .A2(net1642),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14207_ (.A1(_09794_),
    .A2(_09807_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14208_ (.A1(_09784_),
    .A2(_09814_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14209_ (.A1(net1666),
    .A2(_09824_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14210_ (.A1(net1660),
    .A2(_09827_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14211_ (.I0(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .I1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .S(net1751),
    .Z(_09834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14212_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net1839),
    .B1(_09834_),
    .B2(net2032),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _14213_ (.I0(_08606_),
    .I1(_09374_),
    .S(net1836),
    .Z(_09835_));
 gf180mcu_fd_sc_mcu9t5v0__inv_20 clkload33 (.I(clknet_2_3_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14215_ (.A1(net1607),
    .A2(_09835_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14216_ (.A1(_09789_),
    .A2(_09832_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14217_ (.A1(_09776_),
    .A2(_09821_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14218_ (.A1(net1653),
    .A2(_09817_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14219_ (.A1(_09798_),
    .A2(net1645),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _14220_ (.I(_09814_),
    .ZN(_09837_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14221_ (.A1(net1603),
    .A2(_09837_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14222_ (.A1(net1657),
    .A2(net1598),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14223_ (.A1(net1667),
    .A2(net1636),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _14224_ (.I(_09674_),
    .ZN(_09838_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14225_ (.A1(_09838_),
    .A2(net1836),
    .ZN(_09839_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14226_ (.A1(net1670),
    .A2(net1583),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14227_ (.A1(net1812),
    .A2(net1811),
    .ZN(_09840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14228_ (.I0(_09840_),
    .I1(net1717),
    .S(net1836),
    .Z(_09841_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload34 (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _14230_ (.A1(_08793_),
    .A2(_09745_),
    .Z(_09843_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14231_ (.A1(net2143),
    .A2(_09749_),
    .B(_09843_),
    .ZN(_09844_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14232_ (.I(net1630),
    .ZN(_09845_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14233_ (.A1(_09841_),
    .A2(_09845_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14234_ (.I0(net2191),
    .I1(_09421_),
    .S(net1836),
    .Z(_09846_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload35 (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14236_ (.A1(net1607),
    .A2(net1629),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14237_ (.A1(net1665),
    .A2(net1634),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14238_ (.A1(net1602),
    .A2(net1635),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14239_ (.A1(_09079_),
    .A2(_09745_),
    .Z(_09848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14240_ (.A1(_07904_),
    .A2(net1838),
    .B(_09848_),
    .ZN(_09849_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload36 (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14242_ (.A1(net1642),
    .A2(net1627),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14243_ (.A1(_07957_),
    .A2(_07961_),
    .A3(_07966_),
    .Z(_09851_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14244_ (.A1(_09223_),
    .A2(_09745_),
    .Z(_09852_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14245_ (.A1(_09851_),
    .A2(net1838),
    .B(_09852_),
    .ZN(_09853_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload37 (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14247_ (.A1(net1650),
    .A2(net1626),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14248_ (.A1(net1655),
    .A2(net1641),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14249_ (.I(net1598),
    .ZN(_09855_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14250_ (.A1(net1605),
    .A2(_09855_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14251_ (.A1(_09784_),
    .A2(net1636),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14252_ (.A1(net2030),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .B1(net1716),
    .B2(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .ZN(_09856_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14253_ (.I(_09856_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14254_ (.A1(net1583),
    .A2(net1630),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14255_ (.A1(net1585),
    .A2(_09841_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14256_ (.A1(net1665),
    .A2(net1629),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14257_ (.A1(_09776_),
    .A2(net1634),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14258_ (.A1(net1601),
    .A2(net1635),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14259_ (.A1(net1645),
    .A2(net1643),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14260_ (.A1(net1650),
    .A2(net1641),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14261_ (.A1(net1655),
    .A2(net1599),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14262_ (.I(net1636),
    .ZN(_09857_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14263_ (.A1(net1605),
    .A2(_09857_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14264_ (.A1(_08649_),
    .A2(net1838),
    .Z(_09858_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14265_ (.A1(_09405_),
    .A2(_09745_),
    .B(_09858_),
    .ZN(_09859_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload38 (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14267_ (.A1(net1657),
    .A2(net1624),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14268_ (.A1(net2030),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A3(_09673_),
    .ZN(_09861_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload39 (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_8 clkload40 (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14271_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(net1716),
    .ZN(_09864_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14272_ (.A1(_09861_),
    .A2(_09864_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload41 (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _14274_ (.A1(net1607),
    .A2(net1583),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14275_ (.A1(_09789_),
    .A2(net1631),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14276_ (.A1(_09776_),
    .A2(net1629),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14277_ (.A1(net1653),
    .A2(net1634),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14278_ (.A1(net1645),
    .A2(net1640),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14279_ (.A1(net1648),
    .A2(net1641),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14280_ (.A1(net1650),
    .A2(net1599),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14281_ (.A1(net1655),
    .A2(net1637),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14282_ (.I(net1624),
    .ZN(_09866_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14283_ (.A1(net1605),
    .A2(_09866_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14284_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(net1716),
    .ZN(_09867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14285_ (.A1(_09861_),
    .A2(_09867_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14286_ (.A1(net1665),
    .A2(net1583),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14287_ (.A1(_09796_),
    .A2(net1631),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14288_ (.A1(net1653),
    .A2(net1629),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14289_ (.A1(net1645),
    .A2(net1639),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14290_ (.A1(net1647),
    .A2(net1641),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14291_ (.A1(net1648),
    .A2(net1599),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14292_ (.A1(net1650),
    .A2(net1637),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14293_ (.A1(net1655),
    .A2(net1624),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14294_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(net1716),
    .ZN(_09868_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14295_ (.A1(_09861_),
    .A2(_09868_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14296_ (.A1(_09776_),
    .A2(net1583),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14297_ (.A1(net1601),
    .A2(net1631),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14298_ (.A1(net1600),
    .A2(net1635),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14299_ (.A1(net1643),
    .A2(net1641),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14300_ (.A1(net1647),
    .A2(net1599),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14301_ (.A1(net1648),
    .A2(net1637),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14302_ (.A1(net1650),
    .A2(net1624),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14303_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(net1716),
    .ZN(_09869_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14304_ (.A1(_09861_),
    .A2(_09869_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14305_ (.A1(net1653),
    .A2(net1583),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14306_ (.A1(_09042_),
    .A2(_09745_),
    .Z(_09870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14307_ (.A1(net1789),
    .A2(_09749_),
    .B(_09870_),
    .ZN(_09871_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14308_ (.I(net1623),
    .ZN(_09872_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14309_ (.A1(net1631),
    .A2(net1594),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14310_ (.A1(net1629),
    .A2(net1628),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14311_ (.A1(net1645),
    .A2(net1634),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14312_ (.A1(net1641),
    .A2(net1640),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14313_ (.A1(net1643),
    .A2(net1599),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14314_ (.A1(net1647),
    .A2(net1637),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14315_ (.A1(net1648),
    .A2(net1624),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14316_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(net1716),
    .ZN(_09873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14317_ (.A1(net1710),
    .A2(_09873_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload42 (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14319_ (.A1(net1583),
    .A2(net1623),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14320_ (.I(net1627),
    .ZN(_09875_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14321_ (.A1(net1631),
    .A2(net1593),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14322_ (.A1(net1645),
    .A2(net1629),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14323_ (.A1(net1641),
    .A2(net1639),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14324_ (.A1(net1640),
    .A2(net1599),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14325_ (.A1(net1643),
    .A2(net1637),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14326_ (.A1(net1647),
    .A2(net1624),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14327_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(net1716),
    .ZN(_09876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14328_ (.A1(net1710),
    .A2(_09876_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14329_ (.A1(net1583),
    .A2(net1627),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14330_ (.A1(net1600),
    .A2(net1631),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14331_ (.A1(net1597),
    .A2(net1635),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14332_ (.A1(net1639),
    .A2(net1599),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14333_ (.A1(net1640),
    .A2(net1637),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14334_ (.A1(net1643),
    .A2(net1624),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14335_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(net1716),
    .ZN(_09877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14336_ (.A1(net1710),
    .A2(_09877_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14337_ (.A1(net1645),
    .A2(net1584),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _14338_ (.A1(_07935_),
    .A2(_07939_),
    .A3(_07944_),
    .Z(_09878_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14339_ (.A1(_09166_),
    .A2(_09745_),
    .Z(_09879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14340_ (.A1(_09878_),
    .A2(_09749_),
    .B(_09879_),
    .ZN(_09880_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14341_ (.I(net1620),
    .ZN(_09881_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14342_ (.A1(net1631),
    .A2(net1592),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14343_ (.A1(net1629),
    .A2(net1626),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14344_ (.A1(net1641),
    .A2(net1634),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14345_ (.A1(_09855_),
    .A2(net1635),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14346_ (.A1(net1639),
    .A2(net1637),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14347_ (.A1(net1640),
    .A2(net1624),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14348_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net1716),
    .ZN(_09882_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14349_ (.A1(net1710),
    .A2(_09882_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1533 (.I(_10262_),
    .Z(net1532));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14351_ (.A1(net1584),
    .A2(net1621),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14352_ (.I(_09853_),
    .ZN(_09884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14353_ (.A1(net1632),
    .A2(net1591),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14354_ (.A1(net1641),
    .A2(net1629),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14355_ (.A1(net1599),
    .A2(net1634),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14356_ (.A1(net1595),
    .A2(net1635),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14357_ (.A1(net1639),
    .A2(net1624),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14358_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net1716),
    .ZN(_09885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14359_ (.A1(net1710),
    .A2(_09885_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14360_ (.A1(net1584),
    .A2(net1626),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14361_ (.A1(net1597),
    .A2(net1632),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14362_ (.A1(net1599),
    .A2(net1629),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14363_ (.A1(net1638),
    .A2(net1634),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14364_ (.A1(net1635),
    .A2(_09866_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14365_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net1716),
    .ZN(_09886_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14366_ (.A1(net1710),
    .A2(_09886_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14367_ (.A1(net1641),
    .A2(net1584),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14368_ (.A1(_09855_),
    .A2(net1632),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14369_ (.A1(net1638),
    .A2(net1629),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14370_ (.A1(net1634),
    .A2(net1624),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14371_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net1716),
    .ZN(_09887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14372_ (.A1(net1710),
    .A2(_09887_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14373_ (.A1(net1599),
    .A2(net1584),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14374_ (.A1(net1595),
    .A2(net1633),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14375_ (.A1(net1629),
    .A2(net1624),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14376_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net1716),
    .ZN(_09888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14377_ (.A1(net1710),
    .A2(_09888_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14378_ (.A1(net1638),
    .A2(net1584),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14379_ (.A1(net1633),
    .A2(_09866_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14380_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net1716),
    .ZN(_09889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14381_ (.A1(net1710),
    .A2(_09889_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14382_ (.A1(net1584),
    .A2(net1624),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14383_ (.A1(_08690_),
    .A2(net1838),
    .Z(_09890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14384_ (.A1(net1719),
    .A2(_09745_),
    .B(_09890_),
    .ZN(_09891_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14385_ (.I(net1619),
    .ZN(_09892_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14386_ (.A1(net1633),
    .A2(_09892_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14387_ (.A1(_09682_),
    .A2(net1839),
    .ZN(_09893_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14388_ (.I(_09893_),
    .ZN(_09894_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14389_ (.A1(net1629),
    .A2(net1582),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14390_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net1716),
    .ZN(_09895_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14391_ (.A1(net1710),
    .A2(_09895_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload44 (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14393_ (.A1(net1584),
    .A2(net1619),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14394_ (.A1(net1633),
    .A2(net1590),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14395_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(net1716),
    .ZN(_09897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14396_ (.A1(net1710),
    .A2(_09897_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14397_ (.A1(net1584),
    .A2(net1582),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _14398_ (.I(net2493),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14399_ (.I(_00750_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14400_ (.A1(_09529_),
    .A2(_09532_),
    .A3(_09533_),
    .A4(_09534_),
    .Z(_09898_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14401_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_09645_),
    .A3(net1826),
    .ZN(_09899_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14402_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(\id_stage_i.controller_i.load_err_q ),
    .Z(_09900_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14403_ (.A1(\id_stage_i.controller_i.exc_req_q ),
    .A2(_09900_),
    .ZN(_09901_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14404_ (.A1(_09898_),
    .A2(_09899_),
    .B(_09901_),
    .ZN(_09902_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14405_ (.I(\cs_registers_i.priv_mode_id_o[1] ),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14406_ (.A1(\cs_registers_i.dcsr_q[12] ),
    .A2(_00953_),
    .ZN(_09903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14407_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_09640_),
    .ZN(_09904_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14408_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_09903_),
    .B(_09904_),
    .ZN(_09905_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14409_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09905_),
    .B(net1932),
    .ZN(_09906_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14410_ (.I(\id_stage_i.controller_i.illegal_insn_q ),
    .ZN(_09907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14411_ (.A1(_09907_),
    .A2(_09620_),
    .ZN(_09908_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14412_ (.A1(_09645_),
    .A2(net1826),
    .A3(_09649_),
    .ZN(_09909_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14413_ (.A1(_09901_),
    .A2(_09906_),
    .A3(_09908_),
    .A4(_09909_),
    .Z(_09910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14414_ (.A1(_09499_),
    .A2(_09910_),
    .Z(_09911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14415_ (.A1(_07631_),
    .A2(_07632_),
    .B(_07645_),
    .ZN(_09912_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _14416_ (.A1(\id_stage_i.id_fsm_q ),
    .A2(_07575_),
    .A3(_09912_),
    .Z(_09913_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14417_ (.A1(_09621_),
    .A2(_09913_),
    .Z(_09914_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14418_ (.I(\id_stage_i.branch_set ),
    .ZN(_09915_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _14419_ (.A1(_09586_),
    .A2(_09587_),
    .A3(_09914_),
    .B(_09915_),
    .ZN(_09916_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14420_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(\id_stage_i.controller_i.instr_fetch_err_i ),
    .ZN(_09917_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14421_ (.A1(net1809),
    .A2(_09917_),
    .Z(_09918_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14422_ (.A1(net65),
    .A2(\cs_registers_i.dcsr_q[2] ),
    .Z(_09919_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14423_ (.I(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .ZN(_09920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14424_ (.A1(_09617_),
    .A2(_09920_),
    .Z(_09921_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14425_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_09921_),
    .Z(_09922_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14426_ (.A1(_09497_),
    .A2(_09922_),
    .Z(_09923_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14427_ (.A1(\cs_registers_i.mie_q[14] ),
    .A2(net140),
    .ZN(_09924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14428_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net146),
    .B1(\cs_registers_i.mie_q[7] ),
    .B2(net147),
    .ZN(_09925_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14429_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net144),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net145),
    .ZN(_09926_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14430_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net142),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net143),
    .ZN(_09927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14431_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net135),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net141),
    .ZN(_09928_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14432_ (.A1(_09925_),
    .A2(_09926_),
    .A3(_09927_),
    .A4(_09928_),
    .Z(_09929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14433_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net138),
    .B1(\cs_registers_i.mie_q[13] ),
    .B2(net139),
    .ZN(_09930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14434_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net136),
    .B1(\cs_registers_i.mie_q[11] ),
    .B2(net137),
    .ZN(_09931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14435_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net148),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net149),
    .ZN(_09932_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14436_ (.A1(_09930_),
    .A2(_09931_),
    .A3(_09932_),
    .Z(_09933_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14437_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(net152),
    .B(net150),
    .ZN(_09934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14438_ (.A1(net134),
    .A2(\cs_registers_i.mie_q[15] ),
    .B1(\cs_registers_i.mie_q[17] ),
    .B2(net151),
    .ZN(_09935_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14439_ (.A1(_09934_),
    .A2(_09935_),
    .Z(_09936_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _14440_ (.A1(_09924_),
    .A2(_09929_),
    .A3(_09933_),
    .A4(_09936_),
    .ZN(_09937_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14441_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_09498_),
    .A3(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_09938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14442_ (.I(\cs_registers_i.nmi_mode_i ),
    .ZN(_09939_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14443_ (.A1(net2038),
    .A2(\cs_registers_i.csr_mstatus_mie_o ),
    .Z(_09940_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14444_ (.A1(_09939_),
    .A2(_09940_),
    .Z(_09941_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14445_ (.I(\cs_registers_i.debug_mode_i ),
    .ZN(_09942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14446_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09942_),
    .Z(_09943_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14447_ (.A1(_09938_),
    .A2(_09941_),
    .A3(_09943_),
    .Z(_09944_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14448_ (.A1(net1808),
    .A2(_09944_),
    .Z(_09945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _14449_ (.A1(_09919_),
    .A2(_09923_),
    .B(_09945_),
    .ZN(_09946_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1532 (.I(_10492_),
    .Z(net1531));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14451_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09498_),
    .B(_09921_),
    .ZN(_09948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14452_ (.A1(_09946_),
    .A2(_09948_),
    .ZN(_09949_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _14453_ (.A1(_09902_),
    .A2(_09911_),
    .B1(_09916_),
    .B2(_09918_),
    .C(_09949_),
    .ZN(_09950_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _14454_ (.A1(_09529_),
    .A2(_09532_),
    .A3(_09533_),
    .A4(_09534_),
    .ZN(_09951_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14455_ (.A1(\id_stage_i.controller_i.exc_req_q ),
    .A2(_09900_),
    .Z(_09952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14456_ (.A1(_09951_),
    .A2(_09646_),
    .B(_09952_),
    .ZN(_09953_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14457_ (.A1(_09617_),
    .A2(_09953_),
    .B(_09497_),
    .ZN(_09954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14458_ (.A1(_09618_),
    .A2(_09954_),
    .B(_09922_),
    .ZN(_09955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload45 (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14460_ (.A1(net1589),
    .A2(net1618),
    .ZN(_09957_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1531 (.I(_10794_),
    .Z(net1530));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload47 (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload48 (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14464_ (.A1(net1809),
    .A2(net176),
    .ZN(_09961_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _14465_ (.A1(_09500_),
    .A2(_09639_),
    .A3(_09899_),
    .A4(_09952_),
    .ZN(_09962_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1530 (.I(_03452_),
    .Z(net1529));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload49 (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _14468_ (.A1(_09499_),
    .A2(_09642_),
    .A3(_09646_),
    .A4(_09901_),
    .Z(_09965_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1529 (.I(_03553_),
    .Z(net1528));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload50 (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1528 (.I(_03906_),
    .Z(net1527));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14472_ (.A1(_09924_),
    .A2(_09929_),
    .A3(_09933_),
    .ZN(_09969_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14473_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(net139),
    .Z(_09970_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14474_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net136),
    .ZN(_09971_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14475_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net2040),
    .Z(_09972_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14476_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(net2042),
    .ZN(_09973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14477_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net2044),
    .Z(_09974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14478_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net2046),
    .ZN(_09975_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14479_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net2047),
    .Z(_09976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14480_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(net2045),
    .B1(_09975_),
    .B2(_09976_),
    .ZN(_09977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14481_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net2043),
    .ZN(_09978_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14482_ (.A1(_09974_),
    .A2(_09977_),
    .B(_09978_),
    .ZN(_09979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14483_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net2041),
    .B1(_09973_),
    .B2(_09979_),
    .ZN(_09980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14484_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(net2039),
    .ZN(_09981_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14485_ (.A1(_09972_),
    .A2(_09980_),
    .B(_09981_),
    .ZN(_09982_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _14486_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(net2049),
    .B1(_09971_),
    .B2(_09982_),
    .ZN(_09983_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14487_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(net2048),
    .B(_09983_),
    .ZN(_09984_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14488_ (.A1(_09970_),
    .A2(_09984_),
    .B(_09924_),
    .ZN(_09985_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14489_ (.A1(net2038),
    .A2(_09939_),
    .ZN(_09986_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14490_ (.A1(_09969_),
    .A2(_09985_),
    .A3(_09986_),
    .ZN(_09987_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14491_ (.A1(_09945_),
    .A2(_09987_),
    .Z(_09988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14492_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[2] ),
    .C(_09988_),
    .ZN(_09989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14493_ (.A1(_09961_),
    .A2(_09989_),
    .ZN(_09990_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14494_ (.A1(_09957_),
    .A2(_09990_),
    .ZN(_09991_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1527 (.I(_03975_),
    .Z(net1526));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload51 (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1526 (.I(_03981_),
    .Z(net1525));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14498_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .A2(net1589),
    .ZN(_09995_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14499_ (.A1(_09991_),
    .A2(_09995_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14500_ (.A1(_09499_),
    .A2(_09952_),
    .Z(_09996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14501_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09996_),
    .Z(_09997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14502_ (.A1(net1809),
    .A2(net1519),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[3] ),
    .C(_09997_),
    .ZN(_09998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14503_ (.I(_09926_),
    .ZN(_09999_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14504_ (.A1(_09999_),
    .A2(_09927_),
    .B(_09925_),
    .ZN(_10000_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14505_ (.A1(_09932_),
    .A2(_10000_),
    .ZN(_10001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14506_ (.A1(_09931_),
    .A2(_10001_),
    .ZN(_10002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14507_ (.A1(net1835),
    .A2(_10002_),
    .ZN(_10003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14508_ (.A1(_09924_),
    .A2(_09986_),
    .Z(_10004_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14509_ (.A1(_09969_),
    .A2(_10003_),
    .A3(_10004_),
    .ZN(_10005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14510_ (.A1(_09945_),
    .A2(_10005_),
    .ZN(_10006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1525 (.I(_04044_),
    .Z(net1524));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14512_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(net1747),
    .ZN(_10008_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _14513_ (.A1(_09998_),
    .A2(_10006_),
    .A3(_10008_),
    .ZN(_10009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14514_ (.A1(_09902_),
    .A2(_09911_),
    .B(_09949_),
    .ZN(_10010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14515_ (.A1(_09916_),
    .A2(_09918_),
    .ZN(_10011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _14516_ (.A1(_10010_),
    .A2(_10011_),
    .ZN(_10012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1524 (.I(_04135_),
    .Z(net1523));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14518_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .I1(_10009_),
    .S(_10012_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14519_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .ZN(_10014_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1523 (.I(_01365_),
    .Z(net1522));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14521_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .ZN(_10016_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload52 (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14523_ (.A1(_10014_),
    .A2(net1589),
    .B(net1834),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload53 (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkload54 (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload55 (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 clkload56 (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14528_ (.A1(net2025),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .Z(_10022_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14529_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .ZN(_10023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14530_ (.A1(_10023_),
    .A2(net112),
    .Z(_10024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14531_ (.A1(net101),
    .A2(_10024_),
    .Z(_10025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14532_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .S(net2025),
    .Z(_10026_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _14533_ (.A1(net2026),
    .A2(_10022_),
    .A3(_10025_),
    .A4(_10026_),
    .Z(_10027_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload57 (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload58 (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1522 (.I(net176),
    .Z(net1521));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14537_ (.A1(net2025),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .Z(_10031_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _14538_ (.A1(_10023_),
    .A2(net109),
    .A3(net108),
    .Z(_10032_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14539_ (.A1(_10031_),
    .A2(_10032_),
    .Z(_10033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14540_ (.A1(_10026_),
    .A2(_10033_),
    .ZN(_10034_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14541_ (.A1(net2026),
    .A2(_10034_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14542_ (.A1(_10027_),
    .A2(_00810_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14543_ (.I(_01132_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14544_ (.I(net154),
    .ZN(_10035_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _14545_ (.A1(net65),
    .A2(core_busy_q),
    .A3(net1808),
    .B(fetch_enable_q),
    .ZN(net155));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14546_ (.A1(_10035_),
    .A2(net155),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1521 (.I(_09706_),
    .Z(net1520));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14548_ (.A1(_09755_),
    .A2(net2475),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14549_ (.A1(net1666),
    .A2(net2475),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14550_ (.A1(_09784_),
    .A2(net2481),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14551_ (.A1(net1606),
    .A2(_09784_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14552_ (.A1(_09794_),
    .A2(net2481),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14553_ (.I(_00990_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14554_ (.A1(net2474),
    .A2(_09803_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14555_ (.A1(net2474),
    .A2(net1642),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14556_ (.A1(net1666),
    .A2(net1627),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14557_ (.A1(_09784_),
    .A2(net1627),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14558_ (.A1(net1668),
    .A2(net1625),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14559_ (.A1(_09817_),
    .A2(net1630),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14560_ (.A1(net1603),
    .A2(_09875_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14561_ (.A1(net1661),
    .A2(net1625),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14562_ (.A1(_09821_),
    .A2(net2481),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14563_ (.A1(_09787_),
    .A2(net1627),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14564_ (.A1(net1666),
    .A2(net1625),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14565_ (.A1(_09832_),
    .A2(_09845_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14566_ (.A1(net1649),
    .A2(net1627),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14567_ (.A1(_09784_),
    .A2(net1625),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14568_ (.A1(_09835_),
    .A2(net2481),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14569_ (.A1(_09776_),
    .A2(_09817_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14570_ (.A1(_09798_),
    .A2(net1627),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14571_ (.A1(net1603),
    .A2(_09884_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14572_ (.A1(net1630),
    .A2(_09846_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14573_ (.A1(net1646),
    .A2(net1627),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14574_ (.A1(net1654),
    .A2(net1625),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14575_ (.A1(net1640),
    .A2(net2477),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14576_ (.A1(net1648),
    .A2(net1621),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14577_ (.A1(net1660),
    .A2(_09891_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1520 (.I(net179),
    .Z(net1519));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14579_ (.A1(net1669),
    .A2(net1582),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14580_ (.A1(net1640),
    .A2(net1628),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14581_ (.A1(net1648),
    .A2(net1626),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14582_ (.A1(net1660),
    .A2(net1582),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14583_ (.A1(net1639),
    .A2(net1628),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14584_ (.A1(net1647),
    .A2(net1626),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14585_ (.A1(net1667),
    .A2(net1582),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14586_ (.A1(net1635),
    .A2(net1593),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14587_ (.A1(net1643),
    .A2(net1626),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14588_ (.A1(net1657),
    .A2(net1582),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14589_ (.A1(net1640),
    .A2(net1626),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14590_ (.A1(net1605),
    .A2(net1590),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14591_ (.A1(net1639),
    .A2(net1626),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14592_ (.A1(net1655),
    .A2(net1582),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14593_ (.A1(net1635),
    .A2(net1591),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14594_ (.A1(net1650),
    .A2(net1582),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14595_ (.A1(net1634),
    .A2(net1626),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14596_ (.A1(net1648),
    .A2(net1582),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14597_ (.A1(net1647),
    .A2(net1582),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14598_ (.A1(net1643),
    .A2(net1582),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14599_ (.A1(net1640),
    .A2(net1582),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14600_ (.A1(net1639),
    .A2(net1582),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14601_ (.A1(net1635),
    .A2(net1590),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14602_ (.A1(net1634),
    .A2(net1582),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14603_ (.A1(net1671),
    .A2(net1660),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14604_ (.A1(net1660),
    .A2(net2475),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14605_ (.A1(net1671),
    .A2(_09784_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14606_ (.A1(net1671),
    .A2(_09787_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14607_ (.A1(net1666),
    .A2(net1664),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14608_ (.A1(net1670),
    .A2(_09794_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14609_ (.A1(net2474),
    .A2(_09798_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14610_ (.A1(net1660),
    .A2(net1622),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14611_ (.I(_00991_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14612_ (.A1(_09798_),
    .A2(net2476),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14613_ (.A1(net1666),
    .A2(net1622),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14614_ (.A1(_09803_),
    .A2(net2476),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14615_ (.A1(_09784_),
    .A2(net2477),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14616_ (.A1(net1642),
    .A2(net2476),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14617_ (.A1(net1603),
    .A2(_09872_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14618_ (.A1(net1661),
    .A2(net1620),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14619_ (.A1(net1670),
    .A2(_09821_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14620_ (.A1(_09787_),
    .A2(net1623),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14621_ (.A1(net1666),
    .A2(net1620),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _14622_ (.I(net1670),
    .ZN(_10037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14623_ (.A1(_10037_),
    .A2(_09832_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14624_ (.A1(net1651),
    .A2(net1623),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14625_ (.A1(_09784_),
    .A2(net1621),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14626_ (.A1(net2474),
    .A2(_09835_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14627_ (.A1(_09798_),
    .A2(net1623),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14628_ (.A1(net1603),
    .A2(_09881_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14629_ (.A1(net2474),
    .A2(_09846_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14630_ (.A1(net1665),
    .A2(_09821_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14631_ (.A1(net1646),
    .A2(net2477),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14632_ (.A1(_09787_),
    .A2(net1620),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14633_ (.A1(_10037_),
    .A2(_09841_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14634_ (.A1(net1642),
    .A2(net1623),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14635_ (.A1(net1649),
    .A2(net1621),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14636_ (.A1(net1653),
    .A2(net1639),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14637_ (.A1(net1646),
    .A2(net1645),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14638_ (.A1(net1667),
    .A2(_09859_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14639_ (.I(_01030_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14640_ (.A1(net1639),
    .A2(net2477),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14641_ (.A1(net1647),
    .A2(net1621),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14642_ (.A1(net1667),
    .A2(net1619),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14643_ (.A1(net1635),
    .A2(net1594),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14644_ (.A1(net1643),
    .A2(net1621),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14645_ (.A1(net1657),
    .A2(net1619),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14646_ (.A1(net1634),
    .A2(net2477),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14647_ (.A1(net1640),
    .A2(net1621),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14648_ (.A1(net1605),
    .A2(_09892_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14649_ (.A1(net1634),
    .A2(net1628),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14650_ (.A1(net1639),
    .A2(net1621),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14651_ (.A1(net1655),
    .A2(net1619),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14652_ (.A1(net1635),
    .A2(net1592),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14653_ (.A1(net1650),
    .A2(net1619),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14654_ (.A1(net1634),
    .A2(net1621),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14655_ (.A1(net1648),
    .A2(net1619),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14656_ (.A1(net1629),
    .A2(net1621),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14657_ (.A1(net1647),
    .A2(net1619),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14658_ (.A1(net1643),
    .A2(net1619),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14659_ (.A1(net1640),
    .A2(net1619),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14660_ (.A1(net1639),
    .A2(net1619),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14661_ (.A1(net1635),
    .A2(_09892_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14662_ (.A1(net1634),
    .A2(net1619),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14663_ (.A1(net1629),
    .A2(net1619),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14664_ (.A1(net1671),
    .A2(net1666),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14665_ (.A1(_10037_),
    .A2(net1604),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14666_ (.A1(net1604),
    .A2(_09845_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14667_ (.A1(net1660),
    .A2(net1659),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14668_ (.A1(_09787_),
    .A2(net1630),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14669_ (.A1(_09755_),
    .A2(net1627),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14670_ (.A1(net1660),
    .A2(net1627),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14671_ (.A1(net1670),
    .A2(_09817_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14672_ (.A1(net1629),
    .A2(net2477),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14673_ (.I(_00103_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14674_ (.I(_00123_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14675_ (.I(_00233_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14676_ (.I(_00260_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14677_ (.I(_00036_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14678_ (.I(_00057_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14679_ (.I(_00070_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14680_ (.I(_00078_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14681_ (.I(_00094_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14682_ (.I(_00115_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14683_ (.I(_00137_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14684_ (.I(_00161_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14685_ (.I(_00177_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14686_ (.I(_00189_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14687_ (.I(_00213_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14688_ (.I(_00226_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14689_ (.I(_00254_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14690_ (.I(_00274_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14691_ (.I(_00285_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14692_ (.I(_00297_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14693_ (.I(_00302_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14694_ (.I(_00316_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14695_ (.I(_00323_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14696_ (.I(_00331_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14697_ (.I(_00339_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14698_ (.I(_00344_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14699_ (.I(_00359_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14700_ (.I(_00374_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14701_ (.I(_00379_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14702_ (.I(_00394_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14703_ (.I(_00405_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14704_ (.I(_00410_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14705_ (.I(_00414_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14706_ (.I(_00429_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14707_ (.I(_00440_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14708_ (.I(_00451_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14709_ (.I(_00465_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14710_ (.I(_00476_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14711_ (.I(_00482_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14712_ (.I(_00489_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14713_ (.I(_00500_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14714_ (.I(_00511_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14715_ (.I(_00518_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14716_ (.I(_00522_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14717_ (.I(_00533_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14718_ (.I(_00544_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14719_ (.I(_00550_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14720_ (.I(_00553_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14721_ (.I(_00565_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14722_ (.I(_00576_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14723_ (.I(_00587_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14724_ (.I(_00592_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14725_ (.I(_00597_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14726_ (.I(_00610_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14727_ (.I(_00616_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14728_ (.I(_00622_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14729_ (.I(_00627_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14730_ (.I(_00641_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14731_ (.I(_00648_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14732_ (.I(_00651_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14733_ (.I(_00656_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14734_ (.I(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14735_ (.I(_00677_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14736_ (.I(_00682_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14737_ (.I(_00696_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14738_ (.I(_00703_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14739_ (.I(_00707_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14740_ (.I(_00720_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14741_ (.I(_00726_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14742_ (.I(_00729_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14743_ (.I(_00742_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14744_ (.I(_00753_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14745_ (.I(_00758_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14746_ (.I(_00765_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14747_ (.I(_00773_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14748_ (.I(_00778_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14749_ (.I(_00785_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14750_ (.I(_00795_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14751_ (.I(_00803_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14752_ (.I(_00047_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14753_ (.I(_00114_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14754_ (.I(_00136_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14755_ (.I(_00160_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14756_ (.I(_00174_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14757_ (.I(_00176_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14758_ (.I(_00188_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14759_ (.I(_00212_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14760_ (.I(_00273_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14761_ (.I(_00296_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14762_ (.I(_00301_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14763_ (.I(_00315_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14764_ (.I(_00330_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14765_ (.I(_00338_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14766_ (.I(_00343_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14767_ (.I(_00358_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14768_ (.I(_00373_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14769_ (.I(_00378_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14770_ (.I(_00393_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14771_ (.I(_00404_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14772_ (.I(_00413_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14773_ (.I(_00428_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14774_ (.I(_00439_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14775_ (.I(_00446_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14776_ (.I(_00448_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14777_ (.I(_00450_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14778_ (.I(_00464_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14779_ (.I(_00475_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14780_ (.I(_00488_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14781_ (.I(_00499_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14782_ (.I(_00510_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14783_ (.I(_00517_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14784_ (.I(_00521_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14785_ (.I(_00532_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14786_ (.I(_00543_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14787_ (.I(_00552_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14788_ (.I(_00564_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14789_ (.I(_00575_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14790_ (.I(_00582_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14791_ (.I(_00586_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14792_ (.I(_00591_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14793_ (.I(_00596_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14794_ (.I(_00609_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14795_ (.I(_00621_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14796_ (.I(_00626_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14797_ (.I(_00640_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14798_ (.I(_00647_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14799_ (.I(_00650_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14800_ (.I(_00655_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14801_ (.I(_00669_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14802_ (.I(_00676_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14803_ (.I(_00681_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14804_ (.I(_00695_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14805_ (.I(_00702_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14806_ (.I(_00706_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14807_ (.I(_00719_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14808_ (.I(_00728_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14809_ (.I(_00741_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14810_ (.I(_00748_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14811_ (.I(_00752_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14812_ (.I(_00757_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14813_ (.I(_00764_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14814_ (.I(_00772_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14815_ (.I(_00784_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 clkload61 (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14817_ (.A1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A2(net1823),
    .Z(_10039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14818_ (.I0(_01145_),
    .I1(_10039_),
    .S(net1814),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14819_ (.A1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A2(net1823),
    .Z(_10040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14820_ (.I0(_01151_),
    .I1(_10040_),
    .S(net1814),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14821_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(net1823),
    .Z(_10041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14822_ (.I0(_01158_),
    .I1(_10041_),
    .S(net1814),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14823_ (.A1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A2(net1823),
    .Z(_10042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14824_ (.I0(_01165_),
    .I1(_10042_),
    .S(net1814),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14825_ (.A1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A2(net1823),
    .Z(_10043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14826_ (.I0(_01172_),
    .I1(_10043_),
    .S(net1814),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14827_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(net1823),
    .Z(_10044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14828_ (.I0(net1691),
    .I1(_10044_),
    .S(net1814),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14829_ (.A1(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A2(net1823),
    .Z(_10045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14830_ (.I0(net1690),
    .I1(_10045_),
    .S(net1814),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14831_ (.A1(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .A2(net1823),
    .Z(_10046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14832_ (.I0(_01193_),
    .I1(_10046_),
    .S(net1814),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14833_ (.A1(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .A2(net1823),
    .Z(_10047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14834_ (.I0(net1689),
    .I1(_10047_),
    .S(net1814),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14835_ (.A1(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A2(net1823),
    .Z(_10048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload59 (.I(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14837_ (.I0(net1688),
    .I1(_10048_),
    .S(net1814),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload60 (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14839_ (.A1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .A2(net1823),
    .Z(_10051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14840_ (.I0(net1695),
    .I1(_10051_),
    .S(net1814),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14841_ (.A1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A2(net1823),
    .Z(_10052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14842_ (.I0(_01226_),
    .I1(_10052_),
    .S(net1814),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14843_ (.A1(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .A2(net1823),
    .Z(_10053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14844_ (.I0(_01228_),
    .I1(_10053_),
    .S(net1814),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14845_ (.A1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A2(net1823),
    .Z(_10054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14846_ (.I0(net1685),
    .I1(_10054_),
    .S(net1814),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14847_ (.A1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A2(net1823),
    .Z(_10055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14848_ (.I0(net1684),
    .I1(_10055_),
    .S(net1814),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14849_ (.A1(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .A2(net1823),
    .Z(_10056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14850_ (.I0(net1683),
    .I1(_10056_),
    .S(net1814),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14851_ (.A1(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .A2(net1823),
    .Z(_10057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14852_ (.I0(_01256_),
    .I1(_10057_),
    .S(net1814),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14853_ (.A1(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .A2(net1823),
    .Z(_10058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14854_ (.I0(net1682),
    .I1(_10058_),
    .S(net1814),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14855_ (.A1(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .A2(net1823),
    .Z(_10059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14856_ (.I0(net1681),
    .I1(_10059_),
    .S(net1814),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14857_ (.A1(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .A2(net1823),
    .Z(_10060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload67 (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14859_ (.I0(_01277_),
    .I1(_10060_),
    .S(net1814),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload62 (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14861_ (.A1(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .A2(net1823),
    .Z(_10063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14862_ (.I0(net1680),
    .I1(_10063_),
    .S(net1815),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14863_ (.A1(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .A2(net1823),
    .Z(_10064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14864_ (.I0(net1679),
    .I1(_10064_),
    .S(net1815),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14865_ (.A1(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .A2(net1823),
    .Z(_10065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14866_ (.I0(net1678),
    .I1(_10065_),
    .S(net1815),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14867_ (.A1(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .A2(net1823),
    .Z(_10066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14868_ (.I0(net1677),
    .I1(_10066_),
    .S(net1815),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14869_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net1823),
    .Z(_10067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14870_ (.I0(_01312_),
    .I1(_10067_),
    .S(net1815),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14871_ (.A1(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .A2(net1823),
    .Z(_10068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14872_ (.I0(_01319_),
    .I1(_10068_),
    .S(net1814),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14873_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net1823),
    .Z(_10069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14874_ (.I0(_01326_),
    .I1(_10069_),
    .S(net1814),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14875_ (.A1(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .A2(net1823),
    .Z(_10070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14876_ (.I0(net1676),
    .I1(_10070_),
    .S(net1814),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14877_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net1823),
    .Z(_10071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14878_ (.I0(net1675),
    .I1(_10071_),
    .S(net1814),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _14879_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(net1823),
    .Z(_10072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14880_ (.I0(_01347_),
    .I1(_10072_),
    .S(net1814),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload66 (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload65 (.I(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14883_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14884_ (.I(_00015_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14885_ (.A1(_09755_),
    .A2(net1664),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14886_ (.I(_00038_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14887_ (.A1(net1660),
    .A2(net1652),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14888_ (.I(_00061_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14889_ (.I(_00080_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14890_ (.I(_00075_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14891_ (.A1(net1668),
    .A2(net1644),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14892_ (.I(_00120_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14893_ (.I(_00099_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14894_ (.A1(net1668),
    .A2(net1620),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14895_ (.I(_00127_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14896_ (.I(_00126_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14897_ (.I(_00147_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14898_ (.I(_00143_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14899_ (.I(_00150_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14900_ (.A1(net1668),
    .A2(_09824_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14901_ (.I(_00195_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14902_ (.I(_00200_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14903_ (.I(_00204_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14904_ (.I(_00256_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14905_ (.I(_00228_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14906_ (.A1(net1669),
    .A2(_09859_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14907_ (.I(_00236_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14908_ (.A1(net1669),
    .A2(_09891_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14909_ (.I(_00263_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14910_ (.I(_00321_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14911_ (.I(_00327_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14912_ (.I(_00289_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14913_ (.I(_00371_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14914_ (.I(_00366_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14915_ (.I(_00370_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14916_ (.I(_00401_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14917_ (.I(_00407_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14918_ (.I(_00436_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14919_ (.I(_00443_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14920_ (.I(_00472_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14921_ (.I(_00479_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14922_ (.I(_00507_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14923_ (.I(_00514_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14924_ (.I(_00540_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14925_ (.I(_00547_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14926_ (.I(_00572_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14927_ (.I(_00579_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14928_ (.I(_00606_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14929_ (.I(_00613_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14930_ (.I(_00637_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14931_ (.I(_00644_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14932_ (.I(_00666_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14933_ (.I(_00673_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _14934_ (.I(_00584_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14935_ (.I(_00692_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14936_ (.I(_00699_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14937_ (.I(_00716_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14938_ (.I(_00723_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14939_ (.I(_00738_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14940_ (.I(_00745_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14941_ (.I(_00761_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14942_ (.I(_00749_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14943_ (.I(_00769_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14944_ (.I(_00781_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14945_ (.I(_00789_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14946_ (.I(net2150),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14947_ (.A1(_09498_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .ZN(_10074_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14948_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(_09921_),
    .ZN(_10075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14949_ (.A1(_10074_),
    .A2(_10075_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_10076_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload64 (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload63 (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _14952_ (.A1(net2023),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(_09950_),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .ZN(_10079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14953_ (.A1(_10076_),
    .A2(_10079_),
    .ZN(_10080_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14954_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_10080_),
    .Z(_10081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _14955_ (.I(_10081_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14956_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net2185),
    .ZN(_10082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14957_ (.A1(net2028),
    .A2(net1786),
    .B(_10082_),
    .ZN(_10083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14958_ (.I0(net2119),
    .I1(net1694),
    .S(_07742_),
    .Z(_10084_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14959_ (.A1(_08187_),
    .A2(_10083_),
    .B(_10084_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14960_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .B2(_08197_),
    .ZN(_10085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14961_ (.A1(_07804_),
    .A2(_08228_),
    .B1(net1780),
    .B2(net2028),
    .C(_10085_),
    .ZN(_10086_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _14962_ (.A1(_08187_),
    .A2(_10086_),
    .Z(_10087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14963_ (.I0(net1694),
    .I1(net2119),
    .S(_07808_),
    .Z(_10088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _14964_ (.A1(_10087_),
    .A2(_10088_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14965_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .B2(_08197_),
    .ZN(_10089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14966_ (.A1(net1794),
    .A2(_08228_),
    .B1(_08315_),
    .B2(net2028),
    .C(_10089_),
    .ZN(_10090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_20 clkload68 (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14968_ (.I0(net1694),
    .I1(net2119),
    .S(_07831_),
    .Z(_10092_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14969_ (.A1(_08187_),
    .A2(_10090_),
    .B(_10092_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14970_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .B2(net1824),
    .ZN(_10093_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _14971_ (.A1(net1792),
    .A2(_08200_),
    .ZN(_10094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _14972_ (.A1(net2028),
    .A2(net1778),
    .B(_10093_),
    .C(_10094_),
    .ZN(_10095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14973_ (.I0(net2119),
    .I1(net1694),
    .S(_01173_),
    .Z(_10096_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14974_ (.A1(_08187_),
    .A2(_10095_),
    .B(_10096_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14975_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1790),
    .ZN(_10097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14976_ (.A1(net2028),
    .A2(net1777),
    .B(_10097_),
    .ZN(_10098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14977_ (.I0(net2119),
    .I1(net1694),
    .S(_01180_),
    .Z(_10099_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14978_ (.A1(_08187_),
    .A2(_10098_),
    .B(_10099_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14979_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .B2(net1824),
    .ZN(_10100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14980_ (.A1(_09549_),
    .A2(_08228_),
    .B1(net1776),
    .B2(net2028),
    .C(_10100_),
    .ZN(_10101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14981_ (.I0(net1694),
    .I1(_08218_),
    .S(_01191_),
    .Z(_10102_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14982_ (.A1(_08187_),
    .A2(_10101_),
    .B(_10102_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14983_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .B2(_08197_),
    .ZN(_10103_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14984_ (.A1(_07924_),
    .A2(_08228_),
    .B1(net1775),
    .B2(net2028),
    .C(_10103_),
    .ZN(_10104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14985_ (.I0(_08218_),
    .I1(net1694),
    .S(_07925_),
    .Z(_10105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14986_ (.A1(_08187_),
    .A2(_10104_),
    .B(_10105_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14987_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .B2(_08197_),
    .ZN(_10106_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14988_ (.A1(_07945_),
    .A2(_08228_),
    .B1(net2174),
    .B2(net2028),
    .C(_10106_),
    .ZN(_10107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14989_ (.I0(_08218_),
    .I1(net1694),
    .S(_07946_),
    .Z(_10108_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14990_ (.A1(_08187_),
    .A2(_10107_),
    .B(_10108_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _14991_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .B2(_08197_),
    .ZN(_10109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _14992_ (.A1(_07967_),
    .A2(_08228_),
    .B1(net1735),
    .B2(net2028),
    .C(_10109_),
    .ZN(_10110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14993_ (.I0(_08218_),
    .I1(net1694),
    .S(net1697),
    .Z(_10111_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14994_ (.A1(_08187_),
    .A2(_10110_),
    .B(_10111_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14995_ (.A1(net1841),
    .A2(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net2158),
    .ZN(_10112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _14996_ (.A1(net2028),
    .A2(net1738),
    .B(_10112_),
    .ZN(_10113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _14997_ (.I0(net1693),
    .I1(net1694),
    .S(_07997_),
    .Z(_10114_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _14998_ (.A1(_08187_),
    .A2(_10113_),
    .B(_10114_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _14999_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1755),
    .ZN(_10115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15000_ (.A1(net2028),
    .A2(net1754),
    .B(_10115_),
    .ZN(_10116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15001_ (.I0(net2175),
    .I1(net2111),
    .S(_01341_),
    .Z(_10117_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15002_ (.A1(_08187_),
    .A2(_10116_),
    .B(_10117_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _15003_ (.A1(_08192_),
    .A2(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .B1(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .B2(net1824),
    .C1(_08200_),
    .C2(net1753),
    .ZN(_10118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15004_ (.A1(net2028),
    .A2(net1752),
    .B(_10118_),
    .ZN(_10119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15005_ (.I0(net2175),
    .I1(net2111),
    .S(_01348_),
    .Z(_10120_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15006_ (.A1(_08187_),
    .A2(_10119_),
    .B(_10120_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_1_core_clock (.I(delaynet_0_core_clock),
    .Z(delaynet_1_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_0_core_clock (.I(clk_i),
    .Z(delaynet_0_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15009_ (.A1(net1698),
    .A2(_09627_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15010_ (.A1(net1699),
    .A2(_09627_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15011_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15012_ (.I(_00016_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15013_ (.I(_00020_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15014_ (.A1(net1606),
    .A2(net1660),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15015_ (.I(_00029_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15016_ (.I(_00028_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15017_ (.A1(_09755_),
    .A2(net1652),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15018_ (.I(_00050_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15019_ (.A1(_09755_),
    .A2(net1622),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15020_ (.I(_00049_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15021_ (.I(_00076_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15022_ (.I(_00060_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15023_ (.I(_00100_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15024_ (.I(_00107_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15025_ (.A1(net1660),
    .A2(net1644),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15026_ (.I(_00106_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15027_ (.I(_00148_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15028_ (.I(_00151_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15029_ (.I(_00170_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15030_ (.I(_00179_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15031_ (.A1(net1661),
    .A2(_09814_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15032_ (.I(_00205_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15033_ (.I(_00229_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15034_ (.I(_00202_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15035_ (.I(_00237_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15036_ (.I(_00219_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15037_ (.I(_00264_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15038_ (.A1(net1660),
    .A2(_09859_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15039_ (.I(_00290_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15040_ (.A1(net2030),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B1(net1716),
    .B2(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .ZN(_10123_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15041_ (.I(_10123_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15042_ (.I(_00287_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15043_ (.I(_00333_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15044_ (.I(_00367_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15045_ (.I(_00402_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15046_ (.I(_00361_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15047_ (.I(_00408_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15048_ (.I(_00437_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15049_ (.I(_00396_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15050_ (.I(_00444_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15051_ (.I(_00473_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15052_ (.I(_00431_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15053_ (.I(_00480_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15054_ (.I(_00508_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15055_ (.I(_00467_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15056_ (.I(_00515_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15057_ (.I(_00541_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15058_ (.I(_00502_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15059_ (.I(_00548_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15060_ (.I(_00573_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15061_ (.I(_00535_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15062_ (.I(_00580_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15063_ (.I(_00607_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15064_ (.I(_00567_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15065_ (.I(_00614_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15066_ (.I(_00638_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15067_ (.I(_00600_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15068_ (.I(_00645_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15069_ (.I(_00667_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15070_ (.I(_00631_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15071_ (.I(_00674_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15072_ (.I(_00693_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15073_ (.I(_00660_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15074_ (.I(_00700_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15075_ (.I(_00717_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15076_ (.I(_00685_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15077_ (.I(_00724_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15078_ (.I(_00739_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15079_ (.I(_00709_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15080_ (.I(_00746_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15081_ (.I(_00762_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15082_ (.I(_00731_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15083_ (.I(_00770_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15084_ (.I(_00782_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15085_ (.I(_00790_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15086_ (.I(_00808_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15087_ (.I(net2068),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15088_ (.I(net2096),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15089_ (.I(net2176),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15090_ (.I(_01243_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15091_ (.I(_01250_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15092_ (.I(_01257_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15093_ (.I(net2482),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15094_ (.I(_01271_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15095_ (.I(_01278_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15096_ (.I(_01285_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15097_ (.I(_01292_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15098_ (.I(_01299_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15099_ (.I(_01306_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15100_ (.I(_01313_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15101_ (.I(_01320_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15102_ (.I(_01327_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15103_ (.I(_01334_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1519 (.I(_10268_),
    .Z(net1518));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15105_ (.I(_00989_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15106_ (.I(_00993_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15107_ (.I(_01003_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15108_ (.I(_01007_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15109_ (.I(_01019_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15110_ (.I(_01025_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15111_ (.I(_01031_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15112_ (.I(_00978_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15113_ (.I(_00983_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15114_ (.I(_00997_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15115_ (.I(_01014_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15116_ (.I(_01037_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15117_ (.A1(_07566_),
    .A2(_07557_),
    .Z(_10124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15118_ (.A1(_07711_),
    .A2(_10124_),
    .Z(_10125_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15119_ (.A1(_08121_),
    .A2(_10125_),
    .Z(_10126_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_2_core_clock (.I(delaynet_1_core_clock),
    .Z(delaynet_2_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15121_ (.A1(_07599_),
    .A2(_09699_),
    .Z(_10128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15122_ (.A1(_10125_),
    .A2(_10128_),
    .Z(_10129_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15123_ (.A1(_07652_),
    .A2(_10129_),
    .B(net2099),
    .ZN(_10130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15124_ (.A1(_07553_),
    .A2(net31),
    .ZN(_10131_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15125_ (.A1(_10130_),
    .A2(_10131_),
    .Z(_10132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15126_ (.I0(_10126_),
    .I1(\load_store_unit_i.data_type_q[2] ),
    .S(_10132_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15127_ (.A1(_08158_),
    .A2(_10125_),
    .Z(_10133_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_3_core_clock (.I(delaynet_2_core_clock),
    .Z(delaynet_3_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15129_ (.I0(_10133_),
    .I1(\load_store_unit_i.data_type_q[1] ),
    .S(_10132_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15130_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .S(_09688_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15131_ (.I0(net2032),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_09688_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 delaybuf_4_core_clock (.I(delaynet_3_core_clock),
    .Z(delaynet_4_core_clock));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1518 (.I(_10754_),
    .Z(net1517));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15134_ (.I0(net2031),
    .I1(net2029),
    .S(_09700_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1517 (.I(_10773_),
    .Z(net1516));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15136_ (.A1(_09699_),
    .A2(net1750),
    .ZN(_10138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15137_ (.I0(net2028),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .S(_10138_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15138_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .S(_10138_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15139_ (.I(net1705),
    .ZN(_10139_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2052 (.I(net178),
    .Z(net2051));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15141_ (.I(_00950_),
    .ZN(_10141_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2053 (.I(net2177),
    .Z(net2052));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2054 (.I(net2177),
    .Z(net2053));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15144_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01139_),
    .Z(_10144_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15145_ (.A1(_10139_),
    .A2(_10144_),
    .ZN(_10145_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15146_ (.A1(net1611),
    .A2(_01159_),
    .B(_09627_),
    .ZN(_10146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15147_ (.A1(_01166_),
    .A2(_09627_),
    .ZN(_10147_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15148_ (.A1(_10146_),
    .A2(_10147_),
    .ZN(_10148_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _15149_ (.A1(net1703),
    .A2(net1586),
    .A3(_09627_),
    .Z(_10149_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2055 (.I(_08549_),
    .Z(net2054));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer2056 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(net2055));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15152_ (.I(\cs_registers_i.mhpmcounter[1856] ),
    .ZN(_10152_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2057 (.I(net2057),
    .Z(net2056));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15154_ (.A1(net1702),
    .A2(_09627_),
    .Z(_10154_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15155_ (.A1(net1612),
    .A2(_07773_),
    .A3(_10154_),
    .A4(_09544_),
    .ZN(_10155_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 split2058 (.I(_08942_),
    .Z(net2057));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15157_ (.A1(_07859_),
    .A2(net1610),
    .A3(_09627_),
    .Z(_10157_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15158_ (.A1(_09575_),
    .A2(_09553_),
    .A3(_10157_),
    .Z(_10158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15159_ (.A1(_10155_),
    .A2(_10158_),
    .ZN(_10159_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 rebuffer2059 (.I(net2156),
    .Z(net2058));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15161_ (.A1(_09551_),
    .A2(_09553_),
    .A3(_10157_),
    .Z(_10161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15162_ (.A1(_10155_),
    .A2(_10161_),
    .ZN(_10162_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2060 (.I(_08548_),
    .Z(net2059));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15164_ (.I(\cs_registers_i.mhpmcounter[1888] ),
    .ZN(_10164_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15165_ (.A1(_10152_),
    .A2(_10159_),
    .B1(_10162_),
    .B2(_10164_),
    .ZN(_10165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15166_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .ZN(_10166_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2062 (.I(net1799),
    .Z(net2061));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15168_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .ZN(_10168_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15169_ (.A1(net1700),
    .A2(_09627_),
    .Z(_10169_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15170_ (.A1(net1699),
    .A2(net1698),
    .A3(_01212_),
    .A4(_09627_),
    .Z(_10170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15171_ (.A1(net1696),
    .A2(_09575_),
    .A3(_10170_),
    .Z(_10171_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15172_ (.A1(_07773_),
    .A2(_09590_),
    .A3(_09591_),
    .ZN(_10172_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15173_ (.A1(_10169_),
    .A2(_10171_),
    .A3(_10172_),
    .ZN(_10173_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _15174_ (.A1(_10166_),
    .A2(_10159_),
    .B1(_10162_),
    .B2(_10168_),
    .C(_10173_),
    .ZN(_10174_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15175_ (.A1(_09562_),
    .A2(_09563_),
    .A3(_09567_),
    .B(_09627_),
    .ZN(_10175_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15176_ (.A1(_10149_),
    .A2(_10165_),
    .B1(_10174_),
    .B2(_10175_),
    .ZN(_10176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15177_ (.A1(net1700),
    .A2(_09568_),
    .Z(_10177_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15178_ (.A1(net1701),
    .A2(_10177_),
    .A3(_09577_),
    .A4(_09579_),
    .Z(_10178_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15179_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(_10178_),
    .ZN(_10179_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15180_ (.A1(net1611),
    .A2(_09568_),
    .A3(_10154_),
    .Z(_10180_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15181_ (.A1(net1701),
    .A2(_09625_),
    .ZN(_10181_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15182_ (.A1(net1610),
    .A2(_09628_),
    .A3(_09603_),
    .A4(_10181_),
    .Z(_10182_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15183_ (.A1(_10180_),
    .A2(_10182_),
    .Z(_10183_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer2061 (.I(_08548_),
    .Z(net2060));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2064 (.I(_07610_),
    .Z(net2063));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15186_ (.A1(_09628_),
    .A2(_09629_),
    .A3(_09630_),
    .Z(_10186_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15187_ (.A1(net1612),
    .A2(net1586),
    .A3(_07773_),
    .A4(_10154_),
    .Z(_10187_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15188_ (.A1(_10186_),
    .A2(_10187_),
    .Z(_10188_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2063 (.I(_00861_),
    .Z(net2062));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2067 (.I(_07715_),
    .Z(net2066));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15191_ (.A1(_01198_),
    .A2(_01205_),
    .A3(net1697),
    .A4(_09625_),
    .Z(_10191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15192_ (.A1(net1701),
    .A2(_07859_),
    .B(_09625_),
    .ZN(_10192_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15193_ (.A1(net1610),
    .A2(_09602_),
    .A3(_10191_),
    .A4(_10192_),
    .Z(_10193_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15194_ (.A1(net1703),
    .A2(_09562_),
    .A3(_09563_),
    .A4(_09589_),
    .Z(_10194_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15195_ (.A1(net1702),
    .A2(_09627_),
    .ZN(_10195_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15196_ (.A1(_07773_),
    .A2(_10194_),
    .A3(_10195_),
    .Z(_10196_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15197_ (.A1(_10193_),
    .A2(_10196_),
    .ZN(_10197_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1516 (.I(_03458_),
    .Z(net1515));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15199_ (.A1(net67),
    .A2(net1563),
    .B1(_10188_),
    .B2(\cs_registers_i.dscratch1_q[0] ),
    .C(_10197_),
    .ZN(_10199_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15200_ (.A1(net1611),
    .A2(_01159_),
    .A3(_09598_),
    .B(_09627_),
    .ZN(_10200_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15201_ (.A1(_10186_),
    .A2(_10200_),
    .Z(_10201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2066 (.I(net2204),
    .Z(net2065));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15203_ (.A1(_10146_),
    .A2(_10186_),
    .A3(_10149_),
    .Z(_10203_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2065 (.I(net2063),
    .Z(net2064));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2068 (.I(_07715_),
    .Z(net2067));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15206_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[0] ),
    .ZN(_10206_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15207_ (.A1(_10179_),
    .A2(_10199_),
    .A3(_10206_),
    .Z(_10207_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15208_ (.A1(_07859_),
    .A2(_01180_),
    .A3(net2068),
    .A4(_09627_),
    .Z(_10208_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15209_ (.A1(net1701),
    .A2(net1696),
    .A3(_10170_),
    .A4(_10208_),
    .Z(_10209_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2070 (.I(net1800),
    .Z(net2069));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15211_ (.A1(_10209_),
    .A2(_10187_),
    .Z(_10211_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2069 (.I(_01191_),
    .Z(net2068));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1515 (.I(_04155_),
    .Z(net1514));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15214_ (.A1(_10146_),
    .A2(_10209_),
    .A3(_10149_),
    .Z(_10214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15215_ (.A1(\cs_registers_i.mtval_q[0] ),
    .A2(_10211_),
    .B1(_10214_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .ZN(_10215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15216_ (.A1(_10209_),
    .A2(_10200_),
    .Z(_10216_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1514 (.I(_06906_),
    .Z(net1513));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15218_ (.A1(_07773_),
    .A2(_09569_),
    .A3(_10154_),
    .Z(_10218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15219_ (.A1(_10209_),
    .A2(_10218_),
    .Z(_10219_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2071 (.I(_01228_),
    .Z(net2070));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15221_ (.A1(\cs_registers_i.mscratch_q[0] ),
    .A2(net1554),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_10221_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15222_ (.A1(_10215_),
    .A2(_10221_),
    .Z(_10222_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15223_ (.A1(_10148_),
    .A2(_10176_),
    .B(_10207_),
    .C(_10222_),
    .ZN(_10223_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15224_ (.A1(_01139_),
    .A2(_10223_),
    .Z(_10224_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15225_ (.A1(_10145_),
    .A2(_10224_),
    .Z(_10225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15226_ (.A1(net1697),
    .A2(net1610),
    .Z(_10226_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15227_ (.A1(_10226_),
    .A2(_09622_),
    .A3(_09588_),
    .Z(_10227_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15228_ (.A1(_09584_),
    .A2(_09616_),
    .B(_10227_),
    .C(_09636_),
    .ZN(_10228_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1513 (.I(net183),
    .Z(net1512));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15230_ (.A1(_10178_),
    .A2(net1535),
    .Z(_10230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15231_ (.I0(\cs_registers_i.mcountinhibit_q[0] ),
    .I1(_10225_),
    .S(_10230_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15232_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01151_),
    .Z(_10231_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2072 (.I(_00821_),
    .Z(net2071));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2073 (.I(_01193_),
    .Z(net2072));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15235_ (.A1(\cs_registers_i.mtval_q[2] ),
    .A2(_10211_),
    .B1(_10214_),
    .B2(\cs_registers_i.mcause_q[2] ),
    .C1(_10219_),
    .C2(\cs_registers_i.csr_mepc_o[2] ),
    .ZN(_10234_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2074 (.I(_00849_),
    .Z(net2073));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _15237_ (.A1(net1610),
    .A2(_09602_),
    .A3(_10191_),
    .A4(_10192_),
    .ZN(_10236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15238_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[2] ),
    .C1(_10218_),
    .C2(_10236_),
    .ZN(_10237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15239_ (.A1(\cs_registers_i.mscratch_q[2] ),
    .A2(_10216_),
    .ZN(_10238_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15240_ (.A1(_10186_),
    .A2(_10218_),
    .Z(_10239_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2075 (.I(_08741_),
    .Z(net2074));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2077 (.I(_00877_),
    .Z(net2076));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15243_ (.A1(\cs_registers_i.dscratch1_q[2] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[2] ),
    .C1(net89),
    .C2(net1563),
    .ZN(_10242_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15244_ (.A1(_10238_),
    .A2(_10242_),
    .Z(_10243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15245_ (.A1(_07773_),
    .A2(_10154_),
    .Z(_10244_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15246_ (.A1(net1701),
    .A2(_10177_),
    .A3(_10171_),
    .A4(_10244_),
    .Z(_10245_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2076 (.I(_07993_),
    .Z(net2075));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15248_ (.A1(_10146_),
    .A2(_10147_),
    .Z(_10247_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2078 (.I(net2076),
    .Z(net2077));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 clone2079 (.I(net2090),
    .Z(net2078));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2081 (.I(_08386_),
    .Z(net2080));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2080 (.I(_00873_),
    .Z(net2079));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15253_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1858] ),
    .ZN(_10252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15254_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1890] ),
    .ZN(_10253_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1512 (.I(_10374_),
    .Z(net1511));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15256_ (.A1(_10159_),
    .A2(_10252_),
    .B1(_10253_),
    .B2(_10162_),
    .ZN(_10255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15257_ (.A1(\cs_registers_i.mcountinhibit_q[2] ),
    .A2(_10245_),
    .B1(net1562),
    .B2(_10255_),
    .ZN(_10256_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15258_ (.A1(_10234_),
    .A2(_10237_),
    .A3(_10243_),
    .A4(_10256_),
    .Z(_10257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15259_ (.A1(_10139_),
    .A2(_10231_),
    .B1(_10257_),
    .B2(_01155_),
    .ZN(_10258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15260_ (.I0(\cs_registers_i.mcountinhibit_q[2] ),
    .I1(_10258_),
    .S(_10230_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2082 (.I(\load_store_unit_i.ls_fsm_cs[2] ),
    .Z(net2081));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15262_ (.I(_09601_),
    .ZN(_10260_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15263_ (.A1(_09558_),
    .A2(_10260_),
    .Z(_10261_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15264_ (.A1(_09615_),
    .A2(net1608),
    .A3(_10228_),
    .A4(_10261_),
    .Z(_10262_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15265_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(net1532),
    .Z(_10263_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15266_ (.A1(_09612_),
    .A2(_09613_),
    .A3(_09614_),
    .ZN(_10264_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15267_ (.A1(_10264_),
    .A2(net1535),
    .ZN(_10265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15268_ (.A1(net1532),
    .A2(_10265_),
    .ZN(_10266_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15269_ (.A1(_10263_),
    .A2(_10266_),
    .ZN(_10267_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15270_ (.A1(\cs_registers_i.mcountinhibit_q[0] ),
    .A2(net1532),
    .ZN(_10268_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1511 (.I(_10855_),
    .Z(net1510));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1510 (.I(_10859_),
    .Z(net1509));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15273_ (.A1(net1532),
    .A2(_10265_),
    .Z(_10271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2083 (.I(_00845_),
    .Z(net2082));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15275_ (.A1(_01139_),
    .A2(_10223_),
    .B(_10145_),
    .ZN(_10273_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15276_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(net1518),
    .B1(_10271_),
    .B2(_10273_),
    .ZN(_10274_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15277_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .A2(_10267_),
    .B(_10274_),
    .ZN(_10275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15278_ (.I(_10275_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1508 (.I(_04571_),
    .Z(net1507));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1506 (.I(_05501_),
    .Z(net1505));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1505 (.I(_05592_),
    .Z(net1504));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15282_ (.I0(_00950_),
    .I1(_08009_),
    .S(net2102),
    .Z(_10279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15283_ (.A1(\cs_registers_i.mtval_q[10] ),
    .A2(net1555),
    .Z(_10280_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1503 (.I(_05610_),
    .Z(net1502));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15285_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(_10197_),
    .Z(_10282_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15286_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(net1553),
    .Z(_10283_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1502 (.I(_06466_),
    .Z(net1501));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1504 (.I(_05610_),
    .Z(net1503));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1501 (.I(net182),
    .Z(net1500));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15290_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1866] ),
    .ZN(_10287_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1507 (.I(net1505),
    .Z(net1506));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15292_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1898] ),
    .ZN(_10289_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15293_ (.A1(_10159_),
    .A2(_10287_),
    .B1(_10289_),
    .B2(net1560),
    .ZN(_10290_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15294_ (.A1(net1562),
    .A2(_10290_),
    .ZN(_10291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15295_ (.A1(\cs_registers_i.dscratch0_q[10] ),
    .A2(net1556),
    .ZN(_10292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15296_ (.A1(\cs_registers_i.dscratch1_q[10] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C1(net68),
    .C2(net1563),
    .ZN(_10293_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2085 (.I(_09489_),
    .Z(net2084));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2086 (.I(_09113_),
    .Z(net2085));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15299_ (.A1(\cs_registers_i.mscratch_q[10] ),
    .A2(_10216_),
    .B(_10245_),
    .ZN(_10296_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15300_ (.A1(_10291_),
    .A2(_10292_),
    .A3(_10293_),
    .A4(_10296_),
    .ZN(_10297_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15301_ (.A1(_10280_),
    .A2(_10282_),
    .A3(_10283_),
    .A4(_10297_),
    .Z(_10298_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15302_ (.A1(net1705),
    .A2(_10279_),
    .B1(_10298_),
    .B2(net2102),
    .ZN(_10299_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15303_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .Z(_10300_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15304_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .Z(_10301_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15305_ (.A1(_01369_),
    .A2(_10300_),
    .A3(_10301_),
    .Z(_10302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15306_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(_10302_),
    .ZN(_10303_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _15307_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(_10303_),
    .ZN(_10304_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15308_ (.A1(net1518),
    .A2(_10304_),
    .ZN(_10305_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15309_ (.A1(_10263_),
    .A2(_10266_),
    .Z(_10306_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15310_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .A2(_10306_),
    .ZN(_10307_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15311_ (.A1(_10266_),
    .A2(_10299_),
    .B(_10305_),
    .C(_10307_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15312_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .ZN(_10308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15313_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .Z(_10309_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15314_ (.A1(_10300_),
    .A2(_10301_),
    .A3(_10309_),
    .Z(_10310_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15315_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ),
    .Z(_10311_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15316_ (.A1(_10310_),
    .A2(_10311_),
    .Z(_10312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15317_ (.I0(_10271_),
    .I1(_10312_),
    .S(net1518),
    .Z(_10313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15318_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2159),
    .Z(_10314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15319_ (.A1(_10139_),
    .A2(_10314_),
    .ZN(_10315_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15320_ (.I(\cs_registers_i.mtval_q[11] ),
    .ZN(_10316_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15321_ (.A1(net1701),
    .A2(net1696),
    .A3(_10170_),
    .A4(_10208_),
    .ZN(_10317_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15322_ (.A1(net1611),
    .A2(_10195_),
    .A3(_09590_),
    .Z(_10318_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15323_ (.I(\cs_registers_i.csr_mtvec_o[11] ),
    .ZN(_10319_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _15324_ (.A1(_10316_),
    .A2(_10317_),
    .A3(_10318_),
    .B1(_10193_),
    .B2(_10196_),
    .B3(_10319_),
    .ZN(_10320_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15325_ (.A1(\cs_registers_i.mie_q[15] ),
    .A2(_10180_),
    .A3(_10236_),
    .Z(_10321_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15326_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_10209_),
    .A3(_10218_),
    .Z(_10322_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15327_ (.A1(_10320_),
    .A2(_10321_),
    .A3(_10322_),
    .Z(_10323_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15328_ (.A1(\cs_registers_i.mstatus_q[2] ),
    .A2(_10200_),
    .A3(_10236_),
    .Z(_10324_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15329_ (.A1(net2050),
    .A2(_10180_),
    .A3(_10209_),
    .Z(_10325_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15330_ (.A1(\cs_registers_i.mscratch_q[11] ),
    .A2(_10209_),
    .A3(_10200_),
    .Z(_10326_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15331_ (.A1(_10245_),
    .A2(_10324_),
    .A3(_10325_),
    .A4(_10326_),
    .Z(_10327_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15332_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_10175_),
    .Z(_10328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15333_ (.A1(net1703),
    .A2(_09541_),
    .Z(_10329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15334_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(net1586),
    .A3(_10329_),
    .Z(_10330_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15335_ (.A1(_10328_),
    .A2(_10330_),
    .B(_10155_),
    .C(_10161_),
    .ZN(_10331_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15336_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A2(_10175_),
    .Z(_10332_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15337_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(net1586),
    .A3(_10329_),
    .Z(_10333_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15338_ (.A1(_10332_),
    .A2(_10333_),
    .B(_10155_),
    .C(_10158_),
    .ZN(_10334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15339_ (.A1(_10331_),
    .A2(_10334_),
    .B(_10148_),
    .ZN(_10335_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15340_ (.A1(\cs_registers_i.dscratch1_q[11] ),
    .A2(_10186_),
    .A3(_10187_),
    .Z(_10336_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15341_ (.I(net69),
    .ZN(_10337_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15342_ (.A1(_07773_),
    .A2(_09598_),
    .A3(_10195_),
    .Z(_10338_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15343_ (.A1(net1610),
    .A2(_09628_),
    .A3(_09603_),
    .A4(_10181_),
    .ZN(_10339_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15344_ (.A1(net1611),
    .A2(_10194_),
    .A3(_10195_),
    .Z(_10340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15345_ (.I(\cs_registers_i.csr_depc_o[11] ),
    .ZN(_10341_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _15346_ (.A1(_10337_),
    .A2(_10338_),
    .A3(_10339_),
    .B1(_10340_),
    .B2(_09631_),
    .B3(_10341_),
    .ZN(_10342_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15347_ (.A1(\cs_registers_i.dcsr_q[11] ),
    .A2(_10186_),
    .A3(_10200_),
    .Z(_10343_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15348_ (.A1(\cs_registers_i.dscratch0_q[11] ),
    .A2(_10146_),
    .A3(_10186_),
    .A4(_10149_),
    .Z(_10344_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15349_ (.A1(_10336_),
    .A2(_10342_),
    .A3(_10343_),
    .A4(_10344_),
    .Z(_10345_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15350_ (.A1(_10323_),
    .A2(_10327_),
    .A3(_10335_),
    .A4(_10345_),
    .Z(_10346_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15351_ (.A1(net2159),
    .A2(_10346_),
    .Z(_10347_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15352_ (.A1(_10315_),
    .A2(_10347_),
    .Z(_10348_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15353_ (.A1(_10308_),
    .A2(net1518),
    .A3(_10312_),
    .Z(_10349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15354_ (.A1(_10271_),
    .A2(_10348_),
    .B(_10349_),
    .ZN(_10350_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15355_ (.A1(_10308_),
    .A2(_10313_),
    .B(_10350_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15356_ (.A1(_10159_),
    .A2(net1560),
    .ZN(_10351_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15357_ (.A1(_10338_),
    .A2(_10317_),
    .B(_09626_),
    .ZN(_10352_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15358_ (.A1(net1701),
    .A2(net1696),
    .A3(_09629_),
    .A4(_10170_),
    .Z(_10353_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15359_ (.A1(_07859_),
    .A2(_01180_),
    .A3(_09627_),
    .Z(_10354_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15360_ (.A1(_09628_),
    .A2(_10354_),
    .A3(_09544_),
    .A4(_09545_),
    .Z(_10355_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15361_ (.A1(_10209_),
    .A2(_10353_),
    .A3(_10355_),
    .Z(_10356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15362_ (.A1(_10352_),
    .A2(_10356_),
    .Z(_10357_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15363_ (.A1(net1701),
    .A2(_09570_),
    .A3(_10171_),
    .A4(_10244_),
    .Z(_10358_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15364_ (.I(_10171_),
    .ZN(_10359_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15365_ (.A1(_07773_),
    .A2(_10194_),
    .B(_09598_),
    .C(_09627_),
    .ZN(_10360_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15366_ (.A1(_09625_),
    .A2(_09593_),
    .Z(_10361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15367_ (.A1(_10169_),
    .A2(_10172_),
    .B1(_10360_),
    .B2(_10361_),
    .ZN(_10362_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15368_ (.A1(_10158_),
    .A2(_10161_),
    .B(_10155_),
    .ZN(_10363_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15369_ (.A1(net1699),
    .A2(net1698),
    .A3(_09627_),
    .Z(_10364_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15370_ (.A1(_10364_),
    .A2(_09629_),
    .A3(_09630_),
    .Z(_10365_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15371_ (.A1(net1611),
    .A2(_01159_),
    .B(net1697),
    .C(_09627_),
    .ZN(_10366_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15372_ (.A1(_10180_),
    .A2(_10182_),
    .B1(_10365_),
    .B2(_10366_),
    .ZN(_10367_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15373_ (.A1(_10359_),
    .A2(_10362_),
    .B(_10363_),
    .C(_10367_),
    .ZN(_10368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15374_ (.I(_09636_),
    .ZN(_10369_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15375_ (.A1(_10357_),
    .A2(_10358_),
    .A3(_10368_),
    .B(_10369_),
    .ZN(_10370_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15376_ (.A1(_10226_),
    .A2(_09622_),
    .A3(_09625_),
    .Z(_10371_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15377_ (.A1(_10370_),
    .A2(_10371_),
    .ZN(_10372_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer2087 (.I(\load_store_unit_i.ls_fsm_cs[1] ),
    .Z(net2086));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15379_ (.A1(_10175_),
    .A2(_10351_),
    .A3(_10372_),
    .A4(net1562),
    .ZN(_10374_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2088 (.I(net2086),
    .Z(net2087));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _15381_ (.I(\cs_registers_i.mcountinhibit_q[0] ),
    .ZN(_10376_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15382_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A2(_10376_),
    .Z(_10377_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15383_ (.A1(_10302_),
    .A2(_10311_),
    .A3(_10377_),
    .Z(_10378_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15384_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_10378_),
    .Z(_10379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15385_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1704),
    .Z(_10380_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15386_ (.I(\cs_registers_i.mtval_q[12] ),
    .ZN(_10381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15387_ (.I(\cs_registers_i.csr_mtvec_o[12] ),
    .ZN(_10382_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _15388_ (.A1(_10381_),
    .A2(_10317_),
    .A3(_10318_),
    .B1(_10193_),
    .B2(_10196_),
    .B3(_10382_),
    .ZN(_10383_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15389_ (.A1(\cs_registers_i.mstatus_q[3] ),
    .A2(_10200_),
    .A3(_10236_),
    .Z(_10384_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15390_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(_10209_),
    .A3(_10218_),
    .Z(_10385_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15391_ (.A1(_10383_),
    .A2(_10384_),
    .A3(_10385_),
    .Z(_10386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15392_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_10175_),
    .Z(_10387_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15393_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(net1586),
    .A3(_10329_),
    .Z(_10388_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15394_ (.A1(_10387_),
    .A2(_10388_),
    .B(_10155_),
    .C(_10161_),
    .ZN(_10389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15395_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_10175_),
    .Z(_10390_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15396_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(net1586),
    .A3(_10329_),
    .Z(_10391_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15397_ (.A1(_10390_),
    .A2(_10391_),
    .B(_10155_),
    .C(_10158_),
    .ZN(_10392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15398_ (.A1(_10389_),
    .A2(_10392_),
    .B(_10148_),
    .ZN(_10393_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15399_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_10186_),
    .A3(_10218_),
    .Z(_10394_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15400_ (.I(net70),
    .ZN(_10395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15401_ (.I(\cs_registers_i.dscratch1_q[12] ),
    .ZN(_10396_));
 gf180mcu_fd_sc_mcu9t5v0__oai33_2 _15402_ (.A1(_10395_),
    .A2(_10338_),
    .A3(_10339_),
    .B1(_10318_),
    .B2(_09631_),
    .B3(_10396_),
    .ZN(_10397_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15403_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_10146_),
    .A3(_10186_),
    .A4(_10149_),
    .Z(_10398_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15404_ (.A1(\cs_registers_i.dcsr_q[12] ),
    .A2(_10186_),
    .A3(_10200_),
    .Z(_10399_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15405_ (.A1(_10394_),
    .A2(_10397_),
    .A3(_10398_),
    .A4(_10399_),
    .Z(_10400_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15406_ (.A1(\cs_registers_i.mscratch_q[12] ),
    .A2(_10209_),
    .A3(_10200_),
    .Z(_10401_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15407_ (.A1(_10358_),
    .A2(_10401_),
    .Z(_10402_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15408_ (.A1(_10386_),
    .A2(_10393_),
    .A3(_10400_),
    .A4(_10402_),
    .Z(_10403_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15409_ (.A1(net1705),
    .A2(_10380_),
    .B1(_10403_),
    .B2(net1704),
    .ZN(_10404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15410_ (.A1(_09627_),
    .A2(_09598_),
    .Z(_10405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15411_ (.A1(_07859_),
    .A2(_09627_),
    .Z(_10406_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15412_ (.A1(net1699),
    .A2(net1610),
    .A3(_10406_),
    .A4(_09576_),
    .Z(_10407_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15413_ (.A1(_09551_),
    .A2(_09575_),
    .B(_10155_),
    .C(_10407_),
    .ZN(_10408_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15414_ (.A1(net1701),
    .A2(_10171_),
    .A3(_10244_),
    .Z(_10409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15415_ (.A1(_09570_),
    .A2(_10409_),
    .ZN(_10410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15416_ (.A1(_01187_),
    .A2(_10354_),
    .Z(_10411_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15417_ (.A1(net1696),
    .A2(_09628_),
    .A3(_09544_),
    .A4(_10411_),
    .Z(_10412_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15418_ (.A1(_10209_),
    .A2(_10353_),
    .A3(_10412_),
    .B(_10352_),
    .ZN(_10413_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15419_ (.A1(_10359_),
    .A2(_10362_),
    .Z(_10414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15420_ (.A1(net1610),
    .A2(_09628_),
    .Z(_10415_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15421_ (.A1(_10180_),
    .A2(_10415_),
    .A3(_09603_),
    .A4(_10181_),
    .ZN(_10416_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15422_ (.A1(_01166_),
    .A2(net1696),
    .A3(_09629_),
    .Z(_10417_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15423_ (.A1(_10364_),
    .A2(_10417_),
    .A3(_10366_),
    .ZN(_10418_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15424_ (.A1(_10408_),
    .A2(_10416_),
    .A3(_10418_),
    .Z(_10419_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15425_ (.A1(_10410_),
    .A2(_10413_),
    .A3(_10414_),
    .A4(_10419_),
    .Z(_10420_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15426_ (.A1(_09636_),
    .A2(_10420_),
    .A3(_10371_),
    .Z(_10421_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15427_ (.A1(_10405_),
    .A2(_10408_),
    .A3(_10421_),
    .A4(_10148_),
    .Z(_10422_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15428_ (.A1(_09551_),
    .A2(_10155_),
    .A3(_10407_),
    .ZN(_10423_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15429_ (.A1(_10423_),
    .A2(_10421_),
    .ZN(_10424_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15430_ (.A1(_10422_),
    .A2(_10424_),
    .ZN(_10425_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 split2089 (.I(_00865_),
    .Z(net2088));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1500 (.I(net181),
    .Z(net1499));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15433_ (.I0(_10378_),
    .I1(_10265_),
    .S(net1532),
    .Z(_10428_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15434_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_10428_),
    .ZN(_10429_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15435_ (.A1(net1511),
    .A2(_10379_),
    .B1(_10404_),
    .B2(_10425_),
    .C(_10429_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15436_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2070),
    .Z(_10430_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15437_ (.A1(_10139_),
    .A2(_10430_),
    .Z(_10431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15438_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(net1555),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[13] ),
    .C1(_10197_),
    .C2(\cs_registers_i.csr_mtvec_o[13] ),
    .ZN(_10432_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 rebuffer2091 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .Z(net2090));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1498 (.I(_04697_),
    .Z(net1497));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15441_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1869] ),
    .ZN(_10435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15442_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1901] ),
    .ZN(_10436_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15443_ (.A1(_10159_),
    .A2(_10435_),
    .B1(_10436_),
    .B2(net1560),
    .ZN(_10437_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15444_ (.A1(net1562),
    .A2(_10437_),
    .ZN(_10438_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1497 (.I(_05046_),
    .Z(net1496));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1495 (.I(_05574_),
    .Z(net1494));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1496 (.I(_05574_),
    .Z(net1495));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15448_ (.A1(\cs_registers_i.dscratch1_q[13] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[13] ),
    .C1(net71),
    .C2(net1563),
    .ZN(_10442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15449_ (.A1(\cs_registers_i.dcsr_q[13] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[13] ),
    .ZN(_10443_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15450_ (.A1(_10442_),
    .A2(_10443_),
    .Z(_10444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15451_ (.A1(\cs_registers_i.csr_mepc_o[13] ),
    .A2(net1553),
    .B(_10245_),
    .ZN(_10445_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15452_ (.A1(_10432_),
    .A2(_10438_),
    .A3(_10444_),
    .A4(_10445_),
    .Z(_10446_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15453_ (.A1(_01232_),
    .A2(_10446_),
    .Z(_10447_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15454_ (.A1(_10431_),
    .A2(_10447_),
    .Z(_10448_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15455_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(_10312_),
    .A3(_10377_),
    .ZN(_10449_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15456_ (.A1(_10264_),
    .A2(net1535),
    .Z(_10450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15457_ (.I0(_10449_),
    .I1(_10450_),
    .S(net1532),
    .Z(_10451_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15458_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(_10451_),
    .ZN(_10452_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15459_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(net1532),
    .A3(_10449_),
    .Z(_10453_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15460_ (.A1(_10266_),
    .A2(_10448_),
    .B(_10452_),
    .C(_10453_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15461_ (.A1(_10155_),
    .A2(_10161_),
    .Z(_10454_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15462_ (.A1(_10454_),
    .A2(_10372_),
    .Z(_10455_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15463_ (.A1(net1511),
    .A2(_10455_),
    .ZN(_10456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15464_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1685),
    .Z(_10457_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15465_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(net1555),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .C1(_10197_),
    .C2(\cs_registers_i.csr_mtvec_o[14] ),
    .ZN(_10458_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15466_ (.I(_10458_),
    .ZN(_10459_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1494 (.I(_05579_),
    .Z(net1493));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1493 (.I(_05584_),
    .Z(net1492));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15469_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1870] ),
    .ZN(_10462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15470_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1902] ),
    .ZN(_10463_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15471_ (.A1(_10159_),
    .A2(_10462_),
    .B1(_10463_),
    .B2(net1560),
    .ZN(_10464_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15472_ (.A1(net1562),
    .A2(_10464_),
    .ZN(_10465_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15473_ (.A1(\cs_registers_i.dscratch0_q[14] ),
    .A2(net1556),
    .ZN(_10466_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15474_ (.A1(\cs_registers_i.dscratch1_q[14] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[14] ),
    .C1(net72),
    .C2(net1563),
    .ZN(_10467_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1492 (.I(_05596_),
    .Z(net1491));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15476_ (.A1(\cs_registers_i.mscratch_q[14] ),
    .A2(_10216_),
    .B(_10245_),
    .ZN(_10469_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15477_ (.A1(_10465_),
    .A2(_10466_),
    .A3(_10467_),
    .A4(_10469_),
    .ZN(_10470_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15478_ (.A1(_10459_),
    .A2(_10470_),
    .Z(_10471_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15479_ (.A1(net1705),
    .A2(_10457_),
    .B1(_10471_),
    .B2(net1685),
    .ZN(_10472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15480_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(_10379_),
    .ZN(_10473_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15481_ (.A1(_10175_),
    .A2(_10454_),
    .A3(_10372_),
    .A4(net1562),
    .Z(_10474_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15482_ (.A1(net1511),
    .A2(_10473_),
    .B(_10474_),
    .ZN(_10475_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15483_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A2(_10475_),
    .ZN(_10476_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15484_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .A3(net1511),
    .A4(_10379_),
    .Z(_10477_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15485_ (.A1(_10456_),
    .A2(_10472_),
    .B(_10476_),
    .C(_10477_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15486_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1684),
    .Z(_10478_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15487_ (.A1(\cs_registers_i.mtval_q[15] ),
    .A2(net1555),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[15] ),
    .C1(_10197_),
    .C2(\cs_registers_i.csr_mtvec_o[15] ),
    .ZN(_10479_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1491 (.I(_05600_),
    .Z(net1490));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15489_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1871] ),
    .ZN(_10481_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15490_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1903] ),
    .ZN(_10482_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15491_ (.A1(_10159_),
    .A2(_10481_),
    .B1(_10482_),
    .B2(net1560),
    .ZN(_10483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15492_ (.A1(net1562),
    .A2(_10483_),
    .ZN(_10484_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15493_ (.A1(\cs_registers_i.dscratch1_q[15] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[15] ),
    .C1(net73),
    .C2(net1563),
    .ZN(_10485_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15494_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[15] ),
    .ZN(_10486_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15495_ (.A1(_10485_),
    .A2(_10486_),
    .Z(_10487_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2092 (.I(net2090),
    .Z(net2091));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1499 (.I(_04697_),
    .Z(net1498));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15498_ (.A1(\cs_registers_i.csr_mepc_o[15] ),
    .A2(net1553),
    .B(_10245_),
    .ZN(_10490_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15499_ (.A1(_10479_),
    .A2(_10484_),
    .A3(_10487_),
    .A4(_10490_),
    .Z(_10491_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15500_ (.A1(_10139_),
    .A2(_10478_),
    .B1(_10491_),
    .B2(_01246_),
    .ZN(_10492_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1490 (.I(_05602_),
    .Z(net1489));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15502_ (.A1(_10425_),
    .A2(net1531),
    .ZN(_10494_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15503_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ),
    .Z(_10495_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15504_ (.A1(_10311_),
    .A2(_10495_),
    .Z(_10496_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15505_ (.A1(_10310_),
    .A2(_10496_),
    .Z(_10497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15506_ (.A1(net1518),
    .A2(_10497_),
    .ZN(_10498_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2093 (.I(_08098_),
    .Z(net2092));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15508_ (.I0(_10271_),
    .I1(_10497_),
    .S(net1518),
    .Z(_10500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15509_ (.I0(_10498_),
    .I1(_10500_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .Z(_10501_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15510_ (.A1(_10494_),
    .A2(_10501_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15511_ (.A1(net1511),
    .A2(_10455_),
    .Z(_10502_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1489 (.I(_05606_),
    .Z(net1488));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1488 (.I(_05614_),
    .Z(net1487));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15514_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1683),
    .Z(_10505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15515_ (.A1(_10139_),
    .A2(_10505_),
    .ZN(_10506_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15516_ (.A1(_10180_),
    .A2(_10209_),
    .Z(_10507_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1487 (.I(_05619_),
    .Z(net1486));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1481 (.I(_05664_),
    .Z(net1480));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15519_ (.A1(net135),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[16] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[16] ),
    .ZN(_10510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15520_ (.A1(\cs_registers_i.mtval_q[16] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[16] ),
    .ZN(_10511_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15521_ (.A1(_10180_),
    .A2(_10236_),
    .Z(_10512_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1479 (.I(_05675_),
    .Z(net1478));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15523_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15524_ (.A1(_10511_),
    .A2(_10514_),
    .Z(_10515_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15525_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1872] ),
    .ZN(_10516_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15526_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1904] ),
    .ZN(_10517_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15527_ (.A1(net1561),
    .A2(_10516_),
    .B1(_10517_),
    .B2(net1560),
    .ZN(_10518_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15528_ (.A1(net1562),
    .A2(_10518_),
    .ZN(_10519_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15529_ (.A1(\cs_registers_i.dscratch0_q[16] ),
    .A2(net1556),
    .ZN(_10520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15530_ (.A1(\cs_registers_i.dscratch1_q[16] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .C1(net74),
    .C2(net1563),
    .ZN(_10521_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15531_ (.A1(_10520_),
    .A2(_10521_),
    .Z(_10522_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15532_ (.A1(_10510_),
    .A2(_10515_),
    .A3(_10519_),
    .A4(_10522_),
    .ZN(_10523_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15533_ (.A1(net1683),
    .A2(_10523_),
    .Z(_10524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15534_ (.A1(_10506_),
    .A2(_10524_),
    .ZN(_10525_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15535_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_10302_),
    .A3(_10496_),
    .Z(_10526_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15536_ (.A1(net1518),
    .A2(_10526_),
    .ZN(_10527_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15537_ (.A1(_10263_),
    .A2(_10526_),
    .ZN(_10528_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15538_ (.A1(_10306_),
    .A2(_10528_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .ZN(_10529_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _15539_ (.A1(_10502_),
    .A2(_10525_),
    .B1(_10527_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .C(_10529_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15540_ (.I0(_00950_),
    .I1(_08009_),
    .S(_01256_),
    .Z(_10530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15541_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(net1553),
    .B1(_10197_),
    .B2(\cs_registers_i.csr_mtvec_o[17] ),
    .ZN(_10531_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15542_ (.A1(\cs_registers_i.mtval_q[17] ),
    .A2(net1555),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[17] ),
    .ZN(_10532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15543_ (.A1(_10531_),
    .A2(_10532_),
    .Z(_10533_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15544_ (.A1(net2047),
    .A2(_10507_),
    .B1(_10512_),
    .B2(\cs_registers_i.mie_q[1] ),
    .ZN(_10534_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15545_ (.A1(_10200_),
    .A2(_10236_),
    .Z(_10535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15546_ (.A1(\cs_registers_i.mstatus_q[1] ),
    .A2(_10535_),
    .B(_10245_),
    .ZN(_10536_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15547_ (.A1(_10534_),
    .A2(_10536_),
    .Z(_10537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15548_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1873] ),
    .ZN(_10538_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15549_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1905] ),
    .ZN(_10539_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15550_ (.A1(net1561),
    .A2(_10538_),
    .B1(_10539_),
    .B2(net1560),
    .ZN(_10540_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15551_ (.A1(net1562),
    .A2(_10540_),
    .ZN(_10541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15552_ (.A1(\cs_registers_i.dscratch0_q[17] ),
    .A2(net1556),
    .ZN(_10542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15553_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .C1(net75),
    .C2(net1563),
    .ZN(_10543_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15554_ (.A1(_10542_),
    .A2(_10543_),
    .Z(_10544_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15555_ (.A1(_10533_),
    .A2(_10537_),
    .A3(_10541_),
    .A4(_10544_),
    .ZN(_10545_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15556_ (.A1(net1705),
    .A2(_10530_),
    .B1(_10545_),
    .B2(_01256_),
    .ZN(_10546_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15557_ (.A1(_10376_),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A4(_10497_),
    .ZN(_10547_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15558_ (.A1(net1511),
    .A2(_10547_),
    .B(_10474_),
    .ZN(_10548_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15559_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A2(_10548_),
    .ZN(_10549_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15560_ (.I(_10547_),
    .ZN(_10550_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15561_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A2(net1511),
    .A3(_10550_),
    .Z(_10551_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15562_ (.A1(_10456_),
    .A2(_10546_),
    .B(_10549_),
    .C(_10551_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15563_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1682),
    .Z(_10552_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15564_ (.A1(_10139_),
    .A2(_10552_),
    .ZN(_10553_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15565_ (.A1(net2046),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[18] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[18] ),
    .ZN(_10554_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15566_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[18] ),
    .ZN(_10555_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15567_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10556_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15568_ (.A1(_10555_),
    .A2(_10556_),
    .Z(_10557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15569_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1874] ),
    .ZN(_10558_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15570_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1906] ),
    .ZN(_10559_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15571_ (.A1(net1561),
    .A2(_10558_),
    .B1(_10559_),
    .B2(net1560),
    .ZN(_10560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15572_ (.A1(net1562),
    .A2(_10560_),
    .ZN(_10561_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15573_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(net1556),
    .ZN(_10562_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15574_ (.A1(\cs_registers_i.dscratch1_q[18] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .C1(net76),
    .C2(net1563),
    .ZN(_10563_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15575_ (.A1(_10562_),
    .A2(_10563_),
    .Z(_10564_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15576_ (.A1(_10554_),
    .A2(_10557_),
    .A3(_10561_),
    .A4(_10564_),
    .ZN(_10565_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15577_ (.A1(net1682),
    .A2(_10565_),
    .Z(_10566_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15578_ (.A1(_10553_),
    .A2(_10566_),
    .ZN(_10567_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15579_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A3(_10526_),
    .ZN(_10568_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15580_ (.A1(net1518),
    .A2(_10568_),
    .Z(_10569_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15581_ (.A1(_10306_),
    .A2(_10569_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .ZN(_10570_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15582_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .A2(_10263_),
    .A3(_10568_),
    .Z(_10571_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15583_ (.A1(_10266_),
    .A2(_10567_),
    .B(_10570_),
    .C(_10571_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15584_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1681),
    .Z(_10572_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15585_ (.A1(_10139_),
    .A2(_10572_),
    .ZN(_10573_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15586_ (.A1(net2045),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[19] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[19] ),
    .ZN(_10574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15587_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[19] ),
    .ZN(_10575_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15588_ (.A1(\cs_registers_i.mie_q[3] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10576_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15589_ (.A1(_10575_),
    .A2(_10576_),
    .Z(_10577_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15590_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1875] ),
    .ZN(_10578_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15591_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1907] ),
    .ZN(_10579_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15592_ (.A1(net1561),
    .A2(_10578_),
    .B1(_10579_),
    .B2(net1560),
    .ZN(_10580_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15593_ (.A1(net1562),
    .A2(_10580_),
    .ZN(_10581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15594_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(net1556),
    .ZN(_10582_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15595_ (.A1(\cs_registers_i.dscratch1_q[19] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[19] ),
    .C1(net77),
    .C2(net1563),
    .ZN(_10583_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15596_ (.A1(_10582_),
    .A2(_10583_),
    .Z(_10584_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15597_ (.A1(_10574_),
    .A2(_10577_),
    .A3(_10581_),
    .A4(_10584_),
    .ZN(_10585_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15598_ (.A1(net1681),
    .A2(_10585_),
    .Z(_10586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15599_ (.A1(_10573_),
    .A2(_10586_),
    .Z(_10587_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15600_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ),
    .Z(_10588_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15601_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(_10310_),
    .A3(_10496_),
    .A4(_10588_),
    .Z(_10589_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _15602_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(_10589_),
    .Z(_10590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15603_ (.A1(_10271_),
    .A2(_10587_),
    .B1(_10590_),
    .B2(net1518),
    .ZN(_10591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15604_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(_10306_),
    .ZN(_10592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15605_ (.A1(_10591_),
    .A2(_10592_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15606_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .ZN(_10593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15607_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01145_),
    .Z(_10594_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15608_ (.A1(_10139_),
    .A2(_10594_),
    .ZN(_10595_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15609_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(_10211_),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .ZN(_10596_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15610_ (.A1(\cs_registers_i.mcause_q[1] ),
    .A2(_10214_),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[1] ),
    .ZN(_10597_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15611_ (.A1(_10596_),
    .A2(_10597_),
    .Z(_10598_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15612_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1857] ),
    .ZN(_10599_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15613_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1889] ),
    .ZN(_10600_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15614_ (.A1(_10159_),
    .A2(_10599_),
    .B1(_10600_),
    .B2(_10162_),
    .ZN(_10601_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15615_ (.A1(net1562),
    .A2(_10601_),
    .ZN(_10602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15616_ (.A1(\cs_registers_i.dscratch1_q[1] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[1] ),
    .C1(net78),
    .C2(net1563),
    .ZN(_10603_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15617_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[1] ),
    .ZN(_10604_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15618_ (.A1(_10598_),
    .A2(_10602_),
    .A3(_10603_),
    .A4(_10604_),
    .ZN(_10605_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15619_ (.A1(_01145_),
    .A2(_10605_),
    .Z(_10606_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15620_ (.A1(_10595_),
    .A2(_10606_),
    .Z(_10607_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15621_ (.A1(_01370_),
    .A2(_10263_),
    .B1(_10266_),
    .B2(_10607_),
    .ZN(_10608_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15622_ (.A1(_10593_),
    .A2(_10306_),
    .B(_10608_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15623_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2135),
    .Z(_10609_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15624_ (.A1(_10139_),
    .A2(_10609_),
    .ZN(_10610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15625_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_10211_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[20] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[20] ),
    .ZN(_10611_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15626_ (.A1(net2044),
    .A2(_10507_),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[20] ),
    .ZN(_10612_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15627_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(_10512_),
    .B(_10358_),
    .ZN(_10613_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15628_ (.A1(_10612_),
    .A2(_10613_),
    .Z(_10614_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15629_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1876] ),
    .ZN(_10615_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15630_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1908] ),
    .ZN(_10616_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15631_ (.A1(net1561),
    .A2(_10615_),
    .B1(_10616_),
    .B2(net1560),
    .ZN(_10617_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15632_ (.A1(net1562),
    .A2(_10617_),
    .ZN(_10618_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15633_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(net1556),
    .ZN(_10619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15634_ (.A1(\cs_registers_i.dscratch1_q[20] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .C1(net79),
    .C2(net1563),
    .ZN(_10620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15635_ (.A1(_10619_),
    .A2(_10620_),
    .Z(_10621_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15636_ (.A1(_10611_),
    .A2(_10614_),
    .A3(_10618_),
    .A4(_10621_),
    .Z(_10622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15637_ (.A1(_01281_),
    .A2(_10622_),
    .ZN(_10623_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15638_ (.A1(_10610_),
    .A2(_10623_),
    .Z(_10624_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15639_ (.A1(_10425_),
    .A2(_10624_),
    .ZN(_10625_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15640_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A2(_10526_),
    .A3(_10588_),
    .Z(_10626_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15641_ (.A1(net1518),
    .A2(_10626_),
    .ZN(_10627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15642_ (.I0(_10271_),
    .I1(_10626_),
    .S(net1518),
    .Z(_10628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15643_ (.I0(_10627_),
    .I1(_10628_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .Z(_10629_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15644_ (.A1(_10625_),
    .A2(_10629_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15645_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1680),
    .Z(_10630_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15646_ (.A1(_10139_),
    .A2(_10630_),
    .ZN(_10631_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15647_ (.A1(\cs_registers_i.csr_mepc_o[21] ),
    .A2(net1553),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[21] ),
    .ZN(_10632_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15648_ (.A1(\cs_registers_i.mtval_q[21] ),
    .A2(_10211_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[21] ),
    .ZN(_10633_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15649_ (.A1(_10632_),
    .A2(_10633_),
    .ZN(_10634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15650_ (.A1(net2043),
    .A2(_10507_),
    .B1(_10512_),
    .B2(\cs_registers_i.mie_q[5] ),
    .ZN(_10635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15651_ (.A1(\cs_registers_i.csr_mstatus_tw_o ),
    .A2(_10535_),
    .B(_10245_),
    .ZN(_10636_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15652_ (.A1(_10635_),
    .A2(_10636_),
    .ZN(_10637_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15653_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1877] ),
    .ZN(_10638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15654_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1909] ),
    .ZN(_10639_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15655_ (.A1(_10159_),
    .A2(_10638_),
    .B1(_10639_),
    .B2(net1560),
    .ZN(_10640_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15656_ (.A1(net1562),
    .A2(_10640_),
    .Z(_10641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15657_ (.A1(\cs_registers_i.dscratch0_q[21] ),
    .A2(net1556),
    .ZN(_10642_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15658_ (.A1(\cs_registers_i.dscratch1_q[21] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .C1(net80),
    .C2(net1563),
    .ZN(_10643_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15659_ (.A1(_10642_),
    .A2(_10643_),
    .ZN(_10644_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15660_ (.A1(_10634_),
    .A2(_10637_),
    .A3(_10641_),
    .A4(_10644_),
    .Z(_10645_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15661_ (.A1(net1680),
    .A2(_10645_),
    .Z(_10646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15662_ (.A1(_10631_),
    .A2(_10646_),
    .ZN(_10647_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15663_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A2(_10271_),
    .ZN(_10648_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15664_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ),
    .A3(_10497_),
    .A4(_10588_),
    .Z(_10649_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15665_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(net1518),
    .A3(_10649_),
    .Z(_10650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15666_ (.I0(_10648_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .S(_10650_),
    .Z(_10651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15667_ (.A1(_10425_),
    .A2(_10647_),
    .B(_10651_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15668_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1679),
    .Z(_10652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15669_ (.A1(net2042),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[22] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[22] ),
    .ZN(_10653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15670_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_10211_),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[22] ),
    .ZN(_10654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15671_ (.A1(\cs_registers_i.mie_q[6] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15672_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1878] ),
    .ZN(_10656_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15673_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1910] ),
    .ZN(_10657_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15674_ (.A1(net1561),
    .A2(_10656_),
    .B1(_10657_),
    .B2(net1560),
    .ZN(_10658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15675_ (.A1(\cs_registers_i.dscratch1_q[22] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .C1(net81),
    .C2(net1563),
    .ZN(_10659_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15676_ (.I(_10659_),
    .ZN(_10660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15677_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(net1556),
    .B1(_10658_),
    .B2(net1562),
    .C(_10660_),
    .ZN(_10661_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15678_ (.A1(_10653_),
    .A2(_10654_),
    .A3(_10655_),
    .A4(_10661_),
    .ZN(_10662_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15679_ (.A1(net1705),
    .A2(_10652_),
    .B1(_10662_),
    .B2(net1679),
    .ZN(_10663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15680_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .A2(_10271_),
    .ZN(_10664_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15681_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A3(net1518),
    .A4(_10626_),
    .ZN(_10665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15682_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .I1(_10664_),
    .S(_10665_),
    .Z(_10666_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15683_ (.A1(_10425_),
    .A2(_10663_),
    .B(_10666_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15684_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1678),
    .Z(_10667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15685_ (.A1(net2041),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[23] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[23] ),
    .ZN(_10668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15686_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_10211_),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_10669_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15687_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10670_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15688_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1879] ),
    .ZN(_10671_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15689_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1911] ),
    .ZN(_10672_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15690_ (.A1(net1561),
    .A2(_10671_),
    .B1(_10672_),
    .B2(net1560),
    .ZN(_10673_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15691_ (.A1(\cs_registers_i.dscratch1_q[23] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C1(net82),
    .C2(net1563),
    .ZN(_10674_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15692_ (.I(_10674_),
    .ZN(_10675_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15693_ (.A1(\cs_registers_i.dscratch0_q[23] ),
    .A2(net1556),
    .B1(_10673_),
    .B2(net1562),
    .C(_10675_),
    .ZN(_10676_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15694_ (.A1(_10668_),
    .A2(_10669_),
    .A3(_10670_),
    .A4(_10676_),
    .ZN(_10677_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15695_ (.A1(net1705),
    .A2(_10667_),
    .B1(_10677_),
    .B2(net1678),
    .ZN(_10678_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15696_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .A2(_10271_),
    .ZN(_10679_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15697_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ),
    .Z(_10680_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15698_ (.A1(net1518),
    .A2(_10649_),
    .A3(_10680_),
    .Z(_10681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15699_ (.I0(_10679_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .S(_10681_),
    .Z(_10682_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15700_ (.A1(_10425_),
    .A2(_10678_),
    .B(_10682_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15701_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1677),
    .Z(_10683_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15702_ (.A1(_10139_),
    .A2(_10683_),
    .ZN(_10684_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15703_ (.A1(net2040),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[24] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[24] ),
    .ZN(_10685_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15704_ (.A1(\cs_registers_i.mtval_q[24] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[24] ),
    .ZN(_10686_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15705_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10687_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15706_ (.A1(_10686_),
    .A2(_10687_),
    .Z(_10688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15707_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1880] ),
    .ZN(_10689_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15708_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1912] ),
    .ZN(_10690_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15709_ (.A1(net1561),
    .A2(_10689_),
    .B1(_10690_),
    .B2(net1560),
    .ZN(_10691_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15710_ (.A1(net1562),
    .A2(_10691_),
    .ZN(_10692_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15711_ (.A1(\cs_registers_i.dscratch0_q[24] ),
    .A2(net1556),
    .ZN(_10693_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15712_ (.A1(\cs_registers_i.dscratch1_q[24] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .C1(net83),
    .C2(net1563),
    .ZN(_10694_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15713_ (.A1(_10693_),
    .A2(_10694_),
    .Z(_10695_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15714_ (.A1(_10685_),
    .A2(_10688_),
    .A3(_10692_),
    .A4(_10695_),
    .ZN(_10696_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15715_ (.A1(net1677),
    .A2(_10696_),
    .Z(_10697_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15716_ (.A1(_10684_),
    .A2(_10697_),
    .ZN(_10698_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15717_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(_10266_),
    .ZN(_10699_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15718_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ),
    .A2(_10680_),
    .Z(_10700_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15719_ (.A1(net1518),
    .A2(_10626_),
    .A3(_10700_),
    .ZN(_10701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15720_ (.I0(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .I1(_10699_),
    .S(_10701_),
    .Z(_10702_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15721_ (.A1(_10502_),
    .A2(_10698_),
    .B(_10702_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15722_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A3(_10700_),
    .Z(_10703_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15723_ (.A1(_10649_),
    .A2(_10703_),
    .Z(_10704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15724_ (.I0(_00950_),
    .I1(_08009_),
    .S(_01312_),
    .Z(_10705_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15725_ (.A1(net2039),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[25] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[25] ),
    .ZN(_10706_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15726_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[25] ),
    .ZN(_10707_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15727_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15728_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1881] ),
    .ZN(_10709_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15729_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1913] ),
    .ZN(_10710_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15730_ (.A1(net1561),
    .A2(_10709_),
    .B1(_10710_),
    .B2(net1560),
    .ZN(_10711_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15731_ (.A1(\cs_registers_i.dscratch1_q[25] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .C1(net84),
    .C2(net1563),
    .ZN(_10712_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15732_ (.I(_10712_),
    .ZN(_10713_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15733_ (.A1(\cs_registers_i.dscratch0_q[25] ),
    .A2(net1556),
    .B1(_10711_),
    .B2(net1562),
    .C(_10713_),
    .ZN(_10714_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15734_ (.A1(_10706_),
    .A2(_10707_),
    .A3(_10708_),
    .A4(_10714_),
    .ZN(_10715_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15735_ (.A1(net1705),
    .A2(_10705_),
    .B1(_10715_),
    .B2(_01312_),
    .ZN(_10716_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15736_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ),
    .A2(net1518),
    .A3(_10649_),
    .A4(_10700_),
    .Z(_10717_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15737_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ),
    .A2(_10456_),
    .A3(_10717_),
    .ZN(_10718_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15738_ (.A1(net1518),
    .A2(_10704_),
    .B1(_10716_),
    .B2(_10456_),
    .C(_10718_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15739_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .ZN(_10719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15740_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01319_),
    .Z(_10720_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15741_ (.A1(_10139_),
    .A2(_10720_),
    .ZN(_10721_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15742_ (.A1(net136),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[26] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[26] ),
    .ZN(_10722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15743_ (.A1(\cs_registers_i.mtval_q[26] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[26] ),
    .ZN(_10723_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15744_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10724_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15745_ (.A1(_10723_),
    .A2(_10724_),
    .Z(_10725_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15746_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1882] ),
    .ZN(_10726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15747_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1914] ),
    .ZN(_10727_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15748_ (.A1(net1561),
    .A2(_10726_),
    .B1(_10727_),
    .B2(net1560),
    .ZN(_10728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15749_ (.A1(net1562),
    .A2(_10728_),
    .ZN(_10729_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15750_ (.A1(\cs_registers_i.dscratch0_q[26] ),
    .A2(net1556),
    .ZN(_10730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15751_ (.A1(\cs_registers_i.dscratch1_q[26] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[26] ),
    .C1(net85),
    .C2(net1563),
    .ZN(_10731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15752_ (.A1(_10730_),
    .A2(_10731_),
    .Z(_10732_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15753_ (.A1(_10722_),
    .A2(_10725_),
    .A3(_10729_),
    .A4(_10732_),
    .ZN(_10733_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15754_ (.A1(_01319_),
    .A2(_10733_),
    .Z(_10734_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15755_ (.A1(_10721_),
    .A2(_10734_),
    .Z(_10735_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1477 (.I(_05681_),
    .Z(net1476));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15757_ (.A1(_10626_),
    .A2(_10703_),
    .Z(_10737_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _15758_ (.A1(_10719_),
    .A2(_10737_),
    .ZN(_10738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15759_ (.A1(_10271_),
    .A2(_10735_),
    .B1(_10738_),
    .B2(net1518),
    .ZN(_10739_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15760_ (.A1(_10719_),
    .A2(_10267_),
    .B(_10739_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15761_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A2(_10271_),
    .ZN(_10740_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15762_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(net1518),
    .A3(_10704_),
    .Z(_10741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15763_ (.I0(_10740_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .S(_10741_),
    .Z(_10742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15764_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01326_),
    .Z(_10743_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15765_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(_10211_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[27] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[27] ),
    .ZN(_10744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15766_ (.A1(net2049),
    .A2(_10507_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[27] ),
    .ZN(_10745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15767_ (.A1(\cs_registers_i.mie_q[11] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10746_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15768_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1883] ),
    .ZN(_10747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15769_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1915] ),
    .ZN(_10748_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15770_ (.A1(net1561),
    .A2(_10747_),
    .B1(_10748_),
    .B2(net1560),
    .ZN(_10749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15771_ (.A1(\cs_registers_i.dscratch1_q[27] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .C1(net86),
    .C2(net1563),
    .ZN(_10750_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15772_ (.I(_10750_),
    .ZN(_10751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15773_ (.A1(\cs_registers_i.dscratch0_q[27] ),
    .A2(net1556),
    .B1(_10749_),
    .B2(net1562),
    .C(_10751_),
    .ZN(_10752_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15774_ (.A1(_10744_),
    .A2(_10745_),
    .A3(_10746_),
    .A4(_10752_),
    .Z(_10753_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15775_ (.A1(_10139_),
    .A2(_10743_),
    .B1(_10753_),
    .B2(_01330_),
    .ZN(_10754_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1475 (.I(_05685_),
    .Z(net1474));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15777_ (.A1(_10502_),
    .A2(net1517),
    .ZN(_10756_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15778_ (.A1(_10742_),
    .A2(_10756_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15779_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .Z(_10757_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15780_ (.A1(_10376_),
    .A2(_10737_),
    .A3(_10757_),
    .ZN(_10758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15781_ (.I0(_10758_),
    .I1(_10450_),
    .S(net1532),
    .Z(_10759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15782_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(_10759_),
    .ZN(_10760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15783_ (.A1(net2048),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[28] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[28] ),
    .ZN(_10761_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15784_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(_10211_),
    .B1(net1558),
    .B2(\cs_registers_i.csr_mtvec_o[28] ),
    .ZN(_10762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15785_ (.A1(\cs_registers_i.mie_q[12] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15786_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1884] ),
    .ZN(_10764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15787_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1916] ),
    .ZN(_10765_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15788_ (.A1(net1561),
    .A2(_10764_),
    .B1(_10765_),
    .B2(net1560),
    .ZN(_10766_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15789_ (.A1(\cs_registers_i.dscratch1_q[28] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .C1(net87),
    .C2(net1563),
    .ZN(_10767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15790_ (.I(_10767_),
    .ZN(_10768_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15791_ (.A1(\cs_registers_i.dscratch0_q[28] ),
    .A2(net1556),
    .B1(_10766_),
    .B2(net1562),
    .C(_10768_),
    .ZN(_10769_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15792_ (.A1(_10761_),
    .A2(_10762_),
    .A3(_10763_),
    .A4(_10769_),
    .Z(_10770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15793_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1676),
    .Z(_10771_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15794_ (.A1(net1705),
    .A2(_10771_),
    .ZN(_10772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15795_ (.A1(_01337_),
    .A2(_10770_),
    .B(_10772_),
    .ZN(_10773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1473 (.I(_05693_),
    .Z(net1472));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15797_ (.A1(_10271_),
    .A2(net1516),
    .ZN(_10775_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15798_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(net1532),
    .A3(_10758_),
    .Z(_10776_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15799_ (.A1(_10760_),
    .A2(_10775_),
    .A3(_10776_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15800_ (.I0(_00950_),
    .I1(_08009_),
    .S(net1675),
    .Z(_10777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15801_ (.A1(net139),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[29] ),
    .C1(net1553),
    .C2(\cs_registers_i.csr_mepc_o[29] ),
    .ZN(_10778_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15802_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_10211_),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[29] ),
    .ZN(_10779_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15803_ (.A1(\cs_registers_i.mie_q[13] ),
    .A2(_10512_),
    .B(_10245_),
    .ZN(_10780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15804_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1885] ),
    .ZN(_10781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15805_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1917] ),
    .ZN(_10782_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15806_ (.A1(net1561),
    .A2(_10781_),
    .B1(_10782_),
    .B2(net1560),
    .ZN(_10783_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15807_ (.A1(\cs_registers_i.dscratch1_q[29] ),
    .A2(net1559),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .C1(net88),
    .C2(net1563),
    .ZN(_10784_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15808_ (.I(_10784_),
    .ZN(_10785_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15809_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(net1556),
    .B1(_10783_),
    .B2(net1562),
    .C(_10785_),
    .ZN(_10786_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15810_ (.A1(_10778_),
    .A2(_10779_),
    .A3(_10780_),
    .A4(_10786_),
    .ZN(_10787_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15811_ (.A1(net1705),
    .A2(_10777_),
    .B1(_10787_),
    .B2(net1675),
    .ZN(_10788_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15812_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .A2(_10271_),
    .ZN(_10789_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15813_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A2(net1518),
    .A3(_10704_),
    .A4(_10757_),
    .Z(_10790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15814_ (.I0(_10789_),
    .I1(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .S(_10790_),
    .Z(_10791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15815_ (.A1(_10425_),
    .A2(_10788_),
    .B(_10791_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15816_ (.I(_10258_),
    .ZN(_10792_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15817_ (.A1(_10175_),
    .A2(net1562),
    .ZN(_10793_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _15818_ (.A1(_10423_),
    .A2(_10421_),
    .A3(_10793_),
    .ZN(_10794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15819_ (.A1(_10376_),
    .A2(_01369_),
    .B(net1532),
    .ZN(_10795_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15820_ (.A1(net1530),
    .A2(_10795_),
    .Z(_10796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15821_ (.A1(_01369_),
    .A2(net1518),
    .Z(_10797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15822_ (.I0(_10796_),
    .I1(_10797_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .Z(_10798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15823_ (.A1(_10792_),
    .A2(_10425_),
    .B(_10798_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15824_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .ZN(_10799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15825_ (.A1(\cs_registers_i.mtval_q[30] ),
    .A2(net1555),
    .B1(net1557),
    .B2(\cs_registers_i.csr_mtvec_o[30] ),
    .C1(_10512_),
    .C2(\cs_registers_i.mie_q[14] ),
    .ZN(_10800_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15826_ (.A1(net140),
    .A2(_10507_),
    .B1(net1554),
    .B2(\cs_registers_i.mscratch_q[30] ),
    .ZN(_10801_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15827_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(net1553),
    .B(_10358_),
    .ZN(_10802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15828_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1886] ),
    .ZN(_10803_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15829_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(net1609),
    .B1(net1564),
    .B2(\cs_registers_i.mhpmcounter[1918] ),
    .ZN(_10804_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15830_ (.A1(_10159_),
    .A2(_10803_),
    .B1(_10804_),
    .B2(net1560),
    .ZN(_10805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15831_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_10188_),
    .B(_10201_),
    .ZN(_10806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15832_ (.A1(net90),
    .A2(net1563),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .ZN(_10807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15833_ (.A1(_10806_),
    .A2(_10807_),
    .ZN(_10808_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15834_ (.A1(\cs_registers_i.dscratch0_q[30] ),
    .A2(net1556),
    .B1(_10805_),
    .B2(net1562),
    .C(_10808_),
    .ZN(_10809_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15835_ (.A1(_10800_),
    .A2(_10801_),
    .A3(_10802_),
    .A4(_10809_),
    .Z(_10810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15836_ (.I0(_00950_),
    .I1(_08009_),
    .S(_01347_),
    .Z(_10811_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15837_ (.A1(net1705),
    .A2(_10811_),
    .ZN(_10812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15838_ (.A1(_01351_),
    .A2(_10810_),
    .B(_10812_),
    .ZN(_10813_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15839_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ),
    .Z(_10814_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15840_ (.A1(_10737_),
    .A2(_10814_),
    .Z(_10815_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _15841_ (.A1(_10799_),
    .A2(_10815_),
    .ZN(_10816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15842_ (.A1(_10271_),
    .A2(_10813_),
    .B1(_10816_),
    .B2(net1518),
    .ZN(_10817_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15843_ (.A1(_10799_),
    .A2(_10267_),
    .B(_10817_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15844_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .ZN(_10818_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15845_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ),
    .A2(_10814_),
    .Z(_10819_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15846_ (.A1(_10704_),
    .A2(_10819_),
    .Z(_10820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15847_ (.I0(_10271_),
    .I1(_10820_),
    .S(net1518),
    .Z(_10821_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15848_ (.A1(_10818_),
    .A2(_10820_),
    .Z(_10822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15849_ (.A1(\cs_registers_i.mcause_q[5] ),
    .A2(_10214_),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[31] ),
    .ZN(_10823_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15850_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(net1555),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[31] ),
    .ZN(_10824_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15851_ (.A1(_10823_),
    .A2(_10824_),
    .ZN(_10825_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15852_ (.A1(_09628_),
    .A2(_10417_),
    .Z(_10826_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15853_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_10826_),
    .A3(_10218_),
    .Z(_10827_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15854_ (.A1(_10180_),
    .A2(_10415_),
    .A3(_09603_),
    .A4(_10181_),
    .Z(_10828_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15855_ (.A1(net91),
    .A2(_10828_),
    .Z(_10829_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15856_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_10826_),
    .A3(_10187_),
    .Z(_10830_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15857_ (.A1(_10827_),
    .A2(_10829_),
    .A3(_10830_),
    .Z(_10831_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _15858_ (.I(\cs_registers_i.dscratch0_q[31] ),
    .ZN(_10832_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15859_ (.A1(_10146_),
    .A2(_10149_),
    .Z(_10833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15860_ (.A1(_10826_),
    .A2(_10833_),
    .ZN(_10834_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15861_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_10197_),
    .ZN(_10835_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15862_ (.A1(_10177_),
    .A2(_10409_),
    .ZN(_10836_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _15863_ (.A1(_10832_),
    .A2(_10834_),
    .B(_10835_),
    .C(_10836_),
    .ZN(_10837_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15864_ (.A1(_09575_),
    .A2(_10155_),
    .A3(_10407_),
    .ZN(_10838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15865_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1887] ),
    .ZN(_10839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15866_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(net1609),
    .B1(net1565),
    .B2(\cs_registers_i.mhpmcounter[1919] ),
    .ZN(_10840_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15867_ (.A1(_10838_),
    .A2(_10839_),
    .B1(_10840_),
    .B2(_10423_),
    .ZN(_10841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15868_ (.A1(net1562),
    .A2(_10841_),
    .Z(_10842_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _15869_ (.A1(_10825_),
    .A2(_10831_),
    .A3(_10837_),
    .A4(_10842_),
    .ZN(_10843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15870_ (.I0(_08008_),
    .I1(_10141_),
    .S(_09470_),
    .Z(_10844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15871_ (.A1(_10139_),
    .A2(_10844_),
    .Z(_10845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15872_ (.A1(_09470_),
    .A2(_10843_),
    .B(_10845_),
    .ZN(_10846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15873_ (.A1(net1518),
    .A2(_10822_),
    .B1(_10846_),
    .B2(_10425_),
    .ZN(_10847_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15874_ (.A1(_10818_),
    .A2(_10821_),
    .B(_10847_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1464 (.I(_05715_),
    .Z(net1463));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15876_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A2(_10737_),
    .A3(_10819_),
    .Z(_10849_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _15877_ (.A1(_10162_),
    .A2(_10370_),
    .A3(_10371_),
    .A4(_10793_),
    .ZN(_10850_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15878_ (.A1(_10376_),
    .A2(_10850_),
    .Z(_10851_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15879_ (.A1(_10849_),
    .A2(_10851_),
    .ZN(_10852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15880_ (.I0(_10849_),
    .I1(_10852_),
    .S(_10168_),
    .Z(_10853_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1462 (.I(_05719_),
    .Z(net1461));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _15882_ (.A1(net1518),
    .A2(_10850_),
    .ZN(_10855_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1461 (.I(_05723_),
    .Z(net1460));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15884_ (.A1(_10225_),
    .A2(net1530),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .ZN(_10857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15885_ (.A1(net1532),
    .A2(_10853_),
    .B(_10857_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15886_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .A3(_10820_),
    .ZN(_10858_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _15887_ (.A1(_10376_),
    .A2(_10850_),
    .ZN(_10859_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1460 (.I(net185),
    .Z(net1459));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15889_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(net1509),
    .A3(_10858_),
    .ZN(_10861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15890_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(_10858_),
    .B(_10861_),
    .ZN(_10862_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1459 (.I(net184),
    .Z(net1458));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15892_ (.A1(net1530),
    .A2(_10607_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .ZN(_10864_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15893_ (.A1(net1532),
    .A2(_10862_),
    .B(_10864_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _15894_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A3(_10849_),
    .ZN(_10865_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15895_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(net1509),
    .A3(_10865_),
    .ZN(_10866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15896_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A2(_10865_),
    .B(_10866_),
    .ZN(_10867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15897_ (.A1(_10258_),
    .A2(net1530),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .ZN(_10868_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15898_ (.A1(net1532),
    .A2(_10867_),
    .B(_10868_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15899_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .A4(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ),
    .Z(_10869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15900_ (.A1(_10819_),
    .A2(_10869_),
    .Z(_10870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15901_ (.A1(_10704_),
    .A2(_10870_),
    .Z(_10871_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15902_ (.A1(_10851_),
    .A2(_10871_),
    .ZN(_10872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15903_ (.I0(_10872_),
    .I1(_10871_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .Z(_10873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15904_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2103),
    .Z(_10874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15905_ (.A1(_10139_),
    .A2(_10874_),
    .ZN(_10875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15906_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(net1555),
    .B1(_10512_),
    .B2(\cs_registers_i.mie_q[17] ),
    .ZN(_10876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15907_ (.A1(net151),
    .A2(_10507_),
    .B1(_10214_),
    .B2(\cs_registers_i.mcause_q[3] ),
    .ZN(_10877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15908_ (.A1(_10876_),
    .A2(_10877_),
    .ZN(_10878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15909_ (.A1(\cs_registers_i.csr_mepc_o[3] ),
    .A2(net1553),
    .B1(_10535_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .ZN(_10879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15910_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_10216_),
    .B(_10245_),
    .ZN(_10880_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15911_ (.A1(_10879_),
    .A2(_10880_),
    .ZN(_10881_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15912_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1859] ),
    .ZN(_10882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15913_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1891] ),
    .ZN(_10883_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15914_ (.A1(_10159_),
    .A2(_10882_),
    .B1(_10883_),
    .B2(_10162_),
    .ZN(_10884_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15915_ (.A1(net1562),
    .A2(_10884_),
    .Z(_10885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15916_ (.A1(\cs_registers_i.dscratch0_q[3] ),
    .A2(net1556),
    .ZN(_10886_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15917_ (.A1(\cs_registers_i.dscratch1_q[3] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[3] ),
    .C1(net92),
    .C2(net1563),
    .ZN(_10887_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15918_ (.A1(_10886_),
    .A2(_10887_),
    .ZN(_10888_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _15919_ (.A1(_10878_),
    .A2(_10881_),
    .A3(_10885_),
    .A4(_10888_),
    .Z(_10889_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15920_ (.A1(net2103),
    .A2(_10889_),
    .Z(_10890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15921_ (.A1(_10875_),
    .A2(_10890_),
    .Z(_10891_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15922_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(net1510),
    .B1(_10891_),
    .B2(net1530),
    .ZN(_10892_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15923_ (.A1(net1532),
    .A2(_10873_),
    .B(_10892_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15924_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ),
    .ZN(_10893_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15925_ (.A1(_10865_),
    .A2(_10893_),
    .Z(_10894_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15926_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(net1509),
    .A3(_10894_),
    .ZN(_10895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15927_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(_10894_),
    .B(_10895_),
    .ZN(_10896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15928_ (.I0(_10141_),
    .I1(_08008_),
    .S(_01165_),
    .Z(_10897_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15929_ (.A1(_10139_),
    .A2(_10897_),
    .ZN(_10898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15930_ (.A1(\cs_registers_i.mtval_q[4] ),
    .A2(_10211_),
    .B1(_10214_),
    .B2(\cs_registers_i.mcause_q[4] ),
    .C1(_10216_),
    .C2(\cs_registers_i.mscratch_q[4] ),
    .ZN(_10899_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15931_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(_10826_),
    .A3(_10218_),
    .Z(_10900_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15932_ (.A1(\cs_registers_i.dscratch1_q[4] ),
    .A2(_10826_),
    .A3(_10187_),
    .Z(_10901_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _15933_ (.A1(net93),
    .A2(_10828_),
    .B(_10900_),
    .C(_10901_),
    .ZN(_10902_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15934_ (.A1(\cs_registers_i.dscratch0_q[4] ),
    .A2(_10826_),
    .A3(_10833_),
    .Z(_10903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _15935_ (.A1(_10177_),
    .A2(_10409_),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .C(_10903_),
    .ZN(_10904_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15936_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1860] ),
    .ZN(_10905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15937_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1892] ),
    .ZN(_10906_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15938_ (.A1(_10838_),
    .A2(_10905_),
    .B1(_10906_),
    .B2(_10423_),
    .ZN(_10907_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15939_ (.A1(net1562),
    .A2(_10907_),
    .ZN(_10908_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15940_ (.A1(_10899_),
    .A2(_10902_),
    .A3(_10904_),
    .A4(_10908_),
    .ZN(_10909_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15941_ (.A1(_01165_),
    .A2(_10909_),
    .Z(_10910_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15942_ (.A1(_10898_),
    .A2(_10910_),
    .Z(_10911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15943_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .A2(net1510),
    .B1(_10911_),
    .B2(net1530),
    .ZN(_10912_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15944_ (.A1(net1532),
    .A2(_10896_),
    .B(_10912_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15945_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ),
    .Z(_10913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15946_ (.A1(_10871_),
    .A2(_10913_),
    .ZN(_10914_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _15947_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(net1509),
    .A3(_10914_),
    .ZN(_10915_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15948_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_10914_),
    .B(_10915_),
    .ZN(_10916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15949_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1692),
    .Z(_10917_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15950_ (.A1(_09602_),
    .A2(_09613_),
    .A3(_09614_),
    .Z(_10918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15951_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1861] ),
    .ZN(_10919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15952_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1893] ),
    .ZN(_10920_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _15953_ (.A1(_09612_),
    .A2(_09613_),
    .A3(_09614_),
    .Z(_10921_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15954_ (.A1(_10918_),
    .A2(_10919_),
    .B1(_10920_),
    .B2(_10921_),
    .ZN(_10922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15955_ (.A1(_09569_),
    .A2(_09579_),
    .A3(_09582_),
    .Z(_10923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15956_ (.A1(\cs_registers_i.csr_mepc_o[5] ),
    .A2(_10923_),
    .B(_10178_),
    .ZN(_10924_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15957_ (.A1(_09558_),
    .A2(_09582_),
    .A3(net1608),
    .Z(_10925_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15958_ (.A1(net1612),
    .A2(net1586),
    .Z(_10926_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15959_ (.A1(_10926_),
    .A2(_09579_),
    .A3(_09582_),
    .Z(_10927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15960_ (.A1(\cs_registers_i.mscratch_q[5] ),
    .A2(_10925_),
    .B1(_10927_),
    .B2(\cs_registers_i.mtval_q[5] ),
    .ZN(_10928_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15961_ (.A1(net1696),
    .A2(_09543_),
    .A3(_09552_),
    .A4(_09601_),
    .Z(_10929_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15962_ (.A1(_10929_),
    .A2(_10926_),
    .A3(_09579_),
    .Z(_10930_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15963_ (.A1(net1610),
    .A2(_09601_),
    .Z(_10931_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15964_ (.A1(_09543_),
    .A2(_09603_),
    .A3(_09581_),
    .A4(_10931_),
    .Z(_10932_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15965_ (.A1(\cs_registers_i.dscratch1_q[5] ),
    .A2(_10930_),
    .B1(_10932_),
    .B2(net94),
    .ZN(_10933_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15966_ (.A1(net1586),
    .A2(_10329_),
    .Z(_10934_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15967_ (.A1(_09558_),
    .A2(_10929_),
    .A3(_10934_),
    .Z(_10935_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _15968_ (.A1(_10929_),
    .A2(_09569_),
    .A3(_09579_),
    .Z(_10936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15969_ (.A1(\cs_registers_i.dscratch0_q[5] ),
    .A2(_10935_),
    .B1(_10936_),
    .B2(\cs_registers_i.csr_depc_o[5] ),
    .ZN(_10937_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15970_ (.A1(_10924_),
    .A2(_10928_),
    .A3(_10933_),
    .A4(_10937_),
    .ZN(_10938_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15971_ (.A1(_10261_),
    .A2(_10922_),
    .B(_10938_),
    .ZN(_10939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15972_ (.A1(_10139_),
    .A2(_10917_),
    .B1(_10939_),
    .B2(_01176_),
    .ZN(_10940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15973_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(net1510),
    .B1(_10940_),
    .B2(net1530),
    .ZN(_10941_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15974_ (.A1(net1532),
    .A2(_10916_),
    .B(_10941_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1458 (.I(net157),
    .Z(net1457));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _15976_ (.I0(_10141_),
    .I1(_08008_),
    .S(net1691),
    .Z(_10943_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15977_ (.A1(_10139_),
    .A2(_10943_),
    .ZN(_10944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15978_ (.A1(\cs_registers_i.mtval_q[6] ),
    .A2(_10211_),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[6] ),
    .ZN(_10945_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _15979_ (.A1(\cs_registers_i.mscratch_q[6] ),
    .A2(_10216_),
    .B(_10245_),
    .ZN(_10946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15980_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1862] ),
    .ZN(_10947_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15981_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(net1608),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1894] ),
    .ZN(_10948_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _15982_ (.A1(_10159_),
    .A2(_10947_),
    .B1(_10948_),
    .B2(_10162_),
    .ZN(_10949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15983_ (.A1(net1562),
    .A2(_10949_),
    .ZN(_10950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _15984_ (.A1(\cs_registers_i.dscratch1_q[6] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[6] ),
    .C1(net95),
    .C2(net1563),
    .ZN(_10951_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15985_ (.A1(\cs_registers_i.dcsr_q[6] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[6] ),
    .ZN(_10952_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15986_ (.A1(_10951_),
    .A2(_10952_),
    .Z(_10953_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _15987_ (.A1(_10945_),
    .A2(_10946_),
    .A3(_10950_),
    .A4(_10953_),
    .ZN(_10954_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _15988_ (.A1(net1691),
    .A2(_10954_),
    .Z(_10955_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _15989_ (.A1(_10944_),
    .A2(_10955_),
    .Z(_10956_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1463 (.I(_05719_),
    .Z(net1462));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _15991_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(net1510),
    .B1(_10956_),
    .B2(net1530),
    .ZN(_10958_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1457 (.I(net160),
    .Z(net1456));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1456 (.I(_08838_),
    .Z(net1455));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _15994_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_10703_),
    .A3(_10870_),
    .A4(_10913_),
    .Z(_10961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15995_ (.A1(_10626_),
    .A2(_10961_),
    .ZN(_10962_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15996_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(_10962_),
    .ZN(_10963_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _15997_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A2(net1509),
    .A3(_10962_),
    .B(_10963_),
    .ZN(_10964_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15998_ (.A1(net1511),
    .A2(_10964_),
    .ZN(_10965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _15999_ (.A1(_10958_),
    .A2(_10965_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16000_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .A3(_10871_),
    .A4(_10913_),
    .ZN(_10966_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16001_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(net1509),
    .A3(_10966_),
    .ZN(_10967_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16002_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(_10966_),
    .B(_10967_),
    .ZN(_10968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16003_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2116),
    .Z(_10969_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16004_ (.A1(_10139_),
    .A2(_10969_),
    .ZN(_10970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16005_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(net1553),
    .B1(_10535_),
    .B2(\cs_registers_i.mstatus_q[4] ),
    .C1(_10512_),
    .C2(\cs_registers_i.mie_q[16] ),
    .ZN(_10971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16006_ (.A1(\cs_registers_i.mtval_q[7] ),
    .A2(net1555),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[7] ),
    .ZN(_10972_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16007_ (.A1(net152),
    .A2(_10507_),
    .B(_10245_),
    .ZN(_10973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16008_ (.A1(_10972_),
    .A2(_10973_),
    .Z(_10974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16009_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1863] ),
    .ZN(_10975_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16010_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1895] ),
    .ZN(_10976_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16011_ (.A1(_10159_),
    .A2(_10975_),
    .B1(_10976_),
    .B2(net1560),
    .ZN(_10977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16012_ (.A1(net1562),
    .A2(_10977_),
    .ZN(_10978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16013_ (.A1(\cs_registers_i.dscratch1_q[7] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .C1(net96),
    .C2(net1563),
    .ZN(_10979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16014_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[7] ),
    .ZN(_10980_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16015_ (.A1(_10979_),
    .A2(_10980_),
    .Z(_10981_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16016_ (.A1(_10971_),
    .A2(_10974_),
    .A3(_10978_),
    .A4(_10981_),
    .ZN(_10982_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16017_ (.A1(net2116),
    .A2(_10982_),
    .Z(_10983_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16018_ (.A1(_10970_),
    .A2(_10983_),
    .Z(_10984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16019_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(net1510),
    .B1(_10984_),
    .B2(net1530),
    .ZN(_10985_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16020_ (.A1(net1532),
    .A2(_10968_),
    .B(_10985_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16021_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A2(_10309_),
    .Z(_10986_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _16022_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(_10986_),
    .Z(_10987_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16023_ (.A1(_10271_),
    .A2(_10891_),
    .B1(_10987_),
    .B2(net1518),
    .ZN(_10988_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16024_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(_10306_),
    .ZN(_10989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16025_ (.A1(_10988_),
    .A2(_10989_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16026_ (.A1(_10626_),
    .A2(_10961_),
    .Z(_10990_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16027_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ),
    .Z(_10991_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16028_ (.A1(_10990_),
    .A2(_10991_),
    .ZN(_10992_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16029_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(_10992_),
    .ZN(_10993_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16030_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(net1509),
    .A3(_10992_),
    .Z(_10994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16031_ (.A1(_10993_),
    .A2(_10994_),
    .Z(_10995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16032_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2072),
    .Z(_10996_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16033_ (.A1(_10139_),
    .A2(_10996_),
    .Z(_10997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16034_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(net1555),
    .B1(_10216_),
    .B2(\cs_registers_i.mscratch_q[8] ),
    .C1(_10197_),
    .C2(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_10998_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16035_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1864] ),
    .ZN(_10999_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16036_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1896] ),
    .ZN(_11000_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16037_ (.A1(_10159_),
    .A2(_10999_),
    .B1(_11000_),
    .B2(net1560),
    .ZN(_11001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16038_ (.A1(net1562),
    .A2(_11001_),
    .ZN(_11002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16039_ (.A1(\cs_registers_i.dscratch1_q[8] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .C1(net97),
    .C2(net1563),
    .ZN(_11003_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16040_ (.A1(\cs_registers_i.dcsr_q[8] ),
    .A2(_10201_),
    .B1(net1556),
    .B2(\cs_registers_i.dscratch0_q[8] ),
    .ZN(_11004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16041_ (.A1(_11003_),
    .A2(_11004_),
    .Z(_11005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16042_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(net1553),
    .B(_10358_),
    .ZN(_11006_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16043_ (.A1(_10998_),
    .A2(_11002_),
    .A3(_11005_),
    .A4(_11006_),
    .Z(_11007_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16044_ (.A1(_01197_),
    .A2(_11007_),
    .Z(_11008_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16045_ (.A1(_10997_),
    .A2(_11008_),
    .ZN(_11009_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16046_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(net1510),
    .B1(_11009_),
    .B2(net1530),
    .ZN(_11010_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16047_ (.A1(net1532),
    .A2(_10995_),
    .B(_11010_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16048_ (.I0(_10141_),
    .I1(_08008_),
    .S(net2097),
    .Z(_11011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16049_ (.A1(_10139_),
    .A2(_11011_),
    .ZN(_11012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16050_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(net1555),
    .B1(net1553),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .C1(_10197_),
    .C2(\cs_registers_i.csr_mtvec_o[9] ),
    .ZN(_11013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16051_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1865] ),
    .ZN(_11014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16052_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(net1609),
    .B1(_10149_),
    .B2(\cs_registers_i.mhpmcounter[1897] ),
    .ZN(_11015_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16053_ (.A1(_10159_),
    .A2(_11014_),
    .B1(_11015_),
    .B2(net1560),
    .ZN(_11016_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16054_ (.A1(net1562),
    .A2(_11016_),
    .ZN(_11017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16055_ (.A1(\cs_registers_i.dscratch0_q[9] ),
    .A2(net1556),
    .ZN(_11018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _16056_ (.A1(\cs_registers_i.dscratch1_q[9] ),
    .A2(_10188_),
    .B1(net1552),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .C1(net98),
    .C2(net1563),
    .ZN(_11019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16057_ (.A1(\cs_registers_i.mscratch_q[9] ),
    .A2(_10216_),
    .B(_10245_),
    .ZN(_11020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16058_ (.A1(_11018_),
    .A2(_11019_),
    .A3(_11020_),
    .Z(_11021_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16059_ (.A1(_11013_),
    .A2(_11017_),
    .A3(_11021_),
    .ZN(_11022_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16060_ (.A1(net2097),
    .A2(_11022_),
    .Z(_11023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16061_ (.A1(_11012_),
    .A2(_11023_),
    .Z(_11024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16062_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(net1510),
    .B1(_11024_),
    .B2(net1530),
    .ZN(_11025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16063_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(_10991_),
    .Z(_11026_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16064_ (.A1(_10649_),
    .A2(_10961_),
    .A3(_11026_),
    .ZN(_11027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16065_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(_11027_),
    .ZN(_11028_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16066_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(net1509),
    .A3(_11027_),
    .B(_11028_),
    .ZN(_11029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16067_ (.A1(net1511),
    .A2(_11029_),
    .ZN(_11030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16068_ (.A1(_11025_),
    .A2(_11030_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16069_ (.A1(_10280_),
    .A2(_10282_),
    .A3(_10283_),
    .A4(_10297_),
    .ZN(_11031_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16070_ (.A1(net1705),
    .A2(_10279_),
    .ZN(_11032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16071_ (.A1(_01211_),
    .A2(_11031_),
    .B(_11032_),
    .ZN(_11033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16072_ (.A1(_11033_),
    .A2(net1530),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .ZN(_11034_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16073_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A3(_10990_),
    .A4(_10991_),
    .ZN(_11035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16074_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(_11035_),
    .ZN(_11036_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16075_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A2(net1509),
    .A3(_11035_),
    .B(_11036_),
    .ZN(_11037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16076_ (.A1(net1511),
    .A2(_11037_),
    .ZN(_11038_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16077_ (.A1(_11034_),
    .A2(_11038_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16078_ (.A1(_10348_),
    .A2(net1530),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .ZN(_11039_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16079_ (.A1(_10649_),
    .A2(_10961_),
    .A3(_11026_),
    .Z(_11040_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16080_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A3(_11040_),
    .ZN(_11041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16081_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(_11041_),
    .ZN(_11042_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16082_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(net1509),
    .A3(_11041_),
    .B(_11042_),
    .ZN(_11043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16083_ (.A1(net1511),
    .A2(_11043_),
    .ZN(_11044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16084_ (.A1(_11039_),
    .A2(_11044_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16085_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A3(_10990_),
    .A4(_10991_),
    .Z(_11045_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16086_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A3(_11045_),
    .ZN(_11046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16087_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_11046_),
    .ZN(_11047_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16088_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(net1509),
    .A3(_11046_),
    .Z(_11048_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16089_ (.A1(_11047_),
    .A2(_11048_),
    .Z(_11049_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16090_ (.A1(_10386_),
    .A2(_10393_),
    .A3(_10400_),
    .A4(_10402_),
    .ZN(_11050_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16091_ (.A1(net1705),
    .A2(_10380_),
    .ZN(_11051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16092_ (.A1(_01222_),
    .A2(_11050_),
    .B(_11051_),
    .ZN(_11052_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16093_ (.A1(net1530),
    .A2(_11052_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .ZN(_11053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16094_ (.A1(net1532),
    .A2(_11049_),
    .B(_11053_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16095_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A4(_11040_),
    .Z(_11054_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16096_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(_11054_),
    .ZN(_11055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16097_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(_11055_),
    .ZN(_11056_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16098_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .A2(net1509),
    .A3(_11055_),
    .Z(_11057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16099_ (.A1(_11056_),
    .A2(_11057_),
    .Z(_11058_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16100_ (.A1(_10431_),
    .A2(_10447_),
    .ZN(_11059_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1465 (.I(_05715_),
    .Z(net1464));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16102_ (.A1(net1530),
    .A2(_11059_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .ZN(_11061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16103_ (.A1(net1532),
    .A2(_11058_),
    .B(_11061_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16104_ (.A1(_10459_),
    .A2(_10470_),
    .ZN(_11062_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16105_ (.A1(net1705),
    .A2(_10457_),
    .ZN(_11063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16106_ (.A1(_01239_),
    .A2(_11062_),
    .B(_11063_),
    .ZN(_11064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16107_ (.A1(net1530),
    .A2(_11064_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .ZN(_11065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16108_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ),
    .Z(_11066_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16109_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A3(_11045_),
    .A4(_11066_),
    .Z(_11067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16110_ (.I(_11067_),
    .ZN(_11068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16111_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_11068_),
    .ZN(_11069_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16112_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(net1509),
    .A3(_11068_),
    .B(_11069_),
    .ZN(_11070_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16113_ (.A1(net1511),
    .A2(_11070_),
    .ZN(_11071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16114_ (.A1(_11065_),
    .A2(_11071_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1467 (.I(_05711_),
    .Z(net1466));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16116_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(_11054_),
    .A3(_11066_),
    .ZN(_11073_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16117_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(net1509),
    .A3(_11073_),
    .ZN(_11074_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16118_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(_11073_),
    .B(_11074_),
    .ZN(_11075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16119_ (.A1(net1530),
    .A2(net1531),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .ZN(_11076_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16120_ (.A1(net1532),
    .A2(_11075_),
    .B(_11076_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16121_ (.A1(_10506_),
    .A2(_10524_),
    .Z(_11077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16122_ (.A1(net1530),
    .A2(_11077_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .ZN(_11078_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16123_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A3(_11067_),
    .ZN(_11079_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16124_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(_11079_),
    .ZN(_11080_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16125_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(net1509),
    .A3(_11079_),
    .B(_11080_),
    .ZN(_11081_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16126_ (.A1(net1511),
    .A2(_11081_),
    .ZN(_11082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16127_ (.A1(_11078_),
    .A2(_11082_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16128_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .ZN(_11083_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16129_ (.A1(_11073_),
    .A2(_11083_),
    .Z(_11084_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16130_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(net1509),
    .A3(_11084_),
    .ZN(_11085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16131_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(_11084_),
    .B(_11085_),
    .ZN(_11086_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16132_ (.A1(_10533_),
    .A2(_10537_),
    .A3(_10541_),
    .A4(_10544_),
    .Z(_11087_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16133_ (.A1(net1705),
    .A2(_10530_),
    .ZN(_11088_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16134_ (.A1(_01260_),
    .A2(_11087_),
    .B(_11088_),
    .ZN(_11089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16135_ (.A1(net1530),
    .A2(_11089_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .ZN(_11090_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16136_ (.A1(net1532),
    .A2(_11086_),
    .B(_11090_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16137_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A3(_01369_),
    .A4(net1518),
    .Z(_11091_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16138_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A2(_10456_),
    .A3(_11091_),
    .Z(_11092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16139_ (.A1(_10898_),
    .A2(_10910_),
    .ZN(_11093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16140_ (.A1(_10456_),
    .A2(_11093_),
    .B1(_11091_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .ZN(_11094_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16141_ (.A1(_11092_),
    .A2(_11094_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16142_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ),
    .A2(_10703_),
    .A3(_10870_),
    .A4(_10913_),
    .Z(_11095_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16143_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ),
    .A2(_10626_),
    .A3(_11095_),
    .A4(_11026_),
    .Z(_11096_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16144_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ),
    .A3(_11096_),
    .A4(_11066_),
    .Z(_11097_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16145_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .Z(_11098_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16146_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ),
    .A3(_11097_),
    .A4(_11098_),
    .Z(_11099_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16147_ (.I(_11099_),
    .ZN(_11100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16148_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(_11100_),
    .ZN(_11101_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16149_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(net1509),
    .A3(_11100_),
    .Z(_11102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16150_ (.A1(_11101_),
    .A2(_11102_),
    .Z(_11103_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16151_ (.A1(_10553_),
    .A2(_10566_),
    .Z(_11104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16152_ (.A1(net1530),
    .A2(_11104_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .ZN(_11105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16153_ (.A1(net1532),
    .A2(_11103_),
    .B(_11105_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16154_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16155_ (.A1(_11084_),
    .A2(_03285_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16156_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(net1509),
    .A3(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16157_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(_03286_),
    .B(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16158_ (.A1(net1530),
    .A2(_10587_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16159_ (.A1(net1532),
    .A2(_03288_),
    .B(_03289_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16160_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16161_ (.A1(_11100_),
    .A2(_03290_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16162_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16163_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(net1509),
    .A3(_03291_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16164_ (.A1(_03292_),
    .A2(_03293_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16165_ (.A1(net1530),
    .A2(_10624_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16166_ (.A1(net1532),
    .A2(_03294_),
    .B(_03295_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16167_ (.A1(_10631_),
    .A2(_10646_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16168_ (.A1(net1530),
    .A2(_03296_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16169_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16170_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16171_ (.A1(_03286_),
    .A2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16172_ (.A1(_10376_),
    .A2(_10850_),
    .B(_03300_),
    .C(_03298_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16173_ (.A1(_03298_),
    .A2(_03300_),
    .B(_03301_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16174_ (.A1(net1511),
    .A2(_03302_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16175_ (.A1(_03297_),
    .A2(_03303_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16176_ (.A1(_10653_),
    .A2(_10654_),
    .A3(_10655_),
    .A4(_10661_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16177_ (.A1(net1705),
    .A2(_10652_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16178_ (.A1(_01295_),
    .A2(_03304_),
    .B(_03305_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16179_ (.A1(net1530),
    .A2(_03306_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16180_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16181_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16182_ (.A1(_11079_),
    .A2(_03308_),
    .A3(_03290_),
    .A4(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16183_ (.I(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16184_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16185_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(net1509),
    .A3(_03311_),
    .B(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16186_ (.A1(net1511),
    .A2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16187_ (.A1(_03307_),
    .A2(_03314_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16188_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A3(_03300_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16189_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16190_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .A2(net1509),
    .A3(_03315_),
    .B(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16191_ (.A1(net1511),
    .A2(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16192_ (.A1(_10668_),
    .A2(_10669_),
    .A3(_10670_),
    .A4(_10676_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16193_ (.A1(net1705),
    .A2(_10667_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16194_ (.A1(_01302_),
    .A2(_03319_),
    .B(_03320_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16195_ (.A1(net1530),
    .A2(_03321_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16196_ (.A1(_03318_),
    .A2(_03322_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16197_ (.A1(_10684_),
    .A2(_10697_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16198_ (.A1(net1530),
    .A2(_03323_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16199_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16200_ (.A1(_03310_),
    .A2(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16201_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(_03326_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16202_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(net1509),
    .A3(_03326_),
    .B(_03327_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16203_ (.A1(net1511),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16204_ (.A1(_03324_),
    .A2(_03329_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16205_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A3(_03300_),
    .A4(_03325_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16206_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(net1509),
    .A3(_03330_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16207_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(_03330_),
    .B(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16208_ (.A1(_10706_),
    .A2(_10707_),
    .A3(_10708_),
    .A4(_10714_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16209_ (.A1(net1705),
    .A2(_10705_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16210_ (.A1(_01316_),
    .A2(_03333_),
    .B(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16211_ (.A1(net1530),
    .A2(_03335_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16212_ (.A1(net1532),
    .A2(_03332_),
    .B(_03336_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16213_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A3(_03310_),
    .A4(_03325_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16214_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(net1509),
    .A3(_03337_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16215_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(_03337_),
    .B(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16216_ (.A1(net1530),
    .A2(_10735_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16217_ (.A1(net1532),
    .A2(_03339_),
    .B(_03340_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16218_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A3(_03300_),
    .A4(_03325_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16219_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A3(_03341_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16220_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(_03342_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16221_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .A2(net1509),
    .A3(_03342_),
    .B(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16222_ (.A1(net1511),
    .A2(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16223_ (.A1(net1530),
    .A2(net1517),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16224_ (.A1(_03345_),
    .A2(_03346_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16225_ (.I(_10940_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16226_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ),
    .A3(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ),
    .A4(_10309_),
    .Z(_03348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16227_ (.A1(_10376_),
    .A2(_03348_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16228_ (.A1(_10422_),
    .A2(_03349_),
    .Z(_03350_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16229_ (.A1(net1530),
    .A2(_03350_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16230_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ),
    .A2(net1532),
    .A3(_03349_),
    .Z(_03352_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16231_ (.A1(_10266_),
    .A2(_03347_),
    .B(_03351_),
    .C(_03352_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16232_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A3(_03310_),
    .A4(_03325_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16233_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ),
    .Z(_03354_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16234_ (.A1(_03353_),
    .A2(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16235_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16236_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(net1509),
    .A3(_03355_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16237_ (.A1(_03356_),
    .A2(_03357_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16238_ (.A1(net1530),
    .A2(net1516),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16239_ (.A1(net1532),
    .A2(_03358_),
    .B(_03359_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16240_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A3(_03341_),
    .A4(_03354_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16241_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(net1509),
    .A3(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16242_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(_03360_),
    .B(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16243_ (.A1(_10778_),
    .A2(_10779_),
    .A3(_10780_),
    .A4(_10786_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16244_ (.A1(net1705),
    .A2(_10777_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16245_ (.A1(_01344_),
    .A2(_03363_),
    .B(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16246_ (.A1(net1530),
    .A2(_03365_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16247_ (.A1(net1532),
    .A2(_03362_),
    .B(_03366_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16248_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A3(_03353_),
    .A4(_03354_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16249_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16250_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .A2(net1509),
    .A3(_03367_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16251_ (.A1(_03368_),
    .A2(_03369_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16252_ (.A1(net1530),
    .A2(_10813_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16253_ (.A1(net1532),
    .A2(_03370_),
    .B(_03371_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16254_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16255_ (.A1(_03360_),
    .A2(_03372_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16256_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(net1509),
    .A3(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16257_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .A2(_03373_),
    .B(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16258_ (.A1(net1530),
    .A2(_10846_),
    .B1(net1510),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16259_ (.A1(net1532),
    .A2(_03375_),
    .B(_03376_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16260_ (.A1(_10944_),
    .A2(_10955_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16261_ (.A1(_10376_),
    .A2(_01369_),
    .A3(_10300_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16262_ (.I0(_03378_),
    .I1(_10450_),
    .S(net1532),
    .Z(_03379_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16263_ (.A1(_01369_),
    .A2(net1518),
    .A3(_10300_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16264_ (.I0(_03379_),
    .I1(_03380_),
    .S(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .Z(_03381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16265_ (.A1(_10425_),
    .A2(_03377_),
    .B(_03381_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16266_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .A2(net1518),
    .A3(_10300_),
    .A4(_10309_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16267_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(_10456_),
    .A3(_03382_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16268_ (.A1(_10970_),
    .A2(_10983_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16269_ (.A1(_10456_),
    .A2(_03384_),
    .B1(_03382_),
    .B2(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16270_ (.A1(_03383_),
    .A2(_03385_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16271_ (.A1(_10997_),
    .A2(_11008_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16272_ (.A1(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ),
    .A2(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16273_ (.A1(_03387_),
    .A2(_03380_),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ),
    .C(_10425_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16274_ (.A1(net1518),
    .A2(_10302_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16275_ (.A1(_10425_),
    .A2(_03386_),
    .B(_03388_),
    .C(_03389_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16276_ (.I(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16277_ (.A1(_03390_),
    .A2(_10310_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16278_ (.A1(_10271_),
    .A2(_11024_),
    .B1(_03391_),
    .B2(net1518),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16279_ (.A1(_03390_),
    .A2(_10267_),
    .B(_03392_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16280_ (.A1(_08179_),
    .A2(_08136_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16281_ (.A1(_08140_),
    .A2(_08148_),
    .A3(_08172_),
    .A4(_08178_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16282_ (.A1(_08208_),
    .A2(_08213_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16283_ (.A1(_08155_),
    .A2(_08169_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1455 (.I(net180),
    .Z(net1454));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16285_ (.A1(_03395_),
    .A2(_03396_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16286_ (.A1(_03394_),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16287_ (.A1(_03393_),
    .A2(_03399_),
    .B(_08217_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16288_ (.I(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16289_ (.A1(_09722_),
    .A2(_09739_),
    .B(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16290_ (.A1(_07599_),
    .A2(_09699_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16291_ (.A1(_07711_),
    .A2(_07645_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16292_ (.A1(_08179_),
    .A2(_08136_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16293_ (.A1(_08208_),
    .A2(_08213_),
    .Z(_03406_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16294_ (.A1(_03406_),
    .A2(_03396_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16295_ (.A1(_03405_),
    .A2(_03407_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16296_ (.A1(_03396_),
    .A2(_03394_),
    .Z(_03409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16297_ (.A1(_03396_),
    .A2(_03394_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16298_ (.I0(_03409_),
    .I1(_03410_),
    .S(_03395_),
    .Z(_03411_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16299_ (.A1(_08179_),
    .A2(_08140_),
    .A3(_08172_),
    .A4(_08178_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16300_ (.A1(_03405_),
    .A2(_03411_),
    .B(_03412_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1469 (.I(_05706_),
    .Z(net1468));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16302_ (.A1(_08127_),
    .A2(net1782),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16303_ (.A1(_03396_),
    .A2(_03394_),
    .B(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16304_ (.A1(_03412_),
    .A2(_03409_),
    .B1(_03416_),
    .B2(_03393_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16305_ (.A1(_03395_),
    .A2(_09470_),
    .A3(_03417_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16306_ (.A1(_03395_),
    .A2(_03417_),
    .B(_09470_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16307_ (.A1(_03418_),
    .A2(_03419_),
    .B(_00941_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16308_ (.A1(_00941_),
    .A2(net2106),
    .A3(net2084),
    .B(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16309_ (.I0(_03408_),
    .I1(_03413_),
    .S(_03421_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16310_ (.A1(_08127_),
    .A2(_03403_),
    .A3(_03404_),
    .A4(_03422_),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16311_ (.A1(net169),
    .A2(_09718_),
    .A3(_09719_),
    .A4(_09721_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16312_ (.A1(_09726_),
    .A2(_09729_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16313_ (.A1(net2065),
    .A2(net2169),
    .A3(net174),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16314_ (.A1(_03425_),
    .A2(_09734_),
    .A3(_09736_),
    .B(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16315_ (.A1(_08127_),
    .A2(_10128_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16316_ (.A1(_03424_),
    .A2(_03427_),
    .B(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16317_ (.A1(_07599_),
    .A2(_09654_),
    .B(_10125_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16318_ (.A1(_07642_),
    .A2(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16319_ (.A1(net2032),
    .A2(_09645_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ),
    .C(net2030),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16320_ (.A1(net1815),
    .A2(_03432_),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16321_ (.I(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16322_ (.A1(_09913_),
    .A2(_03434_),
    .B(_09621_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16323_ (.A1(_03431_),
    .A2(_03435_),
    .B(_09538_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16324_ (.A1(_03402_),
    .A2(_03423_),
    .B(_03429_),
    .C(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16325_ (.A1(_09645_),
    .A2(net1826),
    .A3(_09649_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16326_ (.A1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .A2(\cs_registers_i.mcountinhibit_q[2] ),
    .A3(_09658_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16327_ (.A1(_09699_),
    .A2(_03438_),
    .A3(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16328_ (.A1(_09624_),
    .A2(_10370_),
    .B(_08043_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16329_ (.A1(_03440_),
    .A2(_03441_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16330_ (.A1(_10351_),
    .A2(_10372_),
    .A3(_10149_),
    .A4(net1562),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu9t5v0__or3_4 _16331_ (.A1(_03437_),
    .A2(_03442_),
    .A3(_03443_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16332_ (.A1(net1560),
    .A2(_03443_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16333_ (.A1(_03424_),
    .A2(_03427_),
    .B(_03400_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16334_ (.A1(_08127_),
    .A2(_03403_),
    .A3(_03404_),
    .A4(_03422_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16335_ (.A1(_09722_),
    .A2(_09739_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _16336_ (.A1(_03446_),
    .A2(_03447_),
    .B1(_03428_),
    .B2(_03448_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1454 (.I(_05521_),
    .Z(net1453));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1472 (.I(_05698_),
    .Z(net1471));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16339_ (.A1(_09615_),
    .A2(_10228_),
    .A3(_10934_),
    .A4(_10261_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1453 (.I(_00991_),
    .Z(net1452));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1480 (.I(_05675_),
    .Z(net1479));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16342_ (.A1(_09585_),
    .A2(_09637_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16343_ (.A1(_03436_),
    .A2(_03440_),
    .Z(_03456_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _16344_ (.A1(_03449_),
    .A2(net1529),
    .A3(_03455_),
    .A4(_03456_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16345_ (.A1(_10264_),
    .A2(net1529),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1482 (.I(_05664_),
    .Z(net1481));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16347_ (.A1(_10152_),
    .A2(_03457_),
    .A3(net1515),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16348_ (.A1(\cs_registers_i.mhpmcounter[1856] ),
    .A2(_03444_),
    .B1(_03445_),
    .B2(_10273_),
    .C(_03460_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16349_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(\cs_registers_i.mhpmcounter[1858] ),
    .A3(_01367_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16350_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(\cs_registers_i.mhpmcounter[1861] ),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16351_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(_03461_),
    .A3(_03462_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16352_ (.A1(\cs_registers_i.mhpmcounter[1863] ),
    .A2(\cs_registers_i.mhpmcounter[1864] ),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16353_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_03463_),
    .A3(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16354_ (.A1(net1560),
    .A2(_03443_),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16355_ (.I0(_03465_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16356_ (.I(\cs_registers_i.mhpmcounter[1866] ),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1484 (.I(_05634_),
    .Z(net1483));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16358_ (.A1(_03468_),
    .A2(_03457_),
    .A3(_03465_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16359_ (.A1(_10299_),
    .A2(_03445_),
    .B1(_03467_),
    .B2(_03468_),
    .C(_03470_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16360_ (.A1(net2159),
    .A2(_10346_),
    .B(_10315_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16361_ (.A1(\cs_registers_i.mhpmcounter[1857] ),
    .A2(\cs_registers_i.mhpmcounter[1856] ),
    .A3(\cs_registers_i.mhpmcounter[1858] ),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16362_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(\cs_registers_i.mhpmcounter[1862] ),
    .A3(_03462_),
    .A4(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16363_ (.A1(_03464_),
    .A2(_03473_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16364_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(\cs_registers_i.mhpmcounter[1866] ),
    .A3(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16365_ (.I0(_03475_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16366_ (.I(\cs_registers_i.mhpmcounter[1867] ),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16367_ (.A1(_03437_),
    .A2(_03442_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16368_ (.A1(_10351_),
    .A2(_10372_),
    .A3(_10149_),
    .A4(net1562),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16369_ (.A1(_03477_),
    .A2(_03478_),
    .A3(_03479_),
    .A4(_03475_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16370_ (.A1(_03471_),
    .A2(_03445_),
    .B1(_03476_),
    .B2(_03477_),
    .C(_03480_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16371_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(\cs_registers_i.mhpmcounter[1866] ),
    .A3(_03465_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16372_ (.I0(_03481_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16373_ (.I(\cs_registers_i.mhpmcounter[1868] ),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16374_ (.A1(_03483_),
    .A2(_03478_),
    .A3(_03479_),
    .A4(_03481_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16375_ (.A1(_10404_),
    .A2(_03445_),
    .B1(_03482_),
    .B2(_03483_),
    .C(_03484_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16376_ (.A1(_10264_),
    .A2(net1529),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1452 (.I(net156),
    .Z(net1451));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16378_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(\cs_registers_i.mhpmcounter[1867] ),
    .A3(_03475_),
    .Z(_03487_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _16379_ (.A1(\cs_registers_i.mhpmcounter[1869] ),
    .A2(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16380_ (.A1(\cs_registers_i.mhpmcounter[1869] ),
    .A2(_03485_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16381_ (.A1(_03449_),
    .A2(net1529),
    .A3(_03455_),
    .A4(_03456_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1451 (.I(net159),
    .Z(net1450));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16383_ (.I0(_03488_),
    .I1(_03489_),
    .S(net1389),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16384_ (.A1(_10448_),
    .A2(_03485_),
    .B(_03492_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16385_ (.A1(\cs_registers_i.mhpmcounter[1868] ),
    .A2(\cs_registers_i.mhpmcounter[1869] ),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16386_ (.A1(_03481_),
    .A2(_03493_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1450 (.I(net158),
    .Z(net1449));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16388_ (.A1(\cs_registers_i.mhpmcounter[1870] ),
    .A2(_03485_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16389_ (.A1(_03457_),
    .A2(_03494_),
    .B(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16390_ (.I(\cs_registers_i.mhpmcounter[1870] ),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16391_ (.A1(_03498_),
    .A2(_03457_),
    .A3(_03481_),
    .A4(_03493_),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16392_ (.A1(_11064_),
    .A2(net1515),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16393_ (.A1(_03497_),
    .A2(_03499_),
    .A3(_03500_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16394_ (.A1(\cs_registers_i.mhpmcounter[1867] ),
    .A2(\cs_registers_i.mhpmcounter[1865] ),
    .A3(\cs_registers_i.mhpmcounter[1866] ),
    .A4(\cs_registers_i.mhpmcounter[1870] ),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16395_ (.A1(_03474_),
    .A2(_03493_),
    .A3(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16396_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16397_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(_03502_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1449 (.I(net161),
    .Z(net1448));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16399_ (.A1(_03503_),
    .A2(_03504_),
    .B(_03457_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1448 (.I(net163),
    .Z(net1447));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16401_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(_03485_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1447 (.I(net162),
    .Z(net1446));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16403_ (.A1(net1531),
    .A2(net1515),
    .B1(_03508_),
    .B2(net1389),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16404_ (.A1(_03506_),
    .A2(_03510_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16405_ (.A1(\cs_registers_i.mhpmcounter[1871] ),
    .A2(_03464_),
    .A3(_03493_),
    .A4(_03501_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16406_ (.A1(_03463_),
    .A2(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16407_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16408_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03512_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 rebuffer2094 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .Z(net2093));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16410_ (.A1(_03513_),
    .A2(_03514_),
    .B(net1389),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16411_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03490_),
    .A3(_03485_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16412_ (.A1(_11077_),
    .A2(net1515),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16413_ (.A1(_03516_),
    .A2(_03517_),
    .A3(_03518_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2095 (.I(_08504_),
    .Z(net2094));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16415_ (.A1(_03449_),
    .A2(_03455_),
    .A3(_03456_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16416_ (.A1(_10264_),
    .A2(net1535),
    .A3(_10934_),
    .A4(_10261_),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2096 (.I(_00868_),
    .Z(net2095));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16418_ (.I(_03521_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16419_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03473_),
    .A3(_03511_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16420_ (.A1(_03523_),
    .A2(_03524_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16421_ (.A1(_03520_),
    .A2(_03525_),
    .B(_03485_),
    .C(\cs_registers_i.mhpmcounter[1873] ),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16422_ (.I(\cs_registers_i.mhpmcounter[1873] ),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16423_ (.A1(_03527_),
    .A2(_03524_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16424_ (.A1(_11089_),
    .A2(net1515),
    .B1(_03528_),
    .B2(_03457_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16425_ (.A1(_03526_),
    .A2(_03529_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16426_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03463_),
    .A3(_03511_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16427_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16428_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(_03531_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16429_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(_03531_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16430_ (.A1(_03532_),
    .A2(_03533_),
    .B(_03457_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16431_ (.A1(\cs_registers_i.mhpmcounter[1874] ),
    .A2(_03485_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16432_ (.A1(_11104_),
    .A2(net1515),
    .B1(_03535_),
    .B2(net1389),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16433_ (.A1(_03534_),
    .A2(_03536_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16434_ (.A1(_10573_),
    .A2(_10586_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16435_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(\cs_registers_i.mhpmcounter[1874] ),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16436_ (.A1(\cs_registers_i.mhpmcounter[1872] ),
    .A2(_03473_),
    .A3(_03511_),
    .A4(_03538_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16437_ (.I0(_03539_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16438_ (.I(\cs_registers_i.mhpmcounter[1875] ),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16439_ (.A1(_03524_),
    .A2(_03538_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16440_ (.I(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16441_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(net1389),
    .A3(_03543_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16442_ (.A1(_03537_),
    .A2(_03445_),
    .B1(_03540_),
    .B2(_03541_),
    .C(_03544_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16443_ (.A1(\cs_registers_i.mhpmcounter[1857] ),
    .A2(net1389),
    .A3(_03485_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16444_ (.A1(_01368_),
    .A2(_03457_),
    .B1(net1515),
    .B2(_10607_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16445_ (.A1(_03545_),
    .A2(_03546_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16446_ (.A1(_10610_),
    .A2(_10623_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16447_ (.A1(\cs_registers_i.mhpmcounter[1873] ),
    .A2(\cs_registers_i.mhpmcounter[1874] ),
    .A3(\cs_registers_i.mhpmcounter[1875] ),
    .A4(_03530_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16448_ (.I0(_03548_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16449_ (.I(\cs_registers_i.mhpmcounter[1876] ),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16450_ (.A1(_03550_),
    .A2(_03457_),
    .A3(_03548_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16451_ (.A1(_03547_),
    .A2(_03445_),
    .B1(_03549_),
    .B2(_03550_),
    .C(_03551_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16452_ (.A1(net1612),
    .A2(net2289),
    .A3(_09625_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _16453_ (.A1(_10408_),
    .A2(_10421_),
    .A3(_03552_),
    .A4(_10148_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16454_ (.A1(net1528),
    .A2(_03437_),
    .A3(_03442_),
    .A4(_03543_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16455_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(\cs_registers_i.mhpmcounter[1876] ),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16456_ (.A1(_03554_),
    .A2(_03555_),
    .B(\cs_registers_i.mhpmcounter[1877] ),
    .C(_03485_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16457_ (.A1(_03543_),
    .A2(_03555_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16458_ (.A1(\cs_registers_i.mhpmcounter[1877] ),
    .A2(net1389),
    .A3(_03557_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16459_ (.A1(_03296_),
    .A2(net1515),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16460_ (.A1(_03556_),
    .A2(_03558_),
    .A3(_03559_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16461_ (.A1(\cs_registers_i.mhpmcounter[1876] ),
    .A2(\cs_registers_i.mhpmcounter[1877] ),
    .A3(_03548_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16462_ (.I0(_03560_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16463_ (.I(\cs_registers_i.mhpmcounter[1878] ),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16464_ (.A1(_03562_),
    .A2(_03457_),
    .A3(_03560_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16465_ (.A1(_10663_),
    .A2(_03445_),
    .B1(_03561_),
    .B2(_03562_),
    .C(_03563_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16466_ (.I(\cs_registers_i.mhpmcounter[1877] ),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16467_ (.A1(_03564_),
    .A2(_03562_),
    .A3(_03557_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _16468_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(net1389),
    .A3(_03565_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16469_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_03457_),
    .A3(_03565_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16470_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(_03485_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16471_ (.A1(_10678_),
    .A2(_03485_),
    .B1(_03568_),
    .B2(_03457_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16472_ (.A1(_03566_),
    .A2(_03567_),
    .A3(_03569_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16473_ (.A1(\cs_registers_i.mhpmcounter[1878] ),
    .A2(\cs_registers_i.mhpmcounter[1879] ),
    .A3(_03560_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16474_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16475_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(_03570_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16476_ (.A1(_03571_),
    .A2(_03572_),
    .B(_03457_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16477_ (.A1(\cs_registers_i.mhpmcounter[1880] ),
    .A2(_03485_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16478_ (.A1(_03323_),
    .A2(net1515),
    .B1(_03574_),
    .B2(net1389),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16479_ (.A1(_03573_),
    .A2(_03575_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16480_ (.A1(\cs_registers_i.mhpmcounter[1875] ),
    .A2(\cs_registers_i.mhpmcounter[1876] ),
    .A3(\cs_registers_i.mhpmcounter[1877] ),
    .A4(\cs_registers_i.mhpmcounter[1878] ),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16481_ (.A1(\cs_registers_i.mhpmcounter[1879] ),
    .A2(\cs_registers_i.mhpmcounter[1880] ),
    .A3(_03576_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16482_ (.A1(_03539_),
    .A2(_03577_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16483_ (.I0(_03578_),
    .I1(_03466_),
    .S(_03444_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16484_ (.I(\cs_registers_i.mhpmcounter[1881] ),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16485_ (.A1(_03542_),
    .A2(_03577_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16486_ (.I(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16487_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(net1389),
    .A3(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _16488_ (.A1(_10716_),
    .A2(_03445_),
    .B1(_03579_),
    .B2(_03580_),
    .C(_03583_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16489_ (.I(\cs_registers_i.mhpmcounter[1882] ),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16490_ (.A1(\cs_registers_i.mhpmcounter[1881] ),
    .A2(_03538_),
    .A3(_03577_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16491_ (.A1(_03530_),
    .A2(_03585_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16492_ (.A1(_03584_),
    .A2(_03586_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16493_ (.A1(_03584_),
    .A2(_03586_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16494_ (.A1(_03587_),
    .A2(_03588_),
    .B(_03457_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16495_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(_03485_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16496_ (.A1(_10735_),
    .A2(net1515),
    .B1(_03590_),
    .B2(net1389),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16497_ (.A1(_03589_),
    .A2(_03591_),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16498_ (.A1(_03580_),
    .A2(_03584_),
    .A3(_03582_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16499_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16500_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(_03592_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16501_ (.A1(_03593_),
    .A2(_03594_),
    .B(net1389),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16502_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(net1389),
    .A3(_03485_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16503_ (.A1(net1517),
    .A2(net1515),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16504_ (.A1(_03595_),
    .A2(_03596_),
    .A3(_03597_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16505_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(\cs_registers_i.mhpmcounter[1883] ),
    .A3(_03586_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16506_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(_03598_),
    .Z(_03599_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16507_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(_03598_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16508_ (.A1(_03599_),
    .A2(_03600_),
    .B(_03457_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16509_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(_03485_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16510_ (.A1(net1516),
    .A2(net1515),
    .B1(_03602_),
    .B2(net1389),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16511_ (.A1(_03601_),
    .A2(_03603_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2097 (.I(_01229_),
    .Z(net2096));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16513_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(net1529),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16514_ (.I(net1529),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16515_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(_03606_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16516_ (.I(_03592_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16517_ (.A1(\cs_registers_i.mhpmcounter[1883] ),
    .A2(\cs_registers_i.mhpmcounter[1884] ),
    .A3(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16518_ (.A1(_03449_),
    .A2(_03455_),
    .A3(_03456_),
    .A4(_03609_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16519_ (.I0(_03605_),
    .I1(_03607_),
    .S(_03610_),
    .Z(_03611_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2098 (.I(net1689),
    .Z(net2097));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16521_ (.A1(\cs_registers_i.mhpmcounter[1885] ),
    .A2(_03521_),
    .B1(net1515),
    .B2(_03365_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16522_ (.A1(_03611_),
    .A2(_03613_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16523_ (.A1(\cs_registers_i.mhpmcounter[1858] ),
    .A2(_03485_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16524_ (.I(_01367_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16525_ (.A1(\cs_registers_i.mhpmcounter[1858] ),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16526_ (.I0(_03614_),
    .I1(_03616_),
    .S(_03457_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16527_ (.A1(\cs_registers_i.mhpmcounter[1858] ),
    .A2(_03615_),
    .A3(net1389),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16528_ (.A1(_10792_),
    .A2(_03485_),
    .B(_03617_),
    .C(_03618_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16529_ (.A1(\cs_registers_i.mhpmcounter[1884] ),
    .A2(\cs_registers_i.mhpmcounter[1885] ),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16530_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(_03490_),
    .A3(_03598_),
    .A4(_03619_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16531_ (.A1(_03598_),
    .A2(_03619_),
    .B(\cs_registers_i.mhpmcounter[1886] ),
    .C(_03457_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16532_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(_03485_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16533_ (.A1(_10813_),
    .A2(net1515),
    .B1(_03622_),
    .B2(_03490_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16534_ (.A1(_03620_),
    .A2(_03621_),
    .A3(_03623_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16535_ (.A1(\cs_registers_i.mhpmcounter[1882] ),
    .A2(\cs_registers_i.mhpmcounter[1883] ),
    .A3(\cs_registers_i.mhpmcounter[1884] ),
    .A4(\cs_registers_i.mhpmcounter[1885] ),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16536_ (.A1(\cs_registers_i.mhpmcounter[1886] ),
    .A2(_03624_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16537_ (.A1(_03524_),
    .A2(_03585_),
    .A3(_03625_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16538_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(_03626_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16539_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(_03626_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16540_ (.A1(_03627_),
    .A2(_03628_),
    .B(_03457_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16541_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(_03485_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16542_ (.A1(_10846_),
    .A2(net1515),
    .B1(_03630_),
    .B2(net1389),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16543_ (.A1(_03629_),
    .A2(_03631_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16544_ (.A1(_10264_),
    .A2(net1535),
    .A3(_10934_),
    .A4(_10261_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16545_ (.A1(_03490_),
    .A2(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2099 (.I(\load_store_unit_i.ls_fsm_cs[0] ),
    .Z(net2098));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16547_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(_03586_),
    .A3(_03625_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16548_ (.A1(_10164_),
    .A2(net1529),
    .A3(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16549_ (.A1(_10225_),
    .A2(_03521_),
    .B(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16550_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(_03632_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16551_ (.I(_03635_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16552_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(net1529),
    .A3(_03639_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16553_ (.A1(net1389),
    .A2(_03638_),
    .B(_03640_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16554_ (.A1(_03633_),
    .A2(_03637_),
    .B(_03641_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16555_ (.I(\cs_registers_i.mhpmcounter[1889] ),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16556_ (.A1(_10423_),
    .A2(_10421_),
    .A3(_03552_),
    .A4(_10148_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _16557_ (.A1(net1528),
    .A2(_03437_),
    .A3(_03442_),
    .B(_03643_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16558_ (.A1(_10408_),
    .A2(_10421_),
    .A3(_03552_),
    .A4(_10148_),
    .Z(_03645_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2100 (.I(\load_store_unit_i.ls_fsm_cs[0] ),
    .Z(net2099));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16560_ (.A1(\cs_registers_i.mhpmcounter[1887] ),
    .A2(_03524_),
    .A3(_03585_),
    .A4(_03625_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16561_ (.A1(\cs_registers_i.mhpmcounter[1888] ),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16562_ (.A1(_03645_),
    .A2(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16563_ (.A1(_03644_),
    .A2(_03649_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2101 (.I(_08041_),
    .Z(net2100));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16565_ (.A1(_03642_),
    .A2(\cs_registers_i.mhpmcounter[1888] ),
    .A3(net1529),
    .A4(_03647_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16566_ (.A1(_01145_),
    .A2(_10605_),
    .B(_10595_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16567_ (.A1(_03653_),
    .A2(_03643_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16568_ (.A1(_03644_),
    .A2(_03652_),
    .B(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16569_ (.A1(_03642_),
    .A2(_03650_),
    .B(_03655_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16570_ (.I(\cs_registers_i.mhpmcounter[1890] ),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16571_ (.A1(_03642_),
    .A2(_10164_),
    .A3(_03639_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16572_ (.A1(_03645_),
    .A2(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16573_ (.A1(_03644_),
    .A2(_03658_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16574_ (.A1(\cs_registers_i.mhpmcounter[1890] ),
    .A2(_03657_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16575_ (.A1(_10258_),
    .A2(_03521_),
    .B1(_03660_),
    .B2(net1529),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16576_ (.A1(_03656_),
    .A2(_03659_),
    .B1(_03661_),
    .B2(_03633_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16577_ (.I(\cs_registers_i.mhpmcounter[1891] ),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16578_ (.A1(_03642_),
    .A2(_03656_),
    .A3(_03648_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16579_ (.A1(_03645_),
    .A2(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16580_ (.A1(_03644_),
    .A2(_03664_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16581_ (.A1(\cs_registers_i.mhpmcounter[1891] ),
    .A2(_03663_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16582_ (.A1(_10264_),
    .A2(_03606_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16583_ (.A1(net1529),
    .A2(_03666_),
    .B1(_03667_),
    .B2(_10891_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16584_ (.A1(_03662_),
    .A2(_03665_),
    .B1(_03668_),
    .B2(_03633_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16585_ (.I(\cs_registers_i.mhpmcounter[1892] ),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16586_ (.A1(\cs_registers_i.mhpmcounter[1889] ),
    .A2(\cs_registers_i.mhpmcounter[1888] ),
    .A3(\cs_registers_i.mhpmcounter[1891] ),
    .A4(\cs_registers_i.mhpmcounter[1890] ),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16587_ (.A1(_03635_),
    .A2(_03670_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16588_ (.A1(net1528),
    .A2(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16589_ (.A1(_03644_),
    .A2(_03672_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16590_ (.A1(_03669_),
    .A2(net1529),
    .A3(_03671_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16591_ (.A1(_10911_),
    .A2(_03521_),
    .B(_03674_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16592_ (.A1(_03669_),
    .A2(_03673_),
    .B1(_03675_),
    .B2(_03633_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16593_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(_03647_),
    .A3(_03670_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16594_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2102 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net2101));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16596_ (.A1(_10940_),
    .A2(_03521_),
    .B1(_03677_),
    .B2(net1529),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16597_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(_03632_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16598_ (.A1(\cs_registers_i.mhpmcounter[1893] ),
    .A2(net1529),
    .A3(_03676_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16599_ (.A1(net1389),
    .A2(_03680_),
    .B(_03681_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16600_ (.A1(_03633_),
    .A2(_03679_),
    .B(_03682_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16601_ (.I(\cs_registers_i.mhpmcounter[1894] ),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16602_ (.A1(\cs_registers_i.mhpmcounter[1892] ),
    .A2(\cs_registers_i.mhpmcounter[1893] ),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16603_ (.A1(_03671_),
    .A2(_03684_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16604_ (.A1(net1528),
    .A2(_03685_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16605_ (.A1(_03644_),
    .A2(_03686_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16606_ (.A1(_03683_),
    .A2(net1529),
    .A3(_03671_),
    .A4(_03684_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16607_ (.A1(_10956_),
    .A2(_03521_),
    .B(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16608_ (.A1(_03683_),
    .A2(_03687_),
    .B1(_03689_),
    .B2(_03633_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16609_ (.A1(\cs_registers_i.mhpmcounter[1894] ),
    .A2(_03670_),
    .A3(_03684_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16610_ (.A1(_03647_),
    .A2(_03690_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16611_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16612_ (.A1(_10984_),
    .A2(_03521_),
    .B1(_03692_),
    .B2(_03479_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16613_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(_03632_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16614_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(net1529),
    .A3(_03691_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16615_ (.A1(net1389),
    .A2(_03694_),
    .B(_03695_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16616_ (.A1(_03633_),
    .A2(_03693_),
    .B(_03696_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16617_ (.I(\cs_registers_i.mhpmcounter[1859] ),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16618_ (.A1(_03697_),
    .A2(_03472_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16619_ (.A1(_03697_),
    .A2(_03472_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16620_ (.A1(_03698_),
    .A2(_03699_),
    .B(_03457_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16621_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(_03485_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16622_ (.A1(_10891_),
    .A2(net1515),
    .B1(_03701_),
    .B2(net1389),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16623_ (.A1(_03700_),
    .A2(_03702_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16624_ (.I(\cs_registers_i.mhpmcounter[1896] ),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16625_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(_03635_),
    .A3(_03690_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16626_ (.A1(_03645_),
    .A2(_03704_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16627_ (.A1(_03644_),
    .A2(_03705_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16628_ (.I(_03704_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16629_ (.A1(_03703_),
    .A2(_03707_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16630_ (.A1(_11009_),
    .A2(_03521_),
    .B1(_03708_),
    .B2(net1529),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16631_ (.A1(_03703_),
    .A2(_03706_),
    .B1(_03709_),
    .B2(_03633_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16632_ (.A1(_03490_),
    .A2(_03632_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1446 (.I(_01010_),
    .Z(net1445));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1445 (.I(_01011_),
    .Z(net1444));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16635_ (.A1(\cs_registers_i.mhpmcounter[1895] ),
    .A2(\cs_registers_i.mhpmcounter[1896] ),
    .A3(_03647_),
    .A4(_03690_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16636_ (.A1(\cs_registers_i.mhpmcounter[1897] ),
    .A2(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16637_ (.I(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16638_ (.A1(_11024_),
    .A2(_03667_),
    .B1(_03715_),
    .B2(net1529),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _16639_ (.A1(_10454_),
    .A2(_10372_),
    .A3(_10149_),
    .A4(net1562),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16640_ (.A1(_03437_),
    .A2(_03442_),
    .A3(_03443_),
    .B(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16641_ (.A1(_03443_),
    .A2(_03713_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16642_ (.A1(_03718_),
    .A2(_03719_),
    .B(\cs_registers_i.mhpmcounter[1897] ),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16643_ (.A1(_03710_),
    .A2(_03716_),
    .B(_03720_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16644_ (.A1(\cs_registers_i.mhpmcounter[1896] ),
    .A2(\cs_registers_i.mhpmcounter[1897] ),
    .A3(_03707_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16645_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16646_ (.A1(_11033_),
    .A2(_03521_),
    .B1(_03722_),
    .B2(net1529),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16647_ (.I(\cs_registers_i.mhpmcounter[1898] ),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16648_ (.A1(_03724_),
    .A2(_03632_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _16649_ (.A1(\cs_registers_i.mhpmcounter[1898] ),
    .A2(_03606_),
    .A3(_03721_),
    .B1(_03725_),
    .B2(_03457_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16650_ (.A1(_03710_),
    .A2(_03723_),
    .B(_03726_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16651_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(\cs_registers_i.mhpmcounter[1898] ),
    .A3(_03714_),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16652_ (.I(_03727_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16653_ (.A1(_10348_),
    .A2(_03667_),
    .B1(_03728_),
    .B2(net1529),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16654_ (.A1(_03724_),
    .A2(_03715_),
    .B(_03479_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16655_ (.A1(_03718_),
    .A2(_03730_),
    .B(\cs_registers_i.mhpmcounter[1899] ),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16656_ (.A1(_03710_),
    .A2(_03729_),
    .B(_03731_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16657_ (.A1(\cs_registers_i.mhpmcounter[1899] ),
    .A2(\cs_registers_i.mhpmcounter[1898] ),
    .A3(_03721_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16658_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(_03732_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16659_ (.A1(_11052_),
    .A2(_03667_),
    .B1(_03733_),
    .B2(net1529),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16660_ (.A1(net1528),
    .A2(_03732_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16661_ (.A1(_03644_),
    .A2(_03735_),
    .B(\cs_registers_i.mhpmcounter[1900] ),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16662_ (.A1(_03710_),
    .A2(_03734_),
    .B(_03736_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16663_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(\cs_registers_i.mhpmcounter[1901] ),
    .A3(_03727_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16664_ (.I(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16665_ (.A1(_11059_),
    .A2(_03667_),
    .B1(_03738_),
    .B2(net1529),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16666_ (.I(\cs_registers_i.mhpmcounter[1900] ),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16667_ (.A1(_03740_),
    .A2(_03728_),
    .B(_03479_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16668_ (.A1(_03718_),
    .A2(_03741_),
    .B(\cs_registers_i.mhpmcounter[1901] ),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16669_ (.A1(_03710_),
    .A2(_03739_),
    .B(_03742_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16670_ (.I(\cs_registers_i.mhpmcounter[1902] ),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16671_ (.A1(\cs_registers_i.mhpmcounter[1900] ),
    .A2(\cs_registers_i.mhpmcounter[1901] ),
    .A3(_03732_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16672_ (.A1(net1528),
    .A2(_03744_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16673_ (.A1(_03644_),
    .A2(_03745_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16674_ (.A1(_03743_),
    .A2(net1529),
    .A3(_03744_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16675_ (.A1(_11064_),
    .A2(_03521_),
    .B(_03747_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _16676_ (.A1(_03743_),
    .A2(_03746_),
    .B1(_03748_),
    .B2(_03633_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16677_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(\cs_registers_i.mhpmcounter[1903] ),
    .A3(_03737_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16678_ (.A1(net1531),
    .A2(_03667_),
    .B1(_03749_),
    .B2(net1529),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16679_ (.A1(_03743_),
    .A2(_03738_),
    .B(_03479_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16680_ (.A1(_03718_),
    .A2(_03751_),
    .B(\cs_registers_i.mhpmcounter[1903] ),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16681_ (.A1(_03710_),
    .A2(_03750_),
    .B(_03752_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16682_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(\cs_registers_i.mhpmcounter[1903] ),
    .A3(\cs_registers_i.mhpmcounter[1904] ),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16683_ (.A1(_03744_),
    .A2(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16684_ (.A1(_11077_),
    .A2(_03667_),
    .B1(_03754_),
    .B2(net1529),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16685_ (.A1(\cs_registers_i.mhpmcounter[1902] ),
    .A2(\cs_registers_i.mhpmcounter[1903] ),
    .A3(_03744_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16686_ (.A1(net1528),
    .A2(_03756_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16687_ (.A1(_03644_),
    .A2(_03757_),
    .B(\cs_registers_i.mhpmcounter[1904] ),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16688_ (.A1(_03710_),
    .A2(_03755_),
    .B(_03758_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16689_ (.A1(\cs_registers_i.mhpmcounter[1905] ),
    .A2(_03753_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16690_ (.A1(_03737_),
    .A2(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16691_ (.A1(_11089_),
    .A2(_03667_),
    .B1(_03760_),
    .B2(net1529),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16692_ (.A1(_03737_),
    .A2(_03753_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16693_ (.A1(_03645_),
    .A2(_03762_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16694_ (.A1(_03644_),
    .A2(_03763_),
    .B(\cs_registers_i.mhpmcounter[1905] ),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16695_ (.A1(_03710_),
    .A2(_03761_),
    .B(_03764_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16696_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(\cs_registers_i.mhpmcounter[1858] ),
    .A3(_01367_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _16697_ (.A1(_03437_),
    .A2(_03442_),
    .A3(_03765_),
    .B(_03479_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16698_ (.I(\cs_registers_i.mhpmcounter[1860] ),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16699_ (.A1(_03717_),
    .A2(_03766_),
    .B(_03767_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _16700_ (.A1(\cs_registers_i.mhpmcounter[1860] ),
    .A2(net1389),
    .A3(_03765_),
    .B1(_03485_),
    .B2(_11093_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16701_ (.A1(_03768_),
    .A2(_03769_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16702_ (.A1(\cs_registers_i.mhpmcounter[1906] ),
    .A2(_03759_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16703_ (.A1(_03744_),
    .A2(_03770_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16704_ (.I(_03771_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16705_ (.A1(_11104_),
    .A2(_03667_),
    .B1(_03772_),
    .B2(net1529),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16706_ (.A1(_03744_),
    .A2(_03759_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16707_ (.A1(_03645_),
    .A2(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16708_ (.A1(_03644_),
    .A2(_03775_),
    .B(\cs_registers_i.mhpmcounter[1906] ),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16709_ (.A1(_03710_),
    .A2(_03773_),
    .B(_03776_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16710_ (.A1(_03737_),
    .A2(_03770_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16711_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2103 (.I(net1688),
    .Z(net2102));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16713_ (.A1(_10587_),
    .A2(_03521_),
    .B1(_03778_),
    .B2(net1529),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16714_ (.A1(_03443_),
    .A2(_03777_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16715_ (.A1(_03718_),
    .A2(_03781_),
    .B(\cs_registers_i.mhpmcounter[1907] ),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16716_ (.A1(_03710_),
    .A2(_03780_),
    .B(_03782_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1444 (.I(_01022_),
    .Z(net1443));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16718_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(\cs_registers_i.mhpmcounter[1908] ),
    .A3(_03771_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16719_ (.A1(_10624_),
    .A2(_03667_),
    .B1(_03784_),
    .B2(net1529),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16720_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(_03771_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16721_ (.A1(_03645_),
    .A2(_03786_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16722_ (.A1(_03644_),
    .A2(_03787_),
    .B(\cs_registers_i.mhpmcounter[1908] ),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16723_ (.A1(_03710_),
    .A2(_03785_),
    .B(_03788_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16724_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(\cs_registers_i.mhpmcounter[1908] ),
    .A3(\cs_registers_i.mhpmcounter[1909] ),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16725_ (.A1(_03777_),
    .A2(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16726_ (.A1(_03296_),
    .A2(_03667_),
    .B1(_03790_),
    .B2(net1529),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16727_ (.A1(\cs_registers_i.mhpmcounter[1907] ),
    .A2(\cs_registers_i.mhpmcounter[1908] ),
    .A3(_03777_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16728_ (.A1(_03443_),
    .A2(_03792_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16729_ (.A1(_03718_),
    .A2(_03793_),
    .B(\cs_registers_i.mhpmcounter[1909] ),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16730_ (.A1(_03710_),
    .A2(_03791_),
    .B(_03794_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16731_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(_03771_),
    .A3(_03789_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16732_ (.I(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16733_ (.A1(_03306_),
    .A2(_03667_),
    .B1(_03796_),
    .B2(net1529),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16734_ (.A1(_03771_),
    .A2(_03789_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16735_ (.A1(_03645_),
    .A2(_03798_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16736_ (.A1(_03644_),
    .A2(_03799_),
    .B(\cs_registers_i.mhpmcounter[1910] ),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16737_ (.A1(_03710_),
    .A2(_03797_),
    .B(_03800_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16738_ (.A1(\cs_registers_i.mhpmcounter[1910] ),
    .A2(_03777_),
    .A3(_03789_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16739_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16740_ (.A1(_03321_),
    .A2(_03667_),
    .B1(_03802_),
    .B2(net1529),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16741_ (.A1(_03443_),
    .A2(_03801_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16742_ (.A1(_03718_),
    .A2(_03804_),
    .B(\cs_registers_i.mhpmcounter[1911] ),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16743_ (.A1(_03710_),
    .A2(_03803_),
    .B(_03805_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _16744_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(\cs_registers_i.mhpmcounter[1912] ),
    .A3(_03795_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16745_ (.A1(_03323_),
    .A2(_03521_),
    .B1(_03806_),
    .B2(net1529),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16746_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(_03795_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16747_ (.A1(_03645_),
    .A2(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16748_ (.A1(_03644_),
    .A2(_03809_),
    .B(\cs_registers_i.mhpmcounter[1912] ),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16749_ (.A1(_03710_),
    .A2(_03807_),
    .B(_03810_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16750_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(\cs_registers_i.mhpmcounter[1912] ),
    .A3(\cs_registers_i.mhpmcounter[1913] ),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16751_ (.A1(_03801_),
    .A2(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16752_ (.A1(_03335_),
    .A2(_03667_),
    .B1(_03812_),
    .B2(net1529),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16753_ (.A1(\cs_registers_i.mhpmcounter[1911] ),
    .A2(\cs_registers_i.mhpmcounter[1912] ),
    .A3(_03801_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16754_ (.A1(_03443_),
    .A2(_03814_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16755_ (.A1(_03718_),
    .A2(_03815_),
    .B(\cs_registers_i.mhpmcounter[1913] ),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16756_ (.A1(_03710_),
    .A2(_03813_),
    .B(_03816_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16757_ (.A1(\cs_registers_i.mhpmcounter[1914] ),
    .A2(_03811_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16758_ (.A1(_03795_),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16759_ (.A1(_10735_),
    .A2(_03667_),
    .B1(_03818_),
    .B2(net1529),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16760_ (.A1(_03795_),
    .A2(_03811_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16761_ (.A1(_03645_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16762_ (.A1(_03644_),
    .A2(_03821_),
    .B(\cs_registers_i.mhpmcounter[1914] ),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16763_ (.A1(_03710_),
    .A2(_03819_),
    .B(_03822_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16764_ (.I(\cs_registers_i.mhpmcounter[1915] ),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16765_ (.A1(_03801_),
    .A2(_03817_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16766_ (.A1(_03823_),
    .A2(net1529),
    .A3(_03824_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16767_ (.A1(net1517),
    .A2(_03521_),
    .B(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16768_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(_03632_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16769_ (.I(_03824_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16770_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(net1529),
    .A3(_03828_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16771_ (.A1(_03490_),
    .A2(_03827_),
    .B(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16772_ (.A1(_03633_),
    .A2(_03826_),
    .B(_03830_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16773_ (.A1(\cs_registers_i.mhpmcounter[1859] ),
    .A2(\cs_registers_i.mhpmcounter[1860] ),
    .A3(_03472_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16774_ (.A1(\cs_registers_i.mhpmcounter[1861] ),
    .A2(net1515),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16775_ (.A1(_03457_),
    .A2(_03831_),
    .B(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16776_ (.A1(\cs_registers_i.mhpmcounter[1861] ),
    .A2(_03457_),
    .A3(_03831_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16777_ (.A1(_03347_),
    .A2(net1515),
    .B(_03833_),
    .C(_03834_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16778_ (.A1(_03795_),
    .A2(_03817_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16779_ (.A1(\cs_registers_i.mhpmcounter[1915] ),
    .A2(\cs_registers_i.mhpmcounter[1916] ),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16780_ (.A1(_03835_),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16781_ (.A1(net1516),
    .A2(_03521_),
    .B1(_03837_),
    .B2(net1529),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16782_ (.A1(_03823_),
    .A2(_03818_),
    .B(_03645_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16783_ (.A1(_03644_),
    .A2(_03839_),
    .B(\cs_registers_i.mhpmcounter[1916] ),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16784_ (.A1(_03710_),
    .A2(_03838_),
    .B(_03840_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16785_ (.A1(\cs_registers_i.mhpmcounter[1917] ),
    .A2(_03836_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16786_ (.A1(_03828_),
    .A2(_03841_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16787_ (.A1(_03365_),
    .A2(_03667_),
    .B1(_03842_),
    .B2(net1529),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16788_ (.A1(_03824_),
    .A2(_03836_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16789_ (.A1(_03645_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16790_ (.A1(_03644_),
    .A2(_03845_),
    .B(\cs_registers_i.mhpmcounter[1917] ),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16791_ (.A1(_03710_),
    .A2(_03843_),
    .B(_03846_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16792_ (.A1(\cs_registers_i.mhpmcounter[1917] ),
    .A2(\cs_registers_i.mhpmcounter[1918] ),
    .A3(_03836_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16793_ (.A1(_03835_),
    .A2(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16794_ (.A1(_10813_),
    .A2(_03521_),
    .B1(_03848_),
    .B2(net1529),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16795_ (.A1(_03818_),
    .A2(_03841_),
    .B(_03645_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16796_ (.A1(_03644_),
    .A2(_03850_),
    .B(\cs_registers_i.mhpmcounter[1918] ),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16797_ (.A1(_03710_),
    .A2(_03849_),
    .B(_03851_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16798_ (.I(\cs_registers_i.mhpmcounter[1919] ),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _16799_ (.A1(_03852_),
    .A2(net1529),
    .A3(_03824_),
    .A4(_03847_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16800_ (.A1(_10846_),
    .A2(_03521_),
    .B(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16801_ (.A1(\cs_registers_i.mhpmcounter[1919] ),
    .A2(_03632_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16802_ (.A1(_03824_),
    .A2(_03847_),
    .B(_03852_),
    .C(_03606_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16803_ (.A1(_03490_),
    .A2(_03855_),
    .B(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16804_ (.A1(_03633_),
    .A2(_03854_),
    .B(_03857_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16805_ (.A1(_03461_),
    .A2(_03462_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16806_ (.A1(\cs_registers_i.mhpmcounter[1862] ),
    .A2(net1515),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16807_ (.A1(_03457_),
    .A2(_03858_),
    .B(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _16808_ (.A1(_03377_),
    .A2(net1515),
    .B1(_03463_),
    .B2(_03457_),
    .C(_03860_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16809_ (.A1(_03523_),
    .A2(_03473_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16810_ (.A1(_03520_),
    .A2(_03861_),
    .B(_03485_),
    .C(\cs_registers_i.mhpmcounter[1863] ),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16811_ (.I(_03473_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16812_ (.A1(\cs_registers_i.mhpmcounter[1863] ),
    .A2(net1389),
    .A3(_03863_),
    .Z(_03864_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _16813_ (.A1(_03384_),
    .A2(_03485_),
    .B(_03862_),
    .C(_03864_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16814_ (.A1(\cs_registers_i.mhpmcounter[1863] ),
    .A2(_03463_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _16815_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(net1515),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16816_ (.A1(_03457_),
    .A2(_03865_),
    .B(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16817_ (.A1(\cs_registers_i.mhpmcounter[1864] ),
    .A2(_03457_),
    .A3(_03865_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _16818_ (.A1(_03386_),
    .A2(net1515),
    .B(_03867_),
    .C(_03868_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16819_ (.A1(_03464_),
    .A2(_03473_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16820_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16821_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_03869_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _16822_ (.A1(_03870_),
    .A2(_03871_),
    .B(_03457_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16823_ (.A1(\cs_registers_i.mhpmcounter[1865] ),
    .A2(_03485_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16824_ (.A1(_11024_),
    .A2(net1515),
    .B1(_03873_),
    .B2(net1389),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16825_ (.A1(_03872_),
    .A2(_03874_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1443 (.I(_01023_),
    .Z(net1442));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16827_ (.A1(_09905_),
    .A2(_09943_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16828_ (.A1(_09497_),
    .A2(_09919_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16829_ (.A1(_03876_),
    .A2(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16830_ (.A1(_09922_),
    .A2(_03878_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16831_ (.A1(_09906_),
    .A2(_09908_),
    .A3(_03438_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16832_ (.A1(_03880_),
    .A2(_09996_),
    .B(_09945_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16833_ (.A1(net1617),
    .A2(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16834_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(_03882_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16835_ (.A1(net1747),
    .A2(net1746),
    .A3(_03883_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16836_ (.A1(\cs_registers_i.dcsr_q[0] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.mstatus_q[2] ),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16837_ (.A1(_03884_),
    .A2(_03885_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _16838_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(_03882_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _16839_ (.A1(net1747),
    .A2(net1746),
    .A3(_03886_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16840_ (.A1(\cs_registers_i.dcsr_q[1] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.mstatus_q[3] ),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16841_ (.A1(_03887_),
    .A2(_03888_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16842_ (.I(\cs_registers_i.dcsr_q[0] ),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16843_ (.A1(_10372_),
    .A2(_10201_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16844_ (.A1(_09558_),
    .A2(net1608),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16845_ (.A1(_10929_),
    .A2(net1535),
    .A3(_03891_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _16846_ (.A1(_10273_),
    .A2(_03653_),
    .A3(_03892_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16847_ (.A1(_03889_),
    .A2(_03890_),
    .B(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1442 (.I(_01027_),
    .Z(net1441));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16849_ (.I0(\cs_registers_i.priv_mode_id_o[0] ),
    .I1(_03894_),
    .S(net1617),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16850_ (.I0(\cs_registers_i.dcsr_q[11] ),
    .I1(_10348_),
    .S(_03892_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16851_ (.I0(\cs_registers_i.dcsr_q[12] ),
    .I1(_11052_),
    .S(_03892_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16852_ (.I0(\cs_registers_i.dcsr_q[13] ),
    .I1(_11059_),
    .S(_03892_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16853_ (.I0(\cs_registers_i.dcsr_q[15] ),
    .I1(net1531),
    .S(_03892_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16854_ (.I(\cs_registers_i.dcsr_q[1] ),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _16855_ (.A1(_03896_),
    .A2(_03890_),
    .B(_03893_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16856_ (.I0(\cs_registers_i.priv_mode_id_o[1] ),
    .I1(_03897_),
    .S(net1617),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16857_ (.I0(\cs_registers_i.dcsr_q[2] ),
    .I1(_10258_),
    .S(_03892_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16858_ (.I(\cs_registers_i.dcsr_q[6] ),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16859_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_09923_),
    .B1(net1617),
    .B2(_03898_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16860_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_03879_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16861_ (.I(net65),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16862_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_09921_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _16863_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_03900_),
    .A3(\cs_registers_i.dcsr_q[2] ),
    .A4(_03901_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _16864_ (.A1(_03899_),
    .A2(_03902_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _16865_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_09923_),
    .B1(net1617),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16866_ (.I(_03903_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2104 (.I(_01158_),
    .Z(net2103));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16868_ (.I0(\cs_registers_i.pc_if_i[10] ),
    .I1(\cs_registers_i.pc_id_i[10] ),
    .S(net1708),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16869_ (.A1(net1535),
    .A2(_10936_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1441 (.I(_01032_),
    .Z(net1440));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16871_ (.I0(\cs_registers_i.csr_depc_o[10] ),
    .I1(_11033_),
    .S(_03906_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16872_ (.I0(_03905_),
    .I1(_03908_),
    .S(net1617),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16873_ (.I0(\cs_registers_i.pc_if_i[11] ),
    .I1(\cs_registers_i.pc_id_i[11] ),
    .S(net1708),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16874_ (.I0(\cs_registers_i.csr_depc_o[11] ),
    .I1(_10348_),
    .S(net1527),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16875_ (.I0(_03909_),
    .I1(_03910_),
    .S(net1617),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16876_ (.I0(\cs_registers_i.pc_if_i[12] ),
    .I1(\cs_registers_i.pc_id_i[12] ),
    .S(net1708),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16877_ (.I0(\cs_registers_i.csr_depc_o[12] ),
    .I1(_11052_),
    .S(net1527),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16878_ (.I0(_03911_),
    .I1(_03912_),
    .S(net1617),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16879_ (.I0(\cs_registers_i.pc_if_i[13] ),
    .I1(\cs_registers_i.pc_id_i[13] ),
    .S(net1708),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16880_ (.I0(\cs_registers_i.csr_depc_o[13] ),
    .I1(_11059_),
    .S(_03906_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16881_ (.I0(_03913_),
    .I1(_03914_),
    .S(net1617),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16882_ (.I0(\cs_registers_i.pc_if_i[14] ),
    .I1(\cs_registers_i.pc_id_i[14] ),
    .S(net1708),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16883_ (.I0(\cs_registers_i.csr_depc_o[14] ),
    .I1(_11064_),
    .S(net1527),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16884_ (.I0(_03915_),
    .I1(_03916_),
    .S(_03879_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16885_ (.I0(\cs_registers_i.pc_if_i[15] ),
    .I1(\cs_registers_i.pc_id_i[15] ),
    .S(net1708),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16886_ (.I0(\cs_registers_i.csr_depc_o[15] ),
    .I1(net1531),
    .S(net1527),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1440 (.I(_01033_),
    .Z(net1439));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16888_ (.I0(_03917_),
    .I1(_03918_),
    .S(_03879_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16889_ (.I0(\cs_registers_i.pc_if_i[16] ),
    .I1(\cs_registers_i.pc_id_i[16] ),
    .S(net1708),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16890_ (.I0(\cs_registers_i.csr_depc_o[16] ),
    .I1(_11077_),
    .S(_03906_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16891_ (.I0(_03920_),
    .I1(_03921_),
    .S(net1617),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16892_ (.I0(\cs_registers_i.pc_if_i[17] ),
    .I1(\cs_registers_i.pc_id_i[17] ),
    .S(net1708),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16893_ (.I0(\cs_registers_i.csr_depc_o[17] ),
    .I1(_11089_),
    .S(net1527),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16894_ (.I0(_03922_),
    .I1(_03923_),
    .S(_03879_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16895_ (.I0(\cs_registers_i.pc_if_i[18] ),
    .I1(\cs_registers_i.pc_id_i[18] ),
    .S(net1708),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16896_ (.I0(\cs_registers_i.csr_depc_o[18] ),
    .I1(_11104_),
    .S(_03906_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16897_ (.I0(_03924_),
    .I1(_03925_),
    .S(net1617),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1439 (.I(_01034_),
    .Z(net1438));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16899_ (.I0(\cs_registers_i.pc_if_i[19] ),
    .I1(\cs_registers_i.pc_id_i[19] ),
    .S(net1708),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16900_ (.I0(\cs_registers_i.csr_depc_o[19] ),
    .I1(_10587_),
    .S(_03906_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16901_ (.I0(_03927_),
    .I1(_03928_),
    .S(_03879_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16902_ (.I0(net2026),
    .I1(\cs_registers_i.pc_id_i[1] ),
    .S(net1708),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1438 (.I(_01035_),
    .Z(net1437));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16904_ (.I0(\cs_registers_i.csr_depc_o[1] ),
    .I1(_10607_),
    .S(net1527),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16905_ (.I0(_03929_),
    .I1(_03931_),
    .S(net1617),
    .Z(_01535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16906_ (.I0(\cs_registers_i.pc_if_i[20] ),
    .I1(\cs_registers_i.pc_id_i[20] ),
    .S(net1708),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16907_ (.I0(\cs_registers_i.csr_depc_o[20] ),
    .I1(_10624_),
    .S(_03906_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16908_ (.I0(_03932_),
    .I1(_03933_),
    .S(net1617),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16909_ (.I0(\cs_registers_i.pc_if_i[21] ),
    .I1(\cs_registers_i.pc_id_i[21] ),
    .S(net1708),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16910_ (.I0(\cs_registers_i.csr_depc_o[21] ),
    .I1(_03296_),
    .S(_03906_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16911_ (.I0(_03934_),
    .I1(_03935_),
    .S(net1617),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16912_ (.I0(\cs_registers_i.pc_if_i[22] ),
    .I1(\cs_registers_i.pc_id_i[22] ),
    .S(net1708),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16913_ (.I0(\cs_registers_i.csr_depc_o[22] ),
    .I1(_03306_),
    .S(_03906_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16914_ (.I0(_03936_),
    .I1(_03937_),
    .S(_03879_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16915_ (.I0(\cs_registers_i.pc_if_i[23] ),
    .I1(\cs_registers_i.pc_id_i[23] ),
    .S(net1708),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16916_ (.I0(\cs_registers_i.csr_depc_o[23] ),
    .I1(_03321_),
    .S(_03906_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16917_ (.I0(_03938_),
    .I1(_03939_),
    .S(net1617),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16918_ (.I0(\cs_registers_i.pc_if_i[24] ),
    .I1(\cs_registers_i.pc_id_i[24] ),
    .S(net1708),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16919_ (.I0(\cs_registers_i.csr_depc_o[24] ),
    .I1(_03323_),
    .S(_03906_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1437 (.I(net165),
    .Z(net1436));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16921_ (.I0(_03940_),
    .I1(_03941_),
    .S(_03879_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16922_ (.I0(\cs_registers_i.pc_if_i[25] ),
    .I1(\cs_registers_i.pc_id_i[25] ),
    .S(net1708),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16923_ (.I0(\cs_registers_i.csr_depc_o[25] ),
    .I1(_03335_),
    .S(_03906_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16924_ (.I0(_03943_),
    .I1(_03944_),
    .S(_03879_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1436 (.I(net164),
    .Z(net1435));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16926_ (.I0(\cs_registers_i.pc_if_i[26] ),
    .I1(\cs_registers_i.pc_id_i[26] ),
    .S(net1708),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16927_ (.I0(\cs_registers_i.csr_depc_o[26] ),
    .I1(_10735_),
    .S(_03906_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16928_ (.I0(_03946_),
    .I1(_03947_),
    .S(_03879_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16929_ (.I0(\cs_registers_i.pc_if_i[27] ),
    .I1(\cs_registers_i.pc_id_i[27] ),
    .S(net1708),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16930_ (.I0(\cs_registers_i.csr_depc_o[27] ),
    .I1(net1517),
    .S(_03906_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16931_ (.I0(_03948_),
    .I1(_03949_),
    .S(_03879_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16932_ (.I0(\cs_registers_i.pc_if_i[28] ),
    .I1(\cs_registers_i.pc_id_i[28] ),
    .S(net1708),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16933_ (.I0(\cs_registers_i.csr_depc_o[28] ),
    .I1(net1516),
    .S(_03906_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16934_ (.I0(_03950_),
    .I1(_03951_),
    .S(_03879_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16935_ (.I0(\cs_registers_i.pc_if_i[29] ),
    .I1(\cs_registers_i.pc_id_i[29] ),
    .S(net1708),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1435 (.I(_09017_),
    .Z(net1434));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16937_ (.I0(\cs_registers_i.csr_depc_o[29] ),
    .I1(_03365_),
    .S(_03906_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16938_ (.I0(_03952_),
    .I1(_03954_),
    .S(_03879_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16939_ (.I0(\cs_registers_i.pc_if_i[2] ),
    .I1(\cs_registers_i.pc_id_i[2] ),
    .S(net1708),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16940_ (.I0(\cs_registers_i.csr_depc_o[2] ),
    .I1(_10258_),
    .S(net1527),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16941_ (.I0(_03955_),
    .I1(_03956_),
    .S(net1617),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16942_ (.I0(\cs_registers_i.pc_if_i[30] ),
    .I1(\cs_registers_i.pc_id_i[30] ),
    .S(net1708),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16943_ (.I0(\cs_registers_i.csr_depc_o[30] ),
    .I1(_10813_),
    .S(_03906_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16944_ (.I0(_03957_),
    .I1(_03958_),
    .S(net1617),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16945_ (.I0(\cs_registers_i.pc_if_i[31] ),
    .I1(\cs_registers_i.pc_id_i[31] ),
    .S(net1708),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16946_ (.I0(\cs_registers_i.csr_depc_o[31] ),
    .I1(_10846_),
    .S(_03906_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16947_ (.I0(_03959_),
    .I1(_03960_),
    .S(net1617),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16948_ (.I0(\cs_registers_i.pc_if_i[3] ),
    .I1(\cs_registers_i.pc_id_i[3] ),
    .S(net1708),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16949_ (.I0(\cs_registers_i.csr_depc_o[3] ),
    .I1(_10891_),
    .S(_03906_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16950_ (.I0(_03961_),
    .I1(_03962_),
    .S(net1617),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16951_ (.I0(\cs_registers_i.pc_if_i[4] ),
    .I1(\cs_registers_i.pc_id_i[4] ),
    .S(net1708),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16952_ (.I0(\cs_registers_i.csr_depc_o[4] ),
    .I1(_10911_),
    .S(net1527),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16953_ (.I0(_03963_),
    .I1(_03964_),
    .S(net1617),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16954_ (.I0(\cs_registers_i.pc_if_i[5] ),
    .I1(\cs_registers_i.pc_id_i[5] ),
    .S(net1708),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16955_ (.I0(\cs_registers_i.csr_depc_o[5] ),
    .I1(_10940_),
    .S(_03906_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16956_ (.I0(_03965_),
    .I1(_03966_),
    .S(net1617),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16957_ (.I0(\cs_registers_i.pc_if_i[6] ),
    .I1(\cs_registers_i.pc_id_i[6] ),
    .S(net1708),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16958_ (.I0(\cs_registers_i.csr_depc_o[6] ),
    .I1(_10956_),
    .S(_03906_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16959_ (.I0(_03967_),
    .I1(_03968_),
    .S(net1617),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16960_ (.I0(\cs_registers_i.pc_if_i[7] ),
    .I1(\cs_registers_i.pc_id_i[7] ),
    .S(net1708),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16961_ (.I0(\cs_registers_i.csr_depc_o[7] ),
    .I1(_10984_),
    .S(net1527),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16962_ (.I0(_03969_),
    .I1(_03970_),
    .S(_03879_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16963_ (.I0(\cs_registers_i.pc_if_i[8] ),
    .I1(\cs_registers_i.pc_id_i[8] ),
    .S(net1708),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16964_ (.I0(\cs_registers_i.csr_depc_o[8] ),
    .I1(_11009_),
    .S(net1527),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16965_ (.I0(_03971_),
    .I1(_03972_),
    .S(_03879_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16966_ (.I0(\cs_registers_i.pc_if_i[9] ),
    .I1(\cs_registers_i.pc_id_i[9] ),
    .S(net1708),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16967_ (.I0(\cs_registers_i.csr_depc_o[9] ),
    .I1(_11024_),
    .S(net1527),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16968_ (.I0(_03973_),
    .I1(_03974_),
    .S(_03879_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16969_ (.A1(net1535),
    .A2(_10935_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1434 (.I(net166),
    .Z(net1433));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16971_ (.I0(\cs_registers_i.dscratch0_q[0] ),
    .I1(_10225_),
    .S(_03975_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16972_ (.I(\cs_registers_i.dscratch0_q[10] ),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16973_ (.I0(_03977_),
    .I1(_10299_),
    .S(net1526),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _16974_ (.I(_03978_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16975_ (.I0(\cs_registers_i.dscratch0_q[11] ),
    .I1(_10348_),
    .S(_03975_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16976_ (.I0(\cs_registers_i.dscratch0_q[12] ),
    .I1(_11052_),
    .S(_03975_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16977_ (.I0(\cs_registers_i.dscratch0_q[13] ),
    .I1(_11059_),
    .S(net1526),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16978_ (.I0(\cs_registers_i.dscratch0_q[14] ),
    .I1(_11064_),
    .S(net1526),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16979_ (.I0(\cs_registers_i.dscratch0_q[15] ),
    .I1(net1531),
    .S(net1526),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16980_ (.I0(\cs_registers_i.dscratch0_q[16] ),
    .I1(_11077_),
    .S(net1526),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16981_ (.I0(\cs_registers_i.dscratch0_q[17] ),
    .I1(_11089_),
    .S(net1526),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16982_ (.I0(\cs_registers_i.dscratch0_q[18] ),
    .I1(_11104_),
    .S(net1526),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16983_ (.I0(\cs_registers_i.dscratch0_q[19] ),
    .I1(_10587_),
    .S(net1526),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone2105 (.I(net2153),
    .Z(net2104));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16985_ (.I0(\cs_registers_i.dscratch0_q[1] ),
    .I1(_10607_),
    .S(net1526),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16986_ (.I0(\cs_registers_i.dscratch0_q[20] ),
    .I1(_10624_),
    .S(net1526),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16987_ (.I0(\cs_registers_i.dscratch0_q[21] ),
    .I1(_03296_),
    .S(net1526),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16988_ (.I0(\cs_registers_i.dscratch0_q[22] ),
    .I1(_03306_),
    .S(net1526),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16989_ (.I0(\cs_registers_i.dscratch0_q[23] ),
    .I1(_03321_),
    .S(net1526),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16990_ (.I0(\cs_registers_i.dscratch0_q[24] ),
    .I1(_03323_),
    .S(net1526),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16991_ (.I0(\cs_registers_i.dscratch0_q[25] ),
    .I1(_03335_),
    .S(net1526),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16992_ (.I0(\cs_registers_i.dscratch0_q[26] ),
    .I1(_10735_),
    .S(net1526),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16993_ (.I0(\cs_registers_i.dscratch0_q[27] ),
    .I1(net1517),
    .S(net1526),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16994_ (.I0(\cs_registers_i.dscratch0_q[28] ),
    .I1(net1516),
    .S(net1526),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2106 (.I(_08544_),
    .Z(net2105));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16996_ (.I0(\cs_registers_i.dscratch0_q[29] ),
    .I1(_03365_),
    .S(net1526),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16997_ (.I0(\cs_registers_i.dscratch0_q[2] ),
    .I1(_10258_),
    .S(net1526),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16998_ (.I0(\cs_registers_i.dscratch0_q[30] ),
    .I1(_10813_),
    .S(net1526),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _16999_ (.I0(\cs_registers_i.dscratch0_q[31] ),
    .I1(_10846_),
    .S(_03975_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17000_ (.I0(\cs_registers_i.dscratch0_q[3] ),
    .I1(_10891_),
    .S(net1526),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17001_ (.I0(\cs_registers_i.dscratch0_q[4] ),
    .I1(_10911_),
    .S(_03975_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17002_ (.I0(\cs_registers_i.dscratch0_q[5] ),
    .I1(_10940_),
    .S(_03975_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17003_ (.I0(\cs_registers_i.dscratch0_q[6] ),
    .I1(_10956_),
    .S(net1526),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17004_ (.I0(\cs_registers_i.dscratch0_q[7] ),
    .I1(_10984_),
    .S(net1526),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17005_ (.I0(\cs_registers_i.dscratch0_q[8] ),
    .I1(_11009_),
    .S(net1526),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17006_ (.I0(\cs_registers_i.dscratch0_q[9] ),
    .I1(_11024_),
    .S(net1526),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17007_ (.A1(net1535),
    .A2(_10930_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1433 (.I(net168),
    .Z(net1432));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17009_ (.I0(\cs_registers_i.dscratch1_q[0] ),
    .I1(_10225_),
    .S(net1525),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17010_ (.I(\cs_registers_i.dscratch1_q[10] ),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17011_ (.I0(_03983_),
    .I1(_10299_),
    .S(net1525),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17012_ (.I(_03984_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17013_ (.I0(\cs_registers_i.dscratch1_q[11] ),
    .I1(_10348_),
    .S(net1525),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17014_ (.I0(\cs_registers_i.dscratch1_q[12] ),
    .I1(_11052_),
    .S(net1525),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17015_ (.I0(\cs_registers_i.dscratch1_q[13] ),
    .I1(_11059_),
    .S(net1525),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17016_ (.I0(\cs_registers_i.dscratch1_q[14] ),
    .I1(_11064_),
    .S(net1525),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17017_ (.I0(\cs_registers_i.dscratch1_q[15] ),
    .I1(net1531),
    .S(net1525),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17018_ (.I0(\cs_registers_i.dscratch1_q[16] ),
    .I1(_11077_),
    .S(net1525),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17019_ (.I0(\cs_registers_i.dscratch1_q[17] ),
    .I1(_11089_),
    .S(net1525),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17020_ (.I0(\cs_registers_i.dscratch1_q[18] ),
    .I1(_11104_),
    .S(net1525),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17021_ (.I0(\cs_registers_i.dscratch1_q[19] ),
    .I1(_10587_),
    .S(net1525),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2107 (.I(_09485_),
    .Z(net2106));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17023_ (.I0(\cs_registers_i.dscratch1_q[1] ),
    .I1(_10607_),
    .S(net1525),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17024_ (.I0(\cs_registers_i.dscratch1_q[20] ),
    .I1(_10624_),
    .S(net1525),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17025_ (.I0(\cs_registers_i.dscratch1_q[21] ),
    .I1(_03296_),
    .S(net1525),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17026_ (.I0(\cs_registers_i.dscratch1_q[22] ),
    .I1(_03306_),
    .S(net1525),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17027_ (.I0(\cs_registers_i.dscratch1_q[23] ),
    .I1(_03321_),
    .S(net1525),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17028_ (.I0(\cs_registers_i.dscratch1_q[24] ),
    .I1(_03323_),
    .S(net1525),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17029_ (.I0(\cs_registers_i.dscratch1_q[25] ),
    .I1(_03335_),
    .S(net1525),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17030_ (.I0(\cs_registers_i.dscratch1_q[26] ),
    .I1(_10735_),
    .S(net1525),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17031_ (.I0(\cs_registers_i.dscratch1_q[27] ),
    .I1(net1517),
    .S(net1525),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17032_ (.I0(\cs_registers_i.dscratch1_q[28] ),
    .I1(net1516),
    .S(net1525),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1432 (.I(net171),
    .Z(net1431));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17034_ (.I0(\cs_registers_i.dscratch1_q[29] ),
    .I1(_03365_),
    .S(net1525),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17035_ (.I0(\cs_registers_i.dscratch1_q[2] ),
    .I1(_10258_),
    .S(net1525),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17036_ (.I0(\cs_registers_i.dscratch1_q[30] ),
    .I1(_10813_),
    .S(net1525),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17037_ (.I0(\cs_registers_i.dscratch1_q[31] ),
    .I1(_10846_),
    .S(net1525),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17038_ (.I0(\cs_registers_i.dscratch1_q[3] ),
    .I1(_10891_),
    .S(net1525),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17039_ (.I0(\cs_registers_i.dscratch1_q[4] ),
    .I1(_10911_),
    .S(net1525),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17040_ (.I0(\cs_registers_i.dscratch1_q[5] ),
    .I1(_10940_),
    .S(net1525),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17041_ (.I0(\cs_registers_i.dscratch1_q[6] ),
    .I1(_10956_),
    .S(net1525),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17042_ (.I0(\cs_registers_i.dscratch1_q[7] ),
    .I1(_10984_),
    .S(net1525),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17043_ (.I0(\cs_registers_i.dscratch1_q[8] ),
    .I1(_11009_),
    .S(net1525),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17044_ (.I0(\cs_registers_i.dscratch1_q[9] ),
    .I1(_11024_),
    .S(net1525),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _17045_ (.A1(_09922_),
    .A2(_03878_),
    .B(_03881_),
    .C(\cs_registers_i.debug_mode_i ),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17046_ (.A1(\cs_registers_i.nmi_mode_i ),
    .A2(net1746),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17047_ (.A1(net1588),
    .A2(_03988_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2205 (.I(net170),
    .Z(net2204));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1430 (.I(net173),
    .Z(net1429));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17050_ (.A1(_09907_),
    .A2(_09651_),
    .A3(_09900_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1429 (.I(_09309_),
    .Z(net1428));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17052_ (.A1(net1840),
    .A2(net1706),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17053_ (.A1(_09908_),
    .A2(_03438_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17054_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09905_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17055_ (.I0(_09640_),
    .I1(_03996_),
    .S(net1932),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17056_ (.A1(_03995_),
    .A2(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17057_ (.A1(_09524_),
    .A2(_09899_),
    .B(_09917_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17058_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_03999_),
    .A3(_09900_),
    .B(_09996_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17059_ (.A1(_03994_),
    .A2(_03998_),
    .B(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17060_ (.A1(_09988_),
    .A2(_04001_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2108 (.I(_00889_),
    .Z(net2107));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1428 (.I(_04881_),
    .Z(net1427));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17063_ (.A1(\cs_registers_i.mstack_cause_q[0] ),
    .A2(net1707),
    .B1(_04002_),
    .B2(net1588),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17064_ (.A1(_10273_),
    .A2(net1580),
    .B(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17065_ (.A1(_10372_),
    .A2(_10214_),
    .B(net1580),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17066_ (.I0(_04006_),
    .I1(\cs_registers_i.mcause_q[0] ),
    .S(_04007_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17067_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_09917_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1427 (.I(_04883_),
    .Z(net1426));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17069_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(_09651_),
    .B(_04008_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17070_ (.A1(_03998_),
    .A2(_04010_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17071_ (.A1(_04000_),
    .A2(_04011_),
    .B(_10006_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17072_ (.A1(\cs_registers_i.mstack_cause_q[1] ),
    .A2(net1707),
    .B1(_04012_),
    .B2(net1588),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17073_ (.A1(_03653_),
    .A2(net1580),
    .B(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17074_ (.I0(_04014_),
    .I1(\cs_registers_i.mcause_q[1] ),
    .S(_04007_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17075_ (.I(net1588),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2109 (.I(net2172),
    .Z(net2108));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17077_ (.A1(_09925_),
    .A2(_09926_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17078_ (.A1(_09931_),
    .A2(_09932_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17079_ (.I(_09935_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17080_ (.A1(net1835),
    .A2(_10004_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _17081_ (.A1(_04017_),
    .A2(_04018_),
    .B1(_09969_),
    .B2(_04019_),
    .C(_04020_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17082_ (.A1(_09499_),
    .A2(net1706),
    .B1(_04021_),
    .B2(_09945_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17083_ (.A1(\cs_registers_i.mstack_cause_q[2] ),
    .A2(net1707),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17084_ (.I(net1580),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17085_ (.A1(_10258_),
    .A2(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17086_ (.A1(_04015_),
    .A2(_04022_),
    .B(_04023_),
    .C(_04025_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17087_ (.I0(_04026_),
    .I1(\cs_registers_i.mcause_q[2] ),
    .S(_04007_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17088_ (.A1(_10875_),
    .A2(_10890_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17089_ (.A1(net1855),
    .A2(_09996_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17090_ (.A1(net2050),
    .A2(\cs_registers_i.mie_q[15] ),
    .A3(_09929_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17091_ (.A1(_09933_),
    .A2(_10004_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17092_ (.A1(_04029_),
    .A2(_04030_),
    .B(_09945_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17093_ (.A1(_09908_),
    .A2(_03438_),
    .A3(_04028_),
    .B(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17094_ (.A1(\cs_registers_i.mstack_cause_q[3] ),
    .A2(net1707),
    .B1(_04032_),
    .B2(net1588),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17095_ (.A1(_04027_),
    .A2(net1580),
    .B(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17096_ (.I0(_04034_),
    .I1(\cs_registers_i.mcause_q[3] ),
    .S(_04007_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17097_ (.I(_09986_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17098_ (.A1(_09969_),
    .A2(_04035_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17099_ (.A1(_09944_),
    .A2(_04036_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17100_ (.A1(\cs_registers_i.mstack_cause_q[4] ),
    .A2(net1707),
    .B(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17101_ (.A1(_11093_),
    .A2(net1580),
    .B(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17102_ (.I0(_04039_),
    .I1(\cs_registers_i.mcause_q[4] ),
    .S(_04007_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17103_ (.A1(_10846_),
    .A2(_04024_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2110 (.I(_00825_),
    .Z(net2109));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17105_ (.A1(\cs_registers_i.mstack_cause_q[5] ),
    .A2(net1707),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17106_ (.A1(_09945_),
    .A2(_04040_),
    .A3(_04042_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17107_ (.I0(_04043_),
    .I1(\cs_registers_i.mcause_q[5] ),
    .S(_04007_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _17108_ (.A1(net1535),
    .A2(_10923_),
    .B(_03989_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2111 (.I(_07630_),
    .Z(net2110));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17110_ (.A1(\cs_registers_i.mstack_epc_q[0] ),
    .A2(net1707),
    .B1(_04044_),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17111_ (.I(_04046_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone2112 (.I(net2148),
    .Z(net2111));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17113_ (.A1(_03905_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[10] ),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17114_ (.A1(_10299_),
    .A2(net1580),
    .B(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17115_ (.I0(_04049_),
    .I1(\cs_registers_i.csr_mepc_o[10] ),
    .S(_04044_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2113 (.I(net2113),
    .Z(net2112));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17117_ (.A1(_03909_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[11] ),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17118_ (.A1(_03471_),
    .A2(net1580),
    .B(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17119_ (.I0(_04052_),
    .I1(\cs_registers_i.csr_mepc_o[11] ),
    .S(_04044_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17120_ (.A1(_03911_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[12] ),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17121_ (.A1(_10404_),
    .A2(net1580),
    .B(_04053_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17122_ (.I0(_04054_),
    .I1(\cs_registers_i.csr_mepc_o[12] ),
    .S(_04044_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17123_ (.A1(_03913_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[13] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17124_ (.A1(_10448_),
    .A2(net1580),
    .B(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17125_ (.I0(_04056_),
    .I1(\cs_registers_i.csr_mepc_o[13] ),
    .S(net1524),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17126_ (.A1(_03915_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[14] ),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17127_ (.A1(_10472_),
    .A2(net1580),
    .B(_04057_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17128_ (.I0(_04058_),
    .I1(\cs_registers_i.csr_mepc_o[14] ),
    .S(_04044_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17129_ (.I(net1531),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17130_ (.A1(_03917_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[15] ),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17131_ (.A1(_04059_),
    .A2(net1580),
    .B(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17132_ (.I0(_04061_),
    .I1(\cs_registers_i.csr_mepc_o[15] ),
    .S(_04044_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2114 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net2113));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2115 (.I(net2058),
    .Z(net2114));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17135_ (.A1(_03920_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[16] ),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17136_ (.A1(_10525_),
    .A2(net1580),
    .B(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2116 (.I(_07555_),
    .Z(net2115));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17138_ (.I0(_04065_),
    .I1(\cs_registers_i.csr_mepc_o[16] ),
    .S(net1524),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17139_ (.A1(_03922_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[17] ),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17140_ (.A1(_10546_),
    .A2(net1580),
    .B(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17141_ (.I0(_04068_),
    .I1(\cs_registers_i.csr_mepc_o[17] ),
    .S(_04044_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17142_ (.A1(_03924_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[18] ),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17143_ (.A1(_10567_),
    .A2(net1580),
    .B(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17144_ (.I0(_04070_),
    .I1(\cs_registers_i.csr_mepc_o[18] ),
    .S(net1524),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17145_ (.A1(_03927_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[19] ),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17146_ (.A1(_03537_),
    .A2(net1580),
    .B(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17147_ (.I0(_04072_),
    .I1(\cs_registers_i.csr_mepc_o[19] ),
    .S(net1524),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17148_ (.A1(_03929_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[1] ),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17149_ (.A1(_03653_),
    .A2(net1580),
    .B(_04073_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17150_ (.I0(_04074_),
    .I1(\cs_registers_i.csr_mepc_o[1] ),
    .S(_04044_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1426 (.I(_01039_),
    .Z(net1425));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17152_ (.A1(_03932_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[20] ),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17153_ (.A1(_03547_),
    .A2(net1580),
    .B(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17154_ (.I0(_04077_),
    .I1(\cs_registers_i.csr_mepc_o[20] ),
    .S(net1524),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17155_ (.A1(_03934_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[21] ),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17156_ (.A1(_10647_),
    .A2(net1580),
    .B(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17157_ (.I0(_04079_),
    .I1(\cs_registers_i.csr_mepc_o[21] ),
    .S(net1524),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17158_ (.A1(_03936_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[22] ),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17159_ (.A1(_10663_),
    .A2(net1580),
    .B(_04080_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17160_ (.I0(_04081_),
    .I1(\cs_registers_i.csr_mepc_o[22] ),
    .S(net1524),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17161_ (.A1(_03938_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[23] ),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17162_ (.A1(_10678_),
    .A2(net1580),
    .B(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17163_ (.I0(_04083_),
    .I1(\cs_registers_i.csr_mepc_o[23] ),
    .S(net1524),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17164_ (.A1(_03940_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[24] ),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17165_ (.A1(_10698_),
    .A2(net1580),
    .B(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17166_ (.I0(_04085_),
    .I1(\cs_registers_i.csr_mepc_o[24] ),
    .S(net1524),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1425 (.I(_01040_),
    .Z(net1424));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1424 (.I(_01045_),
    .Z(net1423));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17169_ (.A1(_03943_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[25] ),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17170_ (.A1(_10716_),
    .A2(net1580),
    .B(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1423 (.I(_01046_),
    .Z(net1422));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17172_ (.I0(_04089_),
    .I1(\cs_registers_i.csr_mepc_o[25] ),
    .S(net1524),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17173_ (.I(\cs_registers_i.csr_mepc_o[26] ),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17174_ (.A1(_03946_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[26] ),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17175_ (.I(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _17176_ (.A1(_10735_),
    .A2(_04024_),
    .B(net1524),
    .C(_04093_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17177_ (.A1(_04091_),
    .A2(net1524),
    .B(_04094_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17178_ (.I(\cs_registers_i.csr_mepc_o[27] ),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17179_ (.A1(_03948_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[27] ),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17180_ (.I(_04096_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _17181_ (.A1(net1517),
    .A2(_04024_),
    .B(net1524),
    .C(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17182_ (.A1(_04095_),
    .A2(net1524),
    .B(_04098_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17183_ (.I(\cs_registers_i.csr_mepc_o[28] ),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17184_ (.A1(_03950_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[28] ),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17185_ (.I(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _17186_ (.A1(net1516),
    .A2(_04024_),
    .B(net1524),
    .C(_04101_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17187_ (.A1(_04099_),
    .A2(net1524),
    .B(_04102_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17188_ (.A1(_03952_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[29] ),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17189_ (.A1(_10788_),
    .A2(net1580),
    .B(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17190_ (.I0(_04104_),
    .I1(\cs_registers_i.csr_mepc_o[29] ),
    .S(net1524),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17191_ (.A1(_03955_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[2] ),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17192_ (.A1(_04025_),
    .A2(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17193_ (.I0(_04106_),
    .I1(\cs_registers_i.csr_mepc_o[2] ),
    .S(_04044_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _17194_ (.A1(_10800_),
    .A2(_10801_),
    .A3(_10802_),
    .A4(_10809_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17195_ (.A1(net1705),
    .A2(_10811_),
    .B1(_04107_),
    .B2(_01347_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17196_ (.A1(_03957_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[30] ),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17197_ (.A1(_04108_),
    .A2(net1580),
    .B(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17198_ (.I0(_04110_),
    .I1(\cs_registers_i.csr_mepc_o[30] ),
    .S(net1524),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17199_ (.A1(_03959_),
    .A2(net1588),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17200_ (.A1(\cs_registers_i.mstack_epc_q[31] ),
    .A2(net1707),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17201_ (.A1(_04040_),
    .A2(_04111_),
    .A3(_04112_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17202_ (.I0(_04113_),
    .I1(\cs_registers_i.csr_mepc_o[31] ),
    .S(_04044_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17203_ (.A1(_03961_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[3] ),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17204_ (.A1(_04027_),
    .A2(net1580),
    .B(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17205_ (.I0(_04115_),
    .I1(\cs_registers_i.csr_mepc_o[3] ),
    .S(_04044_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17206_ (.A1(_03963_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[4] ),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17207_ (.A1(_11093_),
    .A2(net1580),
    .B(_04116_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17208_ (.I0(_04117_),
    .I1(\cs_registers_i.csr_mepc_o[4] ),
    .S(_04044_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17209_ (.A1(_03965_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[5] ),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17210_ (.A1(_03347_),
    .A2(net1580),
    .B(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17211_ (.I0(_04119_),
    .I1(\cs_registers_i.csr_mepc_o[5] ),
    .S(_04044_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17212_ (.A1(_03967_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[6] ),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17213_ (.A1(_03377_),
    .A2(net1580),
    .B(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17214_ (.I0(_04121_),
    .I1(\cs_registers_i.csr_mepc_o[6] ),
    .S(_04044_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17215_ (.A1(_03969_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[7] ),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17216_ (.A1(_03384_),
    .A2(net1580),
    .B(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17217_ (.I0(_04123_),
    .I1(\cs_registers_i.csr_mepc_o[7] ),
    .S(_04044_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17218_ (.A1(_03971_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[8] ),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17219_ (.A1(_03386_),
    .A2(net1580),
    .B(_04124_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17220_ (.I0(_04125_),
    .I1(\cs_registers_i.csr_mepc_o[8] ),
    .S(_04044_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17221_ (.A1(_11012_),
    .A2(_11023_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17222_ (.A1(_03973_),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_epc_q[9] ),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17223_ (.A1(_04126_),
    .A2(net1580),
    .B(_04127_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17224_ (.I0(_04128_),
    .I1(\cs_registers_i.csr_mepc_o[9] ),
    .S(_04044_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17225_ (.A1(net1701),
    .A2(_07859_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17226_ (.A1(_09588_),
    .A2(_04129_),
    .B(_09577_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17227_ (.A1(_09600_),
    .A2(_04130_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17228_ (.A1(net1535),
    .A2(_04131_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1422 (.I(_01051_),
    .Z(net1421));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1421 (.I(_01052_),
    .Z(net1420));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17231_ (.I0(\cs_registers_i.mie_q[0] ),
    .I1(_11077_),
    .S(_04132_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17232_ (.I0(\cs_registers_i.mie_q[10] ),
    .I1(_10735_),
    .S(_04132_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17233_ (.I0(\cs_registers_i.mie_q[11] ),
    .I1(net1517),
    .S(_04132_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17234_ (.I0(\cs_registers_i.mie_q[12] ),
    .I1(net1516),
    .S(_04132_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17235_ (.I0(\cs_registers_i.mie_q[13] ),
    .I1(_03365_),
    .S(_04132_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17236_ (.I0(\cs_registers_i.mie_q[14] ),
    .I1(_10813_),
    .S(_04132_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17237_ (.I0(\cs_registers_i.mie_q[15] ),
    .I1(_10348_),
    .S(_04132_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17238_ (.I0(\cs_registers_i.mie_q[16] ),
    .I1(_10984_),
    .S(_04132_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17239_ (.I0(\cs_registers_i.mie_q[17] ),
    .I1(_10891_),
    .S(_04132_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17240_ (.I0(\cs_registers_i.mie_q[1] ),
    .I1(_11089_),
    .S(_04132_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17241_ (.I0(\cs_registers_i.mie_q[2] ),
    .I1(_11104_),
    .S(_04132_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17242_ (.I0(\cs_registers_i.mie_q[3] ),
    .I1(_10587_),
    .S(_04132_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17243_ (.I0(\cs_registers_i.mie_q[4] ),
    .I1(_10624_),
    .S(_04132_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17244_ (.I0(\cs_registers_i.mie_q[5] ),
    .I1(_03296_),
    .S(_04132_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17245_ (.I0(\cs_registers_i.mie_q[6] ),
    .I1(_03306_),
    .S(_04132_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17246_ (.I0(\cs_registers_i.mie_q[7] ),
    .I1(_03321_),
    .S(_04132_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17247_ (.I0(\cs_registers_i.mie_q[8] ),
    .I1(_03323_),
    .S(_04132_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17248_ (.I0(\cs_registers_i.mie_q[9] ),
    .I1(_03335_),
    .S(_04132_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17249_ (.A1(net1535),
    .A2(_10925_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2117 (.I(net1690),
    .Z(net2116));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17251_ (.I0(\cs_registers_i.mscratch_q[0] ),
    .I1(_10225_),
    .S(_04135_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17252_ (.I(\cs_registers_i.mscratch_q[10] ),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17253_ (.I0(_04137_),
    .I1(_10299_),
    .S(net1523),
    .Z(_04138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17254_ (.I(_04138_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17255_ (.I0(\cs_registers_i.mscratch_q[11] ),
    .I1(_10348_),
    .S(_04135_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17256_ (.I0(\cs_registers_i.mscratch_q[12] ),
    .I1(_11052_),
    .S(_04135_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17257_ (.I0(\cs_registers_i.mscratch_q[13] ),
    .I1(_11059_),
    .S(_04135_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17258_ (.I0(\cs_registers_i.mscratch_q[14] ),
    .I1(_11064_),
    .S(net1523),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17259_ (.I0(\cs_registers_i.mscratch_q[15] ),
    .I1(net1531),
    .S(_04135_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17260_ (.I0(\cs_registers_i.mscratch_q[16] ),
    .I1(_11077_),
    .S(net1523),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17261_ (.I0(\cs_registers_i.mscratch_q[17] ),
    .I1(_11089_),
    .S(_04135_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17262_ (.I0(\cs_registers_i.mscratch_q[18] ),
    .I1(_11104_),
    .S(net1523),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17263_ (.I0(\cs_registers_i.mscratch_q[19] ),
    .I1(_10587_),
    .S(net1523),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1420 (.I(_01058_),
    .Z(net1419));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17265_ (.I0(\cs_registers_i.mscratch_q[1] ),
    .I1(_10607_),
    .S(_04135_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17266_ (.I0(\cs_registers_i.mscratch_q[20] ),
    .I1(_10624_),
    .S(net1523),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17267_ (.I0(\cs_registers_i.mscratch_q[21] ),
    .I1(_03296_),
    .S(net1523),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17268_ (.I0(\cs_registers_i.mscratch_q[22] ),
    .I1(_03306_),
    .S(net1523),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17269_ (.I0(\cs_registers_i.mscratch_q[23] ),
    .I1(_03321_),
    .S(net1523),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17270_ (.I0(\cs_registers_i.mscratch_q[24] ),
    .I1(_03323_),
    .S(net1523),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17271_ (.I0(\cs_registers_i.mscratch_q[25] ),
    .I1(_03335_),
    .S(net1523),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17272_ (.I0(\cs_registers_i.mscratch_q[26] ),
    .I1(_10735_),
    .S(net1523),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17273_ (.I0(\cs_registers_i.mscratch_q[27] ),
    .I1(net1517),
    .S(net1523),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17274_ (.I0(\cs_registers_i.mscratch_q[28] ),
    .I1(net1516),
    .S(net1523),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1419 (.I(_01063_),
    .Z(net1418));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17276_ (.I0(\cs_registers_i.mscratch_q[29] ),
    .I1(_03365_),
    .S(net1523),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17277_ (.I0(\cs_registers_i.mscratch_q[2] ),
    .I1(_10258_),
    .S(_04135_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17278_ (.I0(\cs_registers_i.mscratch_q[30] ),
    .I1(_10813_),
    .S(net1523),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17279_ (.I0(\cs_registers_i.mscratch_q[31] ),
    .I1(_10846_),
    .S(_04135_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17280_ (.I0(\cs_registers_i.mscratch_q[3] ),
    .I1(_10891_),
    .S(_04135_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17281_ (.I0(\cs_registers_i.mscratch_q[4] ),
    .I1(_10911_),
    .S(_04135_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17282_ (.I0(\cs_registers_i.mscratch_q[5] ),
    .I1(_10940_),
    .S(_04135_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17283_ (.I0(\cs_registers_i.mscratch_q[6] ),
    .I1(_10956_),
    .S(_04135_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17284_ (.I0(\cs_registers_i.mscratch_q[7] ),
    .I1(_10984_),
    .S(_04135_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17285_ (.I0(\cs_registers_i.mscratch_q[8] ),
    .I1(_11009_),
    .S(_04135_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17286_ (.I0(\cs_registers_i.mscratch_q[9] ),
    .I1(_11024_),
    .S(net1523),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1417 (.I(_01069_),
    .Z(net1416));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17288_ (.I0(\cs_registers_i.mstack_cause_q[0] ),
    .I1(\cs_registers_i.mcause_q[0] ),
    .S(net1588),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17289_ (.I0(\cs_registers_i.mstack_cause_q[1] ),
    .I1(\cs_registers_i.mcause_q[1] ),
    .S(net1588),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17290_ (.I0(\cs_registers_i.mstack_cause_q[2] ),
    .I1(\cs_registers_i.mcause_q[2] ),
    .S(net1588),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17291_ (.I0(\cs_registers_i.mstack_cause_q[3] ),
    .I1(\cs_registers_i.mcause_q[3] ),
    .S(net1588),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17292_ (.I0(\cs_registers_i.mstack_cause_q[4] ),
    .I1(\cs_registers_i.mcause_q[4] ),
    .S(net1588),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17293_ (.I0(\cs_registers_i.mstack_cause_q[5] ),
    .I1(\cs_registers_i.mcause_q[5] ),
    .S(net1588),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17294_ (.I0(\cs_registers_i.mstack_q[0] ),
    .I1(\cs_registers_i.mstatus_q[2] ),
    .S(net1588),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1416 (.I(_01070_),
    .Z(net1415));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17296_ (.I0(\cs_registers_i.mstack_q[1] ),
    .I1(\cs_registers_i.mstatus_q[3] ),
    .S(net1588),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17297_ (.I0(\cs_registers_i.mstack_q[2] ),
    .I1(\cs_registers_i.mstatus_q[4] ),
    .S(net1588),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17298_ (.I0(\cs_registers_i.mstack_epc_q[0] ),
    .I1(\cs_registers_i.csr_mepc_o[0] ),
    .S(net1588),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17299_ (.I0(\cs_registers_i.mstack_epc_q[10] ),
    .I1(\cs_registers_i.csr_mepc_o[10] ),
    .S(net1588),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17300_ (.I0(\cs_registers_i.mstack_epc_q[11] ),
    .I1(\cs_registers_i.csr_mepc_o[11] ),
    .S(net1588),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17301_ (.I0(\cs_registers_i.mstack_epc_q[12] ),
    .I1(\cs_registers_i.csr_mepc_o[12] ),
    .S(net1588),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17302_ (.I0(\cs_registers_i.mstack_epc_q[13] ),
    .I1(\cs_registers_i.csr_mepc_o[13] ),
    .S(net1588),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17303_ (.I0(\cs_registers_i.mstack_epc_q[14] ),
    .I1(\cs_registers_i.csr_mepc_o[14] ),
    .S(net1588),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17304_ (.I0(\cs_registers_i.mstack_epc_q[15] ),
    .I1(\cs_registers_i.csr_mepc_o[15] ),
    .S(net1588),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17305_ (.I0(\cs_registers_i.mstack_epc_q[16] ),
    .I1(\cs_registers_i.csr_mepc_o[16] ),
    .S(net1588),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1415 (.I(_01076_),
    .Z(net1414));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17307_ (.I0(\cs_registers_i.mstack_epc_q[17] ),
    .I1(\cs_registers_i.csr_mepc_o[17] ),
    .S(net1588),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17308_ (.I0(\cs_registers_i.mstack_epc_q[18] ),
    .I1(\cs_registers_i.csr_mepc_o[18] ),
    .S(net1588),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17309_ (.I0(\cs_registers_i.mstack_epc_q[19] ),
    .I1(\cs_registers_i.csr_mepc_o[19] ),
    .S(net1588),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17310_ (.I0(\cs_registers_i.mstack_epc_q[1] ),
    .I1(\cs_registers_i.csr_mepc_o[1] ),
    .S(net1588),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17311_ (.I0(\cs_registers_i.mstack_epc_q[20] ),
    .I1(\cs_registers_i.csr_mepc_o[20] ),
    .S(net1588),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17312_ (.I0(\cs_registers_i.mstack_epc_q[21] ),
    .I1(\cs_registers_i.csr_mepc_o[21] ),
    .S(net1588),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17313_ (.I0(\cs_registers_i.mstack_epc_q[22] ),
    .I1(\cs_registers_i.csr_mepc_o[22] ),
    .S(net1588),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17314_ (.I0(\cs_registers_i.mstack_epc_q[23] ),
    .I1(\cs_registers_i.csr_mepc_o[23] ),
    .S(net1588),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17315_ (.I0(\cs_registers_i.mstack_epc_q[24] ),
    .I1(\cs_registers_i.csr_mepc_o[24] ),
    .S(net1588),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17316_ (.I0(\cs_registers_i.mstack_epc_q[25] ),
    .I1(\cs_registers_i.csr_mepc_o[25] ),
    .S(net1588),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1418 (.I(_01064_),
    .Z(net1417));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17318_ (.I0(\cs_registers_i.mstack_epc_q[26] ),
    .I1(\cs_registers_i.csr_mepc_o[26] ),
    .S(net1588),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17319_ (.I0(\cs_registers_i.mstack_epc_q[27] ),
    .I1(\cs_registers_i.csr_mepc_o[27] ),
    .S(net1588),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17320_ (.I0(\cs_registers_i.mstack_epc_q[28] ),
    .I1(\cs_registers_i.csr_mepc_o[28] ),
    .S(net1588),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17321_ (.I0(\cs_registers_i.mstack_epc_q[29] ),
    .I1(\cs_registers_i.csr_mepc_o[29] ),
    .S(net1588),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17322_ (.I0(\cs_registers_i.mstack_epc_q[2] ),
    .I1(\cs_registers_i.csr_mepc_o[2] ),
    .S(net1588),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17323_ (.I0(\cs_registers_i.mstack_epc_q[30] ),
    .I1(\cs_registers_i.csr_mepc_o[30] ),
    .S(net1588),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17324_ (.I0(\cs_registers_i.mstack_epc_q[31] ),
    .I1(\cs_registers_i.csr_mepc_o[31] ),
    .S(net1588),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17325_ (.I0(\cs_registers_i.mstack_epc_q[3] ),
    .I1(\cs_registers_i.csr_mepc_o[3] ),
    .S(net1588),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17326_ (.I0(\cs_registers_i.mstack_epc_q[4] ),
    .I1(\cs_registers_i.csr_mepc_o[4] ),
    .S(net1588),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17327_ (.I0(\cs_registers_i.mstack_epc_q[5] ),
    .I1(\cs_registers_i.csr_mepc_o[5] ),
    .S(net1588),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1414 (.I(_01094_),
    .Z(net1413));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17329_ (.I0(\cs_registers_i.mstack_epc_q[6] ),
    .I1(\cs_registers_i.csr_mepc_o[6] ),
    .S(net1588),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17330_ (.I0(\cs_registers_i.mstack_epc_q[7] ),
    .I1(\cs_registers_i.csr_mepc_o[7] ),
    .S(net1588),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17331_ (.I0(\cs_registers_i.mstack_epc_q[8] ),
    .I1(\cs_registers_i.csr_mepc_o[8] ),
    .S(net1588),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17332_ (.I0(\cs_registers_i.mstack_epc_q[9] ),
    .I1(\cs_registers_i.csr_mepc_o[9] ),
    .S(net1588),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17333_ (.A1(_10372_),
    .A2(_10535_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17334_ (.I0(\cs_registers_i.csr_mstatus_tw_o ),
    .I1(_03296_),
    .S(_04146_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17335_ (.I0(\cs_registers_i.mstatus_q[1] ),
    .I1(_11089_),
    .S(_04146_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1413 (.I(_01099_),
    .Z(net1412));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2118 (.I(_07629_),
    .Z(net2117));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17338_ (.I0(\id_stage_i.controller_i.instr_i[0] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17339_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04149_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17340_ (.A1(_09907_),
    .A2(_03994_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17341_ (.A1(_09942_),
    .A2(_09996_),
    .A3(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17342_ (.A1(_10273_),
    .A2(net1588),
    .B1(_04150_),
    .B2(net1579),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17343_ (.A1(net1535),
    .A2(_10927_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17344_ (.A1(_04015_),
    .A2(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2119 (.I(_07831_),
    .Z(net2118));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17346_ (.I0(\cs_registers_i.mtval_q[0] ),
    .I1(_04153_),
    .S(_04155_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 clone2120 (.A1(net2120),
    .A2(_08215_),
    .B(_08217_),
    .ZN(net2119));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17348_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17349_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(\cs_registers_i.pc_id_i[5] ),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17350_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A4(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17351_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .A3(\cs_registers_i.pc_id_i[8] ),
    .A4(\cs_registers_i.pc_id_i[9] ),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17352_ (.A1(_04160_),
    .A2(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17353_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1412 (.I(_01118_),
    .Z(net1411));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17355_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04158_),
    .C1(_04163_),
    .C2(net1840),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17356_ (.A1(_10299_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17357_ (.I0(\cs_registers_i.mtval_q[10] ),
    .I1(_04166_),
    .S(_04155_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2121 (.I(_08216_),
    .Z(net2120));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17359_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17360_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(\cs_registers_i.pc_id_i[4] ),
    .A3(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A4(_00960_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17361_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_04169_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17362_ (.A1(\cs_registers_i.pc_id_i[10] ),
    .A2(_04161_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17363_ (.A1(_04170_),
    .A2(_04171_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17364_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_04172_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17365_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04168_),
    .C1(_04173_),
    .C2(net1840),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17366_ (.A1(_03471_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17367_ (.I0(\cs_registers_i.mtval_q[11] ),
    .I1(_04175_),
    .S(_04155_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17368_ (.I0(net2021),
    .I1(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17369_ (.A1(_04160_),
    .A2(_04171_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17370_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_04177_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17371_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_04178_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17372_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04176_),
    .C1(_04179_),
    .C2(net1840),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17373_ (.A1(_10404_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04180_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17374_ (.I0(\cs_registers_i.mtval_q[12] ),
    .I1(_04181_),
    .S(_04155_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17375_ (.I0(\id_stage_i.controller_i.instr_i[13] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17376_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[11] ),
    .A3(_04172_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17377_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_04183_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17378_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04182_),
    .C1(_04184_),
    .C2(net1840),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17379_ (.A1(_10448_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17380_ (.I0(\cs_registers_i.mtval_q[13] ),
    .I1(_04186_),
    .S(_04155_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2122 (.I(_08216_),
    .Z(net2121));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17382_ (.I0(\id_stage_i.controller_i.instr_i[14] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17383_ (.I(\cs_registers_i.pc_id_i[14] ),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17384_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[11] ),
    .A3(\cs_registers_i.pc_id_i[13] ),
    .A4(_04177_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17385_ (.A1(_04189_),
    .A2(_04190_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1411 (.I(net167),
    .Z(net1410));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17387_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04188_),
    .C1(_04191_),
    .C2(net1840),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17388_ (.A1(_10472_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17389_ (.I0(\cs_registers_i.mtval_q[14] ),
    .I1(_04194_),
    .S(net1514),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2123 (.I(net1406),
    .Z(net2122));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17391_ (.I0(net2017),
    .I1(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17392_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(\cs_registers_i.pc_id_i[11] ),
    .A3(\cs_registers_i.pc_id_i[13] ),
    .A4(_04172_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17393_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17394_ (.A1(\cs_registers_i.pc_id_i[15] ),
    .A2(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17395_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04196_),
    .C1(_04199_),
    .C2(net1840),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17396_ (.A1(_04059_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04200_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2124 (.I(_08504_),
    .Z(net2123));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17398_ (.I0(\cs_registers_i.mtval_q[15] ),
    .I1(_04201_),
    .S(_04155_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1410 (.I(net172),
    .Z(net1409));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17400_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .A3(_04190_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17401_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(_04204_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2125 (.I(_08391_),
    .Z(net2124));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17403_ (.I(\id_stage_i.controller_i.instr_is_compressed_i ),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17404_ (.A1(_04207_),
    .A2(_04008_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1409 (.I(net2169),
    .Z(net1408));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17406_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net1706),
    .B1(_04205_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1965),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17407_ (.A1(_10525_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17408_ (.I0(\cs_registers_i.mtval_q[16] ),
    .I1(_04211_),
    .S(net1514),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17409_ (.I(\cs_registers_i.pc_id_i[17] ),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17410_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .A3(\cs_registers_i.pc_id_i[16] ),
    .A4(_04197_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17411_ (.A1(_04212_),
    .A2(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17412_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net1706),
    .B1(_04214_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1962),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17413_ (.A1(_10546_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17414_ (.I0(\cs_registers_i.mtval_q[17] ),
    .I1(_04216_),
    .S(net1514),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17415_ (.I(\cs_registers_i.pc_id_i[18] ),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17416_ (.A1(\cs_registers_i.pc_id_i[14] ),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .A3(\cs_registers_i.pc_id_i[16] ),
    .A4(\cs_registers_i.pc_id_i[17] ),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17417_ (.A1(_04190_),
    .A2(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17418_ (.A1(_04217_),
    .A2(_04219_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17419_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net1706),
    .B1(_04220_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1960),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17420_ (.A1(_10567_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17421_ (.I0(\cs_registers_i.mtval_q[18] ),
    .I1(_04222_),
    .S(net1514),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17422_ (.A1(\cs_registers_i.pc_id_i[18] ),
    .A2(_04218_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17423_ (.A1(_04197_),
    .A2(_04223_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17424_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17425_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net1706),
    .B1(_04225_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1958),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17426_ (.A1(_03537_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04226_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17427_ (.I0(\cs_registers_i.mtval_q[19] ),
    .I1(_04227_),
    .S(net1514),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17428_ (.I0(\id_stage_i.controller_i.instr_i[1] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17429_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_04229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17430_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04228_),
    .C1(_04229_),
    .C2(net1840),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17431_ (.A1(_03653_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17432_ (.I0(\cs_registers_i.mtval_q[1] ),
    .I1(_04231_),
    .S(_04155_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17433_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(_04223_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17434_ (.A1(_04190_),
    .A2(_04232_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17435_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(_04233_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17436_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net1706),
    .B1(_04234_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1932),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17437_ (.A1(_03547_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17438_ (.I0(\cs_registers_i.mtval_q[20] ),
    .I1(_04236_),
    .S(net1514),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17439_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(_04197_),
    .A3(_04232_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17440_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(_04237_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17441_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net1706),
    .B1(_04238_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1908),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17442_ (.A1(_10647_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04239_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17443_ (.I0(\cs_registers_i.mtval_q[21] ),
    .I1(_04240_),
    .S(_04155_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17444_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17445_ (.A1(_04233_),
    .A2(_04241_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17446_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(_04242_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17447_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net1706),
    .B1(_04243_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1903),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17448_ (.A1(_10663_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04244_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17449_ (.I0(\cs_registers_i.mtval_q[22] ),
    .I1(_04245_),
    .S(net1514),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1408 (.I(net174),
    .Z(net1407));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17451_ (.I(\cs_registers_i.pc_id_i[23] ),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17452_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(_04197_),
    .A3(_04232_),
    .A4(_04241_),
    .Z(_04248_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17453_ (.A1(_04247_),
    .A2(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17454_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net1706),
    .B1(_04249_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1900),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17455_ (.A1(_10678_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04250_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17456_ (.I0(\cs_registers_i.mtval_q[23] ),
    .I1(_04251_),
    .S(net1514),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2126 (.I(net2124),
    .Z(net2125));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17458_ (.I(\cs_registers_i.pc_id_i[24] ),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17459_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(_04233_),
    .A3(_04241_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17460_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(_04254_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17461_ (.A1(_04253_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17462_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net1706),
    .B1(_04256_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1899),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17463_ (.A1(_10698_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2127 (.I(_07603_),
    .Z(net2126));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17465_ (.I0(\cs_registers_i.mtval_q[24] ),
    .I1(_04258_),
    .S(net1514),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1406 (.I(_04922_),
    .Z(net1405));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17467_ (.I(\cs_registers_i.pc_id_i[25] ),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17468_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(\cs_registers_i.pc_id_i[24] ),
    .A3(_04248_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17469_ (.A1(_04261_),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17470_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net1706),
    .B1(_04263_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1898),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17471_ (.A1(_10716_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17472_ (.I0(\cs_registers_i.mtval_q[25] ),
    .I1(_04265_),
    .S(net1514),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17473_ (.I(\cs_registers_i.pc_id_i[26] ),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17474_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(\cs_registers_i.pc_id_i[24] ),
    .A3(\cs_registers_i.pc_id_i[25] ),
    .A4(_04254_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17475_ (.A1(_04266_),
    .A2(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17476_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net1706),
    .B1(_04268_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1897),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _17477_ (.A1(_10721_),
    .A2(_10734_),
    .A3(_04015_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17478_ (.A1(net1579),
    .A2(_04269_),
    .B(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17479_ (.I0(\cs_registers_i.mtval_q[26] ),
    .I1(_04271_),
    .S(net1514),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17480_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(\cs_registers_i.pc_id_i[24] ),
    .A3(\cs_registers_i.pc_id_i[25] ),
    .A4(\cs_registers_i.pc_id_i[26] ),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17481_ (.A1(_04248_),
    .A2(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17482_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17483_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net1706),
    .B1(_04274_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1896),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17484_ (.A1(net1579),
    .A2(_04275_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17485_ (.A1(net1517),
    .A2(_04015_),
    .B(_04276_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17486_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(net1514),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17487_ (.A1(net1514),
    .A2(_04277_),
    .B(_04278_),
    .ZN(_01774_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17488_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(_04272_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17489_ (.A1(_04254_),
    .A2(_04279_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17490_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_04280_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17491_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net1706),
    .B1(_04281_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1895),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17492_ (.A1(net1579),
    .A2(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17493_ (.A1(net1516),
    .A2(_04015_),
    .B(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17494_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(net1514),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17495_ (.A1(net1514),
    .A2(_04284_),
    .B(_04285_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17496_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(_04279_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17497_ (.A1(_04248_),
    .A2(_04286_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17498_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17499_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net1706),
    .B1(_04288_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1894),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17500_ (.A1(_10788_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04289_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17501_ (.I0(\cs_registers_i.mtval_q[29] ),
    .I1(_04290_),
    .S(net1514),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17502_ (.I0(net2145),
    .I1(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17503_ (.I0(\cs_registers_i.pc_id_i[2] ),
    .I1(_00961_),
    .S(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17504_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04291_),
    .C1(_04292_),
    .C2(net1840),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17505_ (.A1(_10792_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17506_ (.I0(\cs_registers_i.mtval_q[2] ),
    .I1(_04294_),
    .S(_04155_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17507_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(_04286_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17508_ (.A1(_04254_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17509_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(_04296_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17510_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net1706),
    .B1(_04297_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1892),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17511_ (.A1(_04108_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17512_ (.I0(\cs_registers_i.mtval_q[30] ),
    .I1(_04299_),
    .S(net1514),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17513_ (.A1(_09470_),
    .A2(_10843_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17514_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(_04248_),
    .A3(_04295_),
    .Z(_04301_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17515_ (.A1(\cs_registers_i.pc_id_i[31] ),
    .A2(_04301_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17516_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net1706),
    .B1(_04302_),
    .B2(net1840),
    .C1(_04208_),
    .C2(net1891),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _17517_ (.A1(_10845_),
    .A2(_04300_),
    .A3(net1588),
    .B1(net1579),
    .B2(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17518_ (.I0(\cs_registers_i.mtval_q[31] ),
    .I1(_04304_),
    .S(_04155_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17519_ (.I0(net2131),
    .I1(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17520_ (.A1(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A2(_00960_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17521_ (.A1(\cs_registers_i.pc_id_i[3] ),
    .A2(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17522_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04305_),
    .C1(_04307_),
    .C2(net1840),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17523_ (.A1(_04027_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17524_ (.I0(\cs_registers_i.mtval_q[3] ),
    .I1(_04309_),
    .S(_04155_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17525_ (.I0(net2189),
    .I1(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17526_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(\cs_registers_i.pc_id_i[2] ),
    .A3(\cs_registers_i.pc_id_i[3] ),
    .A4(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17527_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_04311_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17528_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04310_),
    .C1(_04312_),
    .C2(net1840),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17529_ (.A1(_11093_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17530_ (.I0(\cs_registers_i.mtval_q[4] ),
    .I1(_04314_),
    .S(_04155_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17531_ (.I0(\id_stage_i.controller_i.instr_i[5] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17532_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_04169_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17533_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04315_),
    .C1(_04316_),
    .C2(net1840),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17534_ (.A1(_03347_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17535_ (.I0(\cs_registers_i.mtval_q[5] ),
    .I1(_04318_),
    .S(_04155_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17536_ (.I0(net2146),
    .I1(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17537_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_04160_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17538_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04319_),
    .C1(_04320_),
    .C2(net1840),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17539_ (.A1(_03377_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17540_ (.I0(\cs_registers_i.mtval_q[6] ),
    .I1(_04322_),
    .S(_04155_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17541_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17542_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(_04170_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17543_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_04324_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17544_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04323_),
    .C1(_04325_),
    .C2(net1840),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17545_ (.A1(_03384_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04326_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17546_ (.I0(\cs_registers_i.mtval_q[7] ),
    .I1(_04327_),
    .S(_04155_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17547_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17548_ (.I(\cs_registers_i.pc_id_i[8] ),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17549_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .A3(_04160_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17550_ (.A1(_04329_),
    .A2(_04330_),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17551_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04328_),
    .C1(_04331_),
    .C2(net1840),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17552_ (.A1(_03386_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17553_ (.I0(\cs_registers_i.mtval_q[8] ),
    .I1(_04333_),
    .S(_04155_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17554_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .I1(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17555_ (.A1(\cs_registers_i.pc_id_i[6] ),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .A3(\cs_registers_i.pc_id_i[8] ),
    .A4(_04170_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17556_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(_04335_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _17557_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(net1706),
    .B1(_04008_),
    .B2(_04334_),
    .C1(_04336_),
    .C2(net1840),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17558_ (.A1(_04126_),
    .A2(net1588),
    .B1(net1579),
    .B2(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17559_ (.I0(\cs_registers_i.mtval_q[9] ),
    .I1(_04338_),
    .S(_04155_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _17560_ (.A1(_07773_),
    .A2(_10194_),
    .A3(_09599_),
    .A4(_04130_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17561_ (.A1(net1535),
    .A2(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1407 (.I(net177),
    .Z(net1406));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17563_ (.A1(_09498_),
    .A2(_09921_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17564_ (.A1(_10372_),
    .A2(net1557),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17565_ (.A1(net1807),
    .A2(_04343_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2128 (.I(_07603_),
    .Z(net2127));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17567_ (.I(\cs_registers_i.csr_mtvec_o[10] ),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1405 (.I(_05206_),
    .Z(net1404));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17569_ (.A1(net6),
    .A2(net1807),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17570_ (.A1(_10299_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04346_),
    .C(_04348_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1404 (.I(_05207_),
    .Z(net1403));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1403 (.I(net2491),
    .Z(net1402));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 clone2129 (.I(net2058),
    .Z(net2128));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17574_ (.A1(net7),
    .A2(net1807),
    .B1(_04343_),
    .B2(_10348_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17575_ (.A1(_10319_),
    .A2(_04344_),
    .B(_04352_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17576_ (.A1(net8),
    .A2(net1807),
    .B1(_04343_),
    .B2(_11052_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17577_ (.A1(_10382_),
    .A2(_04344_),
    .B(_04353_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17578_ (.I(\cs_registers_i.csr_mtvec_o[13] ),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17579_ (.A1(net9),
    .A2(net1807),
    .B1(_04343_),
    .B2(_11059_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17580_ (.A1(_04354_),
    .A2(_04344_),
    .B(_04355_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17581_ (.I(\cs_registers_i.csr_mtvec_o[14] ),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17582_ (.A1(net10),
    .A2(net1807),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17583_ (.A1(_10472_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04356_),
    .C(_04357_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17584_ (.I(\cs_registers_i.csr_mtvec_o[15] ),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17585_ (.A1(net11),
    .A2(net1807),
    .B1(_04343_),
    .B2(net1531),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17586_ (.A1(_04358_),
    .A2(_04344_),
    .B(_04359_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17587_ (.I(\cs_registers_i.csr_mtvec_o[16] ),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17588_ (.A1(net12),
    .A2(net1807),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17589_ (.A1(_10525_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04360_),
    .C(_04361_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17590_ (.I(\cs_registers_i.csr_mtvec_o[17] ),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17591_ (.A1(net13),
    .A2(net1807),
    .B1(_04343_),
    .B2(_11089_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17592_ (.A1(_04362_),
    .A2(_04344_),
    .B(_04363_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17593_ (.I(\cs_registers_i.csr_mtvec_o[18] ),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17594_ (.A1(net14),
    .A2(net1807),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17595_ (.A1(_10567_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04364_),
    .C(_04365_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17596_ (.I(\cs_registers_i.csr_mtvec_o[19] ),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17597_ (.A1(net15),
    .A2(net1807),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17598_ (.A1(_03537_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04366_),
    .C(_04367_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17599_ (.I(\cs_registers_i.csr_mtvec_o[20] ),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17600_ (.A1(net16),
    .A2(net1807),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17601_ (.A1(_03547_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04368_),
    .C(_04369_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17602_ (.I(\cs_registers_i.csr_mtvec_o[21] ),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17603_ (.A1(net17),
    .A2(net1807),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17604_ (.A1(_10647_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04370_),
    .C(_04371_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17605_ (.I(\cs_registers_i.csr_mtvec_o[22] ),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17606_ (.A1(net18),
    .A2(net1807),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17607_ (.A1(_10663_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04372_),
    .C(_04373_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17608_ (.I(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17609_ (.A1(net19),
    .A2(net1807),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17610_ (.A1(_10678_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04374_),
    .C(_04375_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17611_ (.I(\cs_registers_i.csr_mtvec_o[24] ),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17612_ (.A1(net20),
    .A2(net1807),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17613_ (.A1(_10698_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04376_),
    .C(_04377_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17614_ (.I(\cs_registers_i.csr_mtvec_o[25] ),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17615_ (.A1(net21),
    .A2(net1807),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17616_ (.A1(_10716_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04378_),
    .C(_04379_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17617_ (.I(\cs_registers_i.csr_mtvec_o[26] ),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17618_ (.A1(net22),
    .A2(net1807),
    .B1(_04343_),
    .B2(_10735_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17619_ (.A1(_04380_),
    .A2(_04344_),
    .B(_04381_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17620_ (.I(\cs_registers_i.csr_mtvec_o[27] ),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17621_ (.A1(net23),
    .A2(net1807),
    .B1(_04343_),
    .B2(net1517),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17622_ (.A1(_04382_),
    .A2(_04344_),
    .B(_04383_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17623_ (.I(\cs_registers_i.csr_mtvec_o[28] ),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17624_ (.A1(net24),
    .A2(net1807),
    .B1(_04343_),
    .B2(net1516),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17625_ (.A1(_04384_),
    .A2(_04344_),
    .B(_04385_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17626_ (.I(\cs_registers_i.csr_mtvec_o[29] ),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17627_ (.A1(net25),
    .A2(net1807),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17628_ (.A1(_10788_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04386_),
    .C(_04387_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17629_ (.I(\cs_registers_i.csr_mtvec_o[30] ),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17630_ (.A1(net26),
    .A2(net1807),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17631_ (.A1(_04108_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04388_),
    .C(_04389_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17632_ (.I(\cs_registers_i.csr_mtvec_o[31] ),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17633_ (.A1(net27),
    .A2(net1807),
    .B1(_04343_),
    .B2(_10846_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17634_ (.A1(_04390_),
    .A2(_04344_),
    .B(_04391_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17635_ (.I(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _17636_ (.A1(net28),
    .A2(net1807),
    .B1(_04343_),
    .B2(_11009_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17637_ (.A1(_04392_),
    .A2(_04344_),
    .B(_04393_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17638_ (.I(\cs_registers_i.csr_mtvec_o[9] ),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17639_ (.A1(net29),
    .A2(net1807),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17640_ (.A1(_04126_),
    .A2(_04340_),
    .B1(_04344_),
    .B2(_04394_),
    .C(_04395_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2130 (.I(_09191_),
    .Z(net2129));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17642_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(net1673),
    .A3(_09700_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17643_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .I1(_09740_),
    .S(_04397_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _17644_ (.A1(net2028),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17645_ (.A1(_09700_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17646_ (.I0(_09700_),
    .I1(_04399_),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17647_ (.A1(_00965_),
    .A2(_04398_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17648_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .I1(_04400_),
    .S(_09700_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17649_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_00966_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17650_ (.A1(_04398_),
    .A2(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17651_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .I1(_04402_),
    .S(_09700_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17652_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17653_ (.A1(_09695_),
    .A2(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17654_ (.A1(_04398_),
    .A2(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17655_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .I1(_04405_),
    .S(_09700_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17656_ (.I(_00966_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17657_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A3(_04406_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17658_ (.A1(_04398_),
    .A2(_04407_),
    .B(_10138_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17659_ (.A1(_04399_),
    .A2(_04407_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17660_ (.I0(_04408_),
    .I1(_04409_),
    .S(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17661_ (.I0(\alu_adder_result_ex[0] ),
    .I1(net1784),
    .S(net1674),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17662_ (.A1(net2028),
    .A2(_09700_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2131 (.I(net1890),
    .Z(net2130));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17664_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .I1(_04410_),
    .S(net1543),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17665_ (.I(net1735),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2132 (.I(net2130),
    .Z(net2131));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17667_ (.I0(_04413_),
    .I1(net1451),
    .S(net1596),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17668_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .I1(_04415_),
    .S(net1543),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17669_ (.I(net1738),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17670_ (.I0(_04416_),
    .I1(net1457),
    .S(net1596),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17671_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .I1(_04417_),
    .S(net1543),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17672_ (.I0(_09830_),
    .I1(net2298),
    .S(net1596),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17673_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .I1(_04418_),
    .S(net1543),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17674_ (.A1(net1813),
    .A2(_08605_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17675_ (.I0(_04419_),
    .I1(net1450),
    .S(net1596),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17676_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .I1(_04420_),
    .S(net1543),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17677_ (.A1(net2292),
    .A2(net1596),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17678_ (.A1(net1733),
    .A2(net1596),
    .B(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17679_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .I1(_04422_),
    .S(net1543),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17680_ (.I0(net1748),
    .I1(net1448),
    .S(net1596),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17681_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .I1(_04423_),
    .S(net1543),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17682_ (.I(net1770),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17683_ (.I0(_04424_),
    .I1(net1446),
    .S(net1596),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17684_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .I1(_04425_),
    .S(net1543),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17685_ (.I(net2288),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17686_ (.I0(net1732),
    .I1(_04426_),
    .S(net1596),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17687_ (.I(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17688_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .I1(_04428_),
    .S(net1543),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17689_ (.I0(net1731),
    .I1(net2171),
    .S(net1596),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17690_ (.I(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17691_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .I1(_04430_),
    .S(net1543),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17692_ (.I(net1730),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2133 (.I(net2130),
    .Z(net2132));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17694_ (.I0(_04431_),
    .I1(net1436),
    .S(net1596),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2134 (.I(net1890),
    .Z(net2133));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17696_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .I1(_04433_),
    .S(net1543),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17697_ (.I(net1786),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17698_ (.I0(net1539),
    .I1(_04435_),
    .S(net1674),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17699_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .I1(_04436_),
    .S(net1543),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17700_ (.I0(net1658),
    .I1(net2278),
    .S(net1596),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17701_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .I1(_04437_),
    .S(net1543),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17702_ (.I(net1727),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17703_ (.I0(_04438_),
    .I1(net1410),
    .S(net1596),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17704_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .I1(_04439_),
    .S(net1543),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17705_ (.I(net1726),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17706_ (.I0(_04440_),
    .I1(net1432),
    .S(net1596),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17707_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .I1(_04441_),
    .S(net1543),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17708_ (.I(net169),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17709_ (.I0(net1725),
    .I1(_04442_),
    .S(net1596),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17710_ (.I(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17711_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .I1(_04444_),
    .S(net1543),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17712_ (.I(net2065),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17713_ (.I0(net1723),
    .I1(_04445_),
    .S(net1596),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17714_ (.I(_04446_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17715_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .I1(_04447_),
    .S(net1543),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17716_ (.A1(net1431),
    .A2(net1596),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17717_ (.A1(net1722),
    .A2(net1596),
    .B(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17718_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .I1(_04449_),
    .S(net1543),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17719_ (.I0(net1721),
    .I1(net2293),
    .S(net1596),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17720_ (.I(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17721_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .I1(_04451_),
    .S(net1543),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17722_ (.I(net1720),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17723_ (.I0(_04452_),
    .I1(net1429),
    .S(net1596),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17724_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .I1(_04453_),
    .S(net1543),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17725_ (.I0(net1712),
    .I1(net2138),
    .S(net1596),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2135 (.I(net2093),
    .Z(net2134));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17727_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .I1(_04454_),
    .S(net1543),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17728_ (.I(net1754),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17729_ (.I0(_04456_),
    .I1(net1408),
    .S(net1596),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17730_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .I1(_04457_),
    .S(net1543),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17731_ (.I(net1781),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17732_ (.I0(_04458_),
    .I1(net1521),
    .S(net1596),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17733_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .I1(_04459_),
    .S(net1543),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17734_ (.I(net1752),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17735_ (.I0(_04460_),
    .I1(net2122),
    .S(net1596),
    .Z(_04461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17736_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .I1(_04461_),
    .S(net1543),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17737_ (.I(net2051),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17738_ (.A1(_04462_),
    .A2(_09673_),
    .B(_09467_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17739_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .I1(_04463_),
    .S(net1543),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17740_ (.I(net1780),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17741_ (.I0(net1519),
    .I1(_04464_),
    .S(net1674),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17742_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .I1(_04465_),
    .S(net1543),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17743_ (.I0(net1715),
    .I1(net1454),
    .S(net1596),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17744_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .I1(_04466_),
    .S(net1543),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17745_ (.I0(_08324_),
    .I1(_08337_),
    .S(net1867),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17746_ (.I0(_04467_),
    .I1(_08334_),
    .S(net1844),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17747_ (.I0(net1499),
    .I1(_04468_),
    .S(net1674),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17748_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .I1(_04469_),
    .S(net1543),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17749_ (.I0(_08348_),
    .I1(_08359_),
    .S(net1867),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17750_ (.I0(_04470_),
    .I1(_08356_),
    .S(net1844),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17751_ (.I0(_04471_),
    .I1(net1500),
    .S(net1596),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17752_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .I1(_04472_),
    .S(net1543),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17753_ (.I0(_08366_),
    .I1(_08376_),
    .S(net1866),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17754_ (.I0(_04473_),
    .I1(_08373_),
    .S(net1844),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17755_ (.I0(net1512),
    .I1(_04474_),
    .S(net1674),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17756_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .I1(_04475_),
    .S(net1543),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17757_ (.I(net1458),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17758_ (.I0(net1775),
    .I1(_04476_),
    .S(net1596),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17759_ (.I(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17760_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .I1(_04478_),
    .S(net1543),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17761_ (.I(net2174),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17762_ (.I0(net1459),
    .I1(_04479_),
    .S(net1674),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17763_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .I1(_04480_),
    .S(net1543),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17764_ (.A1(_08194_),
    .A2(_04411_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2136 (.I(_01277_),
    .Z(net2135));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17766_ (.A1(net2106),
    .A2(net2084),
    .B(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17767_ (.I(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17768_ (.A1(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .A2(net2106),
    .A3(net2084),
    .B(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17769_ (.A1(_09695_),
    .A2(_09696_),
    .A3(_04483_),
    .A4(_04485_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2137 (.I(net1687),
    .Z(net2136));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17771_ (.A1(net2027),
    .A2(_09700_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17772_ (.A1(_00964_),
    .A2(_04488_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17773_ (.A1(_04486_),
    .A2(_04489_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17774_ (.A1(_04481_),
    .A2(_04490_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17775_ (.A1(_04483_),
    .A2(_04485_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone2138 (.I(net2055),
    .Z(net2137));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17777_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_09696_),
    .A3(_04491_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17778_ (.A1(_00967_),
    .A2(_04488_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17779_ (.A1(_04493_),
    .A2(_04494_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17780_ (.A1(_04481_),
    .A2(_04495_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17781_ (.A1(_00969_),
    .A2(_04488_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17782_ (.A1(_04493_),
    .A2(_04496_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17783_ (.A1(_04481_),
    .A2(_04497_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17784_ (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17785_ (.A1(_04498_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17786_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04499_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17787_ (.A1(_04489_),
    .A2(_04500_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17788_ (.A1(_04481_),
    .A2(_04501_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17789_ (.A1(_00968_),
    .A2(_04488_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17790_ (.A1(_04500_),
    .A2(_04502_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17791_ (.A1(_04481_),
    .A2(_04503_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17792_ (.A1(_04494_),
    .A2(_04500_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17793_ (.A1(_04481_),
    .A2(_04504_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17794_ (.A1(_04496_),
    .A2(_04500_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17795_ (.A1(_04481_),
    .A2(_04505_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17796_ (.A1(_04498_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17797_ (.A1(_09695_),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04506_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17798_ (.A1(_04489_),
    .A2(_04507_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17799_ (.A1(_04481_),
    .A2(_04508_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17800_ (.A1(_04502_),
    .A2(_04507_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17801_ (.A1(_04481_),
    .A2(_04509_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17802_ (.A1(_04494_),
    .A2(_04507_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17803_ (.A1(_04481_),
    .A2(_04510_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2139 (.I(net1407),
    .Z(net2138));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17805_ (.A1(_04496_),
    .A2(_04507_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17806_ (.A1(_04481_),
    .A2(_04512_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17807_ (.I(_04481_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17808_ (.A1(_09695_),
    .A2(_00968_),
    .A3(_09696_),
    .A4(_04491_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17809_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .A2(_04513_),
    .B1(_04514_),
    .B2(_04488_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17810_ (.I(_04515_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17811_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17812_ (.A1(_09695_),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04516_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17813_ (.A1(_04489_),
    .A2(_04517_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17814_ (.A1(_04481_),
    .A2(_04518_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17815_ (.A1(_04502_),
    .A2(_04517_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17816_ (.A1(_04481_),
    .A2(_04519_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17817_ (.A1(_04494_),
    .A2(_04517_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17818_ (.A1(_04481_),
    .A2(_04520_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17819_ (.A1(_04496_),
    .A2(_04517_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17820_ (.A1(_04481_),
    .A2(_04521_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17821_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04506_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17822_ (.A1(_04489_),
    .A2(_04522_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17823_ (.A1(_04481_),
    .A2(_04523_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17824_ (.A1(_04502_),
    .A2(_04522_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17825_ (.A1(_04481_),
    .A2(_04524_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17826_ (.A1(_04494_),
    .A2(_04522_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17827_ (.A1(_04481_),
    .A2(_04525_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17828_ (.A1(_04496_),
    .A2(_04522_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17829_ (.A1(_04481_),
    .A2(_04526_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17830_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04516_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17831_ (.A1(_04489_),
    .A2(_04527_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17832_ (.A1(_04481_),
    .A2(_04528_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1402 (.I(_04770_),
    .Z(net1401));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17834_ (.A1(_04502_),
    .A2(_04527_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17835_ (.A1(_04481_),
    .A2(_04530_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17836_ (.A1(_04486_),
    .A2(_04494_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17837_ (.A1(_04481_),
    .A2(_04531_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17838_ (.A1(_04494_),
    .A2(_04527_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17839_ (.A1(_04481_),
    .A2(_04532_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17840_ (.A1(_04496_),
    .A2(_04527_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17841_ (.A1(_04481_),
    .A2(_04533_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17842_ (.A1(_04486_),
    .A2(_04496_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17843_ (.A1(_04481_),
    .A2(_04534_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17844_ (.A1(_09695_),
    .A2(_04483_),
    .A3(_04485_),
    .A4(_04499_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17845_ (.A1(_04489_),
    .A2(_04535_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17846_ (.A1(_04481_),
    .A2(_04536_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17847_ (.A1(_04502_),
    .A2(_04535_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17848_ (.A1(_04481_),
    .A2(_04537_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17849_ (.A1(_04494_),
    .A2(_04535_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17850_ (.A1(_04481_),
    .A2(_04538_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17851_ (.A1(_04496_),
    .A2(_04535_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17852_ (.A1(_04481_),
    .A2(_04539_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17853_ (.A1(_04489_),
    .A2(_04493_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17854_ (.A1(_04481_),
    .A2(_04540_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1401 (.I(_05237_),
    .Z(net1400));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1400 (.I(_05430_),
    .Z(net1399));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _17857_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .A2(_00968_),
    .A3(_09696_),
    .A4(_04491_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17858_ (.A1(_09700_),
    .A2(_04543_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17859_ (.A1(net2028),
    .A2(_09700_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17860_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .A2(_04545_),
    .B(net2027),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17861_ (.A1(_04544_),
    .A2(_04546_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17862_ (.A1(fetch_enable_q),
    .A2(net66),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17863_ (.A1(_07567_),
    .A2(_07643_),
    .B(_07634_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17864_ (.A1(_07586_),
    .A2(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _17865_ (.A1(_09624_),
    .A2(_10370_),
    .B(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17866_ (.A1(_09699_),
    .A2(_03434_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17867_ (.A1(_04549_),
    .A2(_04550_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 rebuffer2140 (.I(net1933),
    .Z(net2139));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer2141 (.I(net2139),
    .Z(net2140));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 rebuffer2142 (.I(net2139),
    .Z(net2141));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17871_ (.I0(net48),
    .I1(net32),
    .S(net1887),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17872_ (.I0(net62),
    .I1(net39),
    .S(net1887),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17873_ (.I(net1886),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2143 (.I(net1933),
    .Z(net2142));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17875_ (.I0(_04555_),
    .I1(_04556_),
    .S(_04557_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17876_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2144 (.I(_07740_),
    .Z(net2143));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2145 (.I(net1893),
    .Z(net2144));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2146 (.I(net1893),
    .Z(net2145));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2147 (.I(net1888),
    .Z(net2146));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 split2148 (.I(net1888),
    .Z(net2147));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2149 (.I(_08185_),
    .Z(net2148));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17883_ (.I0(net62),
    .I1(\load_store_unit_i.rdata_q[8] ),
    .I2(\load_store_unit_i.rdata_q[16] ),
    .I3(net32),
    .S0(net1887),
    .S1(net1886),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17884_ (.I0(net61),
    .I1(net47),
    .I2(net38),
    .I3(net56),
    .S0(net1886),
    .S1(net1887),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17885_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_04568_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _17886_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_04559_),
    .B1(_04560_),
    .B2(_04567_),
    .C(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17887_ (.A1(_04549_),
    .A2(_04550_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2150 (.I(_07570_),
    .Z(net2149));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2151 (.I(_01225_),
    .Z(net2150));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17890_ (.I(_01137_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17891_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_07599_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17892_ (.I(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17893_ (.A1(_04574_),
    .A2(net1611),
    .A3(_01159_),
    .B(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17894_ (.A1(_01166_),
    .A2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2152 (.I(net1931),
    .Z(net2151));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17896_ (.A1(_07773_),
    .A2(_09568_),
    .B(_04575_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17897_ (.A1(net1702),
    .A2(_04580_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 split2153 (.I(net1931),
    .Z(net2152));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17899_ (.A1(_03415_),
    .A2(_03396_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17900_ (.I0(net1691),
    .I1(_01312_),
    .S(net1616),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2154 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net2153));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17902_ (.I0(net1692),
    .I1(_01319_),
    .S(net1616),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17903_ (.I0(_04584_),
    .I1(_04586_),
    .S(net1612),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17904_ (.I0(net2072),
    .I1(net1678),
    .S(net1616),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17905_ (.I0(net2116),
    .I1(net1677),
    .S(net1616),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17906_ (.I0(_04588_),
    .I1(_04589_),
    .S(net1612),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 rebuffer2155 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net2154));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17908_ (.I0(_01145_),
    .I1(_01151_),
    .I2(_01347_),
    .I3(net1675),
    .S0(net1703),
    .S1(net1616),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2160 (.I(net1695),
    .Z(net2159));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17910_ (.I0(net2103),
    .I1(_01165_),
    .I2(net1676),
    .I3(_01326_),
    .S0(net1703),
    .S1(net1616),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17911_ (.I(_01138_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17912_ (.I0(_04595_),
    .I1(net2289),
    .S(_04575_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2159 (.I(net1787),
    .Z(net2158));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2158 (.I(net1774),
    .Z(net2157));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17915_ (.A1(_04574_),
    .A2(_04576_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17916_ (.A1(_07773_),
    .A2(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2157 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net2156));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17918_ (.I0(_04587_),
    .I1(_04590_),
    .I2(_04592_),
    .I3(_04594_),
    .S0(_04596_),
    .S1(_04600_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17919_ (.A1(_04581_),
    .A2(_04602_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17920_ (.A1(_08082_),
    .A2(_08099_),
    .A3(net1616),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17921_ (.A1(_09470_),
    .A2(net1616),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17922_ (.A1(_04604_),
    .A2(_04605_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17923_ (.I0(_01138_),
    .I1(net1586),
    .S(_04575_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2156 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net2155));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17925_ (.A1(_08121_),
    .A2(_08126_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17926_ (.A1(_03395_),
    .A2(_04609_),
    .A3(_03396_),
    .Z(_04610_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17927_ (.A1(net1612),
    .A2(_04600_),
    .A3(_04607_),
    .B(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17928_ (.A1(_01159_),
    .A2(_04580_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2162 (.I(net2160),
    .Z(net2161));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _17930_ (.A1(_04606_),
    .A2(_04611_),
    .B(_04612_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17931_ (.A1(_09470_),
    .A2(_04610_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 rebuffer2161 (.I(net1728),
    .Z(net2160));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17933_ (.A1(_04578_),
    .A2(_04615_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _17934_ (.A1(_04578_),
    .A2(_04603_),
    .A3(_04614_),
    .B(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17935_ (.I0(_01165_),
    .I1(net1692),
    .I2(_01326_),
    .I3(_01319_),
    .S0(net1703),
    .S1(net1616),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17936_ (.I0(_04584_),
    .I1(_04589_),
    .S(net1703),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17937_ (.I0(_01145_),
    .I1(_01139_),
    .I2(_01347_),
    .I3(_00938_),
    .S0(net1612),
    .S1(net1616),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17938_ (.I0(_01151_),
    .I1(net2103),
    .I2(net1675),
    .I3(net1676),
    .S0(net1703),
    .S1(net1616),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17939_ (.I0(_04619_),
    .I1(_04620_),
    .I2(_04621_),
    .I3(_04622_),
    .S0(net1551),
    .S1(_04600_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17940_ (.I0(net2070),
    .I1(net1682),
    .S(net1616),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17941_ (.I0(net1704),
    .I1(net1681),
    .S(net1616),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17942_ (.I0(_04624_),
    .I1(_04625_),
    .S(net1612),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17943_ (.I0(net1685),
    .I1(_01256_),
    .S(net1616),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17944_ (.I0(net1684),
    .I1(net1683),
    .S(net1616),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17945_ (.I0(_04627_),
    .I1(_04628_),
    .S(net1703),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17946_ (.I0(net2097),
    .I1(net1679),
    .S(net1616),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17947_ (.I0(_04588_),
    .I1(_04630_),
    .S(net1703),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17948_ (.I0(net2159),
    .I1(net2135),
    .S(net1616),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17949_ (.I0(net2102),
    .I1(net1680),
    .S(net1616),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17950_ (.I0(_04632_),
    .I1(_04633_),
    .S(net1612),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17951_ (.I0(_04626_),
    .I1(_04629_),
    .I2(_04631_),
    .I3(_04634_),
    .S0(net1551),
    .S1(_04600_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17952_ (.A1(_03415_),
    .A2(_03396_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2163 (.I(net1996),
    .Z(net2162));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17954_ (.I0(net2102),
    .I1(net1680),
    .S(_04636_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17955_ (.I0(net2159),
    .I1(net2135),
    .S(_04636_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17956_ (.I0(_04638_),
    .I1(_04639_),
    .S(net1612),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17957_ (.I0(net2072),
    .I1(net1678),
    .S(_04636_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17958_ (.I0(net2097),
    .I1(net1679),
    .S(_04636_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17959_ (.I0(_04641_),
    .I1(_04642_),
    .S(net1612),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17960_ (.I0(net1685),
    .I1(_01256_),
    .S(_04636_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17961_ (.I0(net1684),
    .I1(net1683),
    .S(_04636_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17962_ (.I0(_04644_),
    .I1(_04645_),
    .S(net1612),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17963_ (.I0(net1704),
    .I1(net1681),
    .S(_04636_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17964_ (.I0(net2070),
    .I1(net1682),
    .S(_04636_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17965_ (.I0(_04647_),
    .I1(_04648_),
    .S(net1612),
    .Z(_04649_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1399 (.I(_04491_),
    .Z(net1398));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17967_ (.I0(_04640_),
    .I1(_04643_),
    .I2(_04646_),
    .I3(_04649_),
    .S0(net1551),
    .S1(_04600_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2164 (.I(net1996),
    .Z(net2163));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _17969_ (.A1(net1701),
    .A2(_04577_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2165 (.I(net1996),
    .Z(net2164));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2166 (.I(net1996),
    .Z(net2165));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _17972_ (.I0(_04615_),
    .I1(_04623_),
    .I2(_04635_),
    .I3(_04651_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2167 (.I(net1996),
    .Z(net2166));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17974_ (.I0(_04618_),
    .I1(_04656_),
    .S(_04583_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17975_ (.A1(net1782),
    .A2(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _17976_ (.A1(_08128_),
    .A2(_03412_),
    .A3(_08216_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2168 (.I(_08448_),
    .Z(net2167));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17978_ (.A1(_08128_),
    .A2(_03396_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17979_ (.A1(_03394_),
    .A2(_04662_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17980_ (.A1(_08127_),
    .A2(_03412_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _17981_ (.A1(_04663_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone2169 (.I(net2090),
    .Z(net2168));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17983_ (.I(_03396_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _17984_ (.I0(_03395_),
    .I1(_08129_),
    .S(_03394_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17985_ (.A1(_04667_),
    .A2(_08217_),
    .A3(_04668_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2170 (.I(net175),
    .Z(net2169));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1398 (.I(_04924_),
    .Z(net1397));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _17988_ (.A1(_08217_),
    .A2(_03394_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2171 (.I(net1889),
    .Z(net2170));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17990_ (.A1(_01195_),
    .A2(net1614),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _17991_ (.A1(_08217_),
    .A2(_03394_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _17992_ (.A1(net1587),
    .A2(_04675_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2172 (.I(_08928_),
    .Z(net2171));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _17994_ (.A1(_01196_),
    .A2(net1578),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _17995_ (.A1(_01199_),
    .A2(net1587),
    .B(_04674_),
    .C(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _17996_ (.A1(net1458),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17997_ (.I(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _17998_ (.A1(_00086_),
    .A2(_01000_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _17999_ (.A1(net2030),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A3(net1751),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18000_ (.A1(net1718),
    .A2(_04683_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1397 (.I(_05290_),
    .Z(net1396));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18002_ (.I0(_04681_),
    .I1(_04682_),
    .S(_04684_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18003_ (.I0(_04680_),
    .I1(_04686_),
    .S(net1815),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18004_ (.A1(_11007_),
    .A2(net1507),
    .A3(_04659_),
    .A4(_04687_),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18005_ (.A1(net1508),
    .A2(_04570_),
    .B(_04688_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2173 (.I(_00889_),
    .Z(net2172));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18007_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18008_ (.A1(net30),
    .A2(\load_store_unit_i.lsu_err_q ),
    .A3(\load_store_unit_i.data_we_q ),
    .A4(_09654_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18009_ (.A1(_09538_),
    .A2(_03433_),
    .B1(_04548_),
    .B2(_09585_),
    .C(_09686_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18010_ (.A1(_09585_),
    .A2(_09637_),
    .B(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18011_ (.A1(_04692_),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18012_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_04695_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18013_ (.A1(_04691_),
    .A2(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2174 (.I(_00857_),
    .Z(net2173));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18015_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .I1(net1392),
    .S(_04697_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18016_ (.I0(net49),
    .I1(net43),
    .S(net1887),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18017_ (.I0(net63),
    .I1(net40),
    .S(net1887),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18018_ (.I0(_04699_),
    .I1(_04700_),
    .S(_04557_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2175 (.I(net1736),
    .Z(net2174));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18020_ (.I0(net63),
    .I1(\load_store_unit_i.rdata_q[9] ),
    .I2(\load_store_unit_i.rdata_q[17] ),
    .I3(net43),
    .S0(net1887),
    .S1(net1886),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18021_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_04701_),
    .B1(_04703_),
    .B2(_04560_),
    .C(_04569_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone2176 (.I(net2180),
    .Z(net2175));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18023_ (.A1(net1612),
    .A2(_04610_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18024_ (.A1(_04604_),
    .A2(_04605_),
    .A3(_04706_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18025_ (.I0(_04587_),
    .I1(_04592_),
    .I2(_04594_),
    .I3(_04707_),
    .S0(_04600_),
    .S1(_04607_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18026_ (.I0(_04625_),
    .I1(_04632_),
    .S(net1612),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18027_ (.I0(_04630_),
    .I1(_04633_),
    .S(net1703),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18028_ (.I0(_04624_),
    .I1(_04627_),
    .S(net1703),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18029_ (.A1(net1611),
    .A2(_04599_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2177 (.I(_01236_),
    .Z(net2176));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18031_ (.I0(_04590_),
    .I1(_04709_),
    .I2(_04710_),
    .I3(_04711_),
    .S0(_04712_),
    .S1(net1551),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18032_ (.I0(_04639_),
    .I1(_04647_),
    .S(net1612),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18033_ (.I0(_04638_),
    .I1(_04642_),
    .S(net1703),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18034_ (.A1(net1703),
    .A2(_04636_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18035_ (.I0(net1684),
    .I1(net1683),
    .S(_04717_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18036_ (.I0(_04644_),
    .I1(_04648_),
    .S(net1703),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18037_ (.I0(_04715_),
    .I1(_04716_),
    .I2(_04718_),
    .I3(_04719_),
    .S0(net1551),
    .S1(_04600_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2178 (.I(_07622_),
    .Z(net2177));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18039_ (.I0(_04615_),
    .I1(_04708_),
    .I2(_04714_),
    .I3(_04720_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18040_ (.A1(net1782),
    .A2(_04583_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18041_ (.A1(_04722_),
    .A2(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2179 (.I(_08383_),
    .Z(net2178));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2180 (.I(net1913),
    .Z(net2179));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2181 (.I(_08218_),
    .Z(net2180));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18045_ (.A1(_09470_),
    .A2(_04610_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18046_ (.A1(_04712_),
    .A2(net1551),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18047_ (.A1(_04581_),
    .A2(_04729_),
    .B(_04578_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18048_ (.I0(_04619_),
    .I1(_04622_),
    .I2(_04631_),
    .I3(_04620_),
    .S0(_04607_),
    .S1(_04712_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18049_ (.A1(_04653_),
    .A2(_04612_),
    .A3(_04731_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18050_ (.I(_04621_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18051_ (.A1(_04578_),
    .A2(_04612_),
    .A3(_04729_),
    .A4(_04733_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18052_ (.A1(_04728_),
    .A2(_04730_),
    .B(_04732_),
    .C(_04734_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18053_ (.A1(_03415_),
    .A2(_08217_),
    .A3(_08170_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18054_ (.A1(_04663_),
    .A2(_04664_),
    .Z(_04737_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18055_ (.A1(_01206_),
    .A2(net1587),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18056_ (.A1(_01202_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01203_),
    .C(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18057_ (.A1(_08455_),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18058_ (.I(_01000_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18059_ (.A1(net1452),
    .A2(_00995_),
    .B(_00994_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18060_ (.I(_00999_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18061_ (.A1(_04741_),
    .A2(_04742_),
    .B(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18062_ (.A1(_01005_),
    .A2(_04744_),
    .Z(_04745_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18063_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(_04745_),
    .S(_04684_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18064_ (.I0(_04740_),
    .I1(_04746_),
    .S(net1815),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18065_ (.A1(net1615),
    .A2(_04735_),
    .B(_04747_),
    .C(_11022_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18066_ (.A1(net1507),
    .A2(_04724_),
    .A3(_04748_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18067_ (.A1(net1508),
    .A2(_04704_),
    .B(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2182 (.I(_07654_),
    .Z(net2181));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18069_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .I1(net1388),
    .S(net1497),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18070_ (.I0(net33),
    .I1(\load_store_unit_i.rdata_q[10] ),
    .I2(\load_store_unit_i.rdata_q[18] ),
    .I3(net54),
    .S0(net1887),
    .S1(net1886),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18071_ (.I0(net50),
    .I1(net54),
    .S(net1887),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18072_ (.I0(net33),
    .I1(net41),
    .S(net1887),
    .Z(_04754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18073_ (.I0(_04753_),
    .I1(_04754_),
    .S(_04557_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18074_ (.A1(net1833),
    .A2(_04752_),
    .B1(_04755_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_04569_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18075_ (.I0(_04615_),
    .I1(_04621_),
    .I2(_04622_),
    .I3(_04619_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18076_ (.I0(_04620_),
    .I1(_04631_),
    .I2(_04634_),
    .I3(_04626_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18077_ (.I0(_04629_),
    .I1(_04646_),
    .I2(_04649_),
    .I3(_04640_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18078_ (.I0(_04615_),
    .I1(_04757_),
    .I2(_04758_),
    .I3(_04759_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18079_ (.I0(_04592_),
    .I1(_04707_),
    .S(_04607_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18080_ (.I0(_04615_),
    .I1(_04761_),
    .S(_04712_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18081_ (.I0(_04587_),
    .I1(_04594_),
    .I2(_04710_),
    .I3(_04590_),
    .S0(_04607_),
    .S1(_04712_),
    .Z(_04763_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18082_ (.A1(_04581_),
    .A2(_04763_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18083_ (.A1(_04612_),
    .A2(_04762_),
    .B(_04764_),
    .C(_04653_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18084_ (.A1(_03396_),
    .A2(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18085_ (.A1(_03396_),
    .A2(_04760_),
    .B(_04766_),
    .C(net1782),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2183 (.I(net2139),
    .Z(net2182));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18087_ (.A1(_00086_),
    .A2(_04741_),
    .B(_04743_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18088_ (.A1(_01005_),
    .A2(_04769_),
    .B(_01004_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18089_ (.A1(_01009_),
    .A2(net1401),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2184 (.I(_07600_),
    .Z(net2183));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18091_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(_04771_),
    .S(_04684_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2185 (.I(net2090),
    .Z(net2184));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2186 (.I(net1796),
    .Z(net2185));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2187 (.I(_00905_),
    .Z(net2186));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18095_ (.A1(_01213_),
    .A2(net1587),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18096_ (.A1(_01209_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01210_),
    .C(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18097_ (.A1(_08509_),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_04778_),
    .C(net1783),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18098_ (.A1(net1783),
    .A2(_04773_),
    .B(_04779_),
    .C(_09585_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18099_ (.A1(_11031_),
    .A2(net1507),
    .A3(_04767_),
    .A4(_04780_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18100_ (.A1(net1508),
    .A2(_04756_),
    .B(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2188 (.I(net1772),
    .Z(net2187));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18102_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .I1(net1381),
    .S(net1498),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18103_ (.I0(net34),
    .I1(\load_store_unit_i.rdata_q[11] ),
    .I2(\load_store_unit_i.rdata_q[19] ),
    .I3(net57),
    .S0(net1887),
    .S1(net1886),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18104_ (.I0(net51),
    .I1(net57),
    .S(net1887),
    .Z(_04785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18105_ (.I0(net34),
    .I1(net42),
    .S(net1887),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18106_ (.I0(_04785_),
    .I1(_04786_),
    .S(_04557_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18107_ (.A1(net1833),
    .A2(_04784_),
    .B1(_04787_),
    .B2(\load_store_unit_i.data_type_q[2] ),
    .C(_04569_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18108_ (.I(_01008_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18109_ (.I(_01009_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18110_ (.A1(_01005_),
    .A2(_04744_),
    .B(_01004_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18111_ (.A1(_04790_),
    .A2(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18112_ (.A1(_04789_),
    .A2(_04792_),
    .Z(_04793_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18113_ (.A1(net1444),
    .A2(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18114_ (.I0(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .I1(_04794_),
    .S(_04684_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18115_ (.A1(_08187_),
    .A2(_04795_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18116_ (.A1(net1457),
    .A2(_04660_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18117_ (.A1(_01216_),
    .A2(net1614),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18118_ (.A1(_01217_),
    .A2(net1578),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18119_ (.A1(_01220_),
    .A2(net1587),
    .B(_04798_),
    .C(_04799_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18120_ (.A1(_04665_),
    .A2(_04800_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18121_ (.A1(_04596_),
    .A2(_04592_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18122_ (.A1(_04607_),
    .A2(_04594_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18123_ (.A1(net1782),
    .A2(_04667_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18124_ (.I(_04804_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18125_ (.A1(_03406_),
    .A2(_04805_),
    .B1(_04596_),
    .B2(net1703),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18126_ (.A1(_04606_),
    .A2(_04600_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _18127_ (.A1(_04600_),
    .A2(_04802_),
    .A3(_04803_),
    .B1(_04806_),
    .B2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18128_ (.I0(_04587_),
    .I1(_04590_),
    .S(net1551),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18129_ (.I0(_04709_),
    .I1(_04710_),
    .S(_04607_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18130_ (.I0(_04809_),
    .I1(_04810_),
    .S(_04712_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18131_ (.I0(_04715_),
    .I1(_04719_),
    .S(_04607_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18132_ (.I0(_04711_),
    .I1(_04718_),
    .S(net1551),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18133_ (.I0(_04812_),
    .I1(_04813_),
    .S(_04600_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18134_ (.I0(_04615_),
    .I1(_04808_),
    .I2(_04811_),
    .I3(_04814_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18135_ (.A1(net1783),
    .A2(_04583_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18136_ (.A1(_04797_),
    .A2(_04801_),
    .A3(_04815_),
    .A4(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18137_ (.A1(_04653_),
    .A2(_04581_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18138_ (.I0(_04621_),
    .I1(_04622_),
    .S(net1551),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18139_ (.I0(_04615_),
    .I1(_04819_),
    .S(_04712_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone2189 (.I(net1944),
    .Z(net2188));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18141_ (.I0(_04619_),
    .I1(_04620_),
    .I2(_04631_),
    .I3(_04634_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18142_ (.A1(_04653_),
    .A2(_04612_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18143_ (.A1(_04578_),
    .A2(_04615_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18144_ (.A1(_04818_),
    .A2(_04820_),
    .B1(_04822_),
    .B2(_04823_),
    .C(_04824_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18145_ (.A1(_04665_),
    .A2(_04800_),
    .B(_04797_),
    .C(net1782),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18146_ (.A1(net1615),
    .A2(_04825_),
    .B1(_04826_),
    .B2(net1783),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18147_ (.A1(_04796_),
    .A2(_04817_),
    .A3(_04827_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18148_ (.A1(_10346_),
    .A2(net1508),
    .A3(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18149_ (.A1(net1508),
    .A2(_04788_),
    .B(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2190 (.I(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net2189));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18151_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .I1(net1376),
    .S(_04697_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18152_ (.I0(net52),
    .I1(net58),
    .S(net1887),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18153_ (.I0(net35),
    .I1(net44),
    .S(net1887),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18154_ (.I0(_04832_),
    .I1(_04833_),
    .S(_04557_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18155_ (.I0(net35),
    .I1(\load_store_unit_i.rdata_q[12] ),
    .I2(\load_store_unit_i.rdata_q[20] ),
    .I3(net58),
    .S0(net1887),
    .S1(net1886),
    .Z(_04835_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2191 (.I(net1771),
    .Z(net2190));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18157_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_04834_),
    .B1(_04835_),
    .B2(net1833),
    .C(_04569_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18158_ (.I(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18159_ (.I0(_04808_),
    .I1(_04811_),
    .S(_04612_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2192 (.I(_08669_),
    .Z(net2191));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18161_ (.A1(_04653_),
    .A2(_04839_),
    .B(_04583_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2193 (.I(net1773),
    .Z(net2192));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18163_ (.A1(_01227_),
    .A2(net1614),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18164_ (.A1(_01224_),
    .A2(net1578),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18165_ (.A1(_01223_),
    .A2(net1587),
    .B(_04843_),
    .C(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18166_ (.A1(net2298),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18167_ (.I0(_04626_),
    .I1(_04629_),
    .I2(_04646_),
    .I3(_04649_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18168_ (.I0(_04615_),
    .I1(_04820_),
    .I2(_04822_),
    .I3(_04847_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18169_ (.A1(net1615),
    .A2(_04848_),
    .B(net1782),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18170_ (.A1(net1783),
    .A2(_04846_),
    .A3(_04849_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18171_ (.A1(_04790_),
    .A2(net1401),
    .B(_04789_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18172_ (.A1(net1444),
    .A2(_04851_),
    .B(net1445),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18173_ (.A1(_01017_),
    .A2(_04852_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18174_ (.I0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .I1(net1391),
    .S(_04684_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18175_ (.A1(_08187_),
    .A2(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18176_ (.A1(_04841_),
    .A2(_04850_),
    .A3(_04855_),
    .B(_11050_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clone2194 (.I(net2005),
    .Z(net2193));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18178_ (.I0(_04838_),
    .I1(_04856_),
    .S(net1507),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2195 (.I(_08817_),
    .Z(net2194));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18180_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .I1(net1375),
    .S(net1497),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18181_ (.I(net1887),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2273 (.I(_08252_),
    .Z(net2272));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18183_ (.A1(_04557_),
    .A2(net1887),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2277 (.I(_06353_),
    .Z(net2276));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18185_ (.A1(net1886),
    .A2(_04860_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18186_ (.A1(\load_store_unit_i.rdata_q[13] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18187_ (.A1(_04860_),
    .A2(net53),
    .B1(net45),
    .B2(_04862_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18188_ (.I0(_04865_),
    .I1(_04866_),
    .S(\load_store_unit_i.data_type_q[2] ),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18189_ (.A1(net1887),
    .A2(net59),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18190_ (.A1(_04867_),
    .A2(_04868_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18191_ (.A1(_04557_),
    .A2(_04860_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18192_ (.A1(net36),
    .A2(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18193_ (.A1(_04860_),
    .A2(_04867_),
    .B1(_04869_),
    .B2(_04557_),
    .C(_04871_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18194_ (.I(\load_store_unit_i.data_type_q[2] ),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18195_ (.A1(_04873_),
    .A2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18196_ (.A1(_04872_),
    .A2(_04874_),
    .B(_04569_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18197_ (.A1(_01230_),
    .A2(net1614),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18198_ (.A1(_01231_),
    .A2(net1578),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18199_ (.A1(_01234_),
    .A2(net1587),
    .B(_04876_),
    .C(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18200_ (.A1(net1450),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18201_ (.I(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18202_ (.A1(_01008_),
    .A2(net1445),
    .A3(_01016_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18203_ (.A1(_01011_),
    .A2(_01010_),
    .B(_01017_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18204_ (.I(_01016_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18205_ (.A1(_04792_),
    .A2(net1427),
    .B1(_04882_),
    .B2(net1426),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18206_ (.A1(net1442),
    .A2(_04884_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18207_ (.I0(_04880_),
    .I1(_04885_),
    .S(_04684_),
    .Z(_04886_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2279 (.I(net1433),
    .Z(net2278));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18209_ (.I0(_04879_),
    .I1(_04886_),
    .S(net1815),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18210_ (.I0(_04709_),
    .I1(_04711_),
    .I2(_04718_),
    .I3(_04719_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18211_ (.I0(_04762_),
    .I1(_04889_),
    .S(_04653_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18212_ (.I0(_04615_),
    .I1(_04763_),
    .S(_04653_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18213_ (.I0(_04890_),
    .I1(_04891_),
    .S(_04581_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18214_ (.I0(_04757_),
    .I1(_04758_),
    .S(_04612_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18215_ (.A1(_04653_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18216_ (.A1(_03396_),
    .A2(_04894_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18217_ (.A1(_03396_),
    .A2(_04892_),
    .B(_04895_),
    .C(net1782),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18218_ (.A1(_10446_),
    .A2(net1507),
    .A3(_04888_),
    .A4(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18219_ (.A1(net1508),
    .A2(_04875_),
    .B(_04897_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2289 (.I(net1447),
    .Z(net2288));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18221_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .I1(net1377),
    .S(net1498),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18222_ (.I0(net55),
    .I1(net60),
    .S(net1887),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18223_ (.I0(net37),
    .I1(net46),
    .S(net1887),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18224_ (.I0(_04900_),
    .I1(_04901_),
    .S(_04557_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18225_ (.I0(net37),
    .I1(\load_store_unit_i.rdata_q[14] ),
    .I2(\load_store_unit_i.rdata_q[22] ),
    .I3(net60),
    .S0(net1887),
    .S1(net1886),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18226_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_04902_),
    .B1(_04903_),
    .B2(_04560_),
    .C(_04569_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2288 (.I(_08819_),
    .Z(net2287));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2290 (.I(_01135_),
    .Z(net2289));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1396 (.I(_03437_),
    .Z(net1395));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18230_ (.A1(_01241_),
    .A2(net1587),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18231_ (.A1(_01237_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01238_),
    .C(_04908_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18232_ (.A1(net2292),
    .A2(_04660_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18233_ (.A1(_04737_),
    .A2(_04909_),
    .B(_04910_),
    .C(net1783),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18234_ (.I(_04723_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18235_ (.A1(_04581_),
    .A2(_04729_),
    .A3(_04733_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18236_ (.A1(_04581_),
    .A2(_04729_),
    .B(_04615_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18237_ (.A1(_04578_),
    .A2(_04913_),
    .A3(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18238_ (.I0(_04626_),
    .I1(_04634_),
    .I2(_04646_),
    .I3(_04629_),
    .S0(_04607_),
    .S1(_04712_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18239_ (.I0(_04731_),
    .I1(_04916_),
    .S(_04612_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18240_ (.A1(_04578_),
    .A2(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18241_ (.I0(_04708_),
    .I1(_04714_),
    .S(_04612_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18242_ (.A1(_04653_),
    .A2(_04919_),
    .B(_04824_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _18243_ (.A1(_04912_),
    .A2(_04915_),
    .A3(_04918_),
    .B1(_04920_),
    .B2(_04583_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18244_ (.A1(_04883_),
    .A2(_04882_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18245_ (.A1(_01023_),
    .A2(_04922_),
    .Z(_04923_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18246_ (.A1(_04770_),
    .A2(_04790_),
    .B(net1427),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18247_ (.A1(_04923_),
    .A2(net1397),
    .B(net1443),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18248_ (.A1(net1441),
    .A2(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18249_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(_04926_),
    .S(_04684_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18250_ (.A1(_08187_),
    .A2(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18251_ (.A1(_04911_),
    .A2(_04921_),
    .B(_04928_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18252_ (.A1(_11062_),
    .A2(net1507),
    .A3(_04929_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18253_ (.A1(net1508),
    .A2(_04904_),
    .B(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2291 (.I(_00833_),
    .Z(net2290));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18255_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .I1(net1371),
    .S(net1497),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1394 (.I(_03449_),
    .Z(net1393));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1393 (.I(_04689_),
    .Z(net1392));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18258_ (.I0(net38),
    .I1(\load_store_unit_i.rdata_q[15] ),
    .I2(\load_store_unit_i.rdata_q[23] ),
    .I3(net61),
    .S0(net1887),
    .S1(net1886),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18259_ (.I0(net56),
    .I1(net61),
    .S(net1887),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18260_ (.I0(net38),
    .I1(net47),
    .S(net1887),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18261_ (.I0(_04936_),
    .I1(_04937_),
    .S(_04557_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18262_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_04938_),
    .Z(_04939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18263_ (.A1(_04560_),
    .A2(_04935_),
    .B(_04939_),
    .C(_04569_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18264_ (.I0(_04623_),
    .I1(_04635_),
    .S(_04612_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18265_ (.I0(_04615_),
    .I1(_04941_),
    .S(_04653_),
    .Z(_04942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18266_ (.A1(_04606_),
    .A2(_04611_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18267_ (.I0(_04810_),
    .I1(_04813_),
    .S(_04712_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18268_ (.I0(_04615_),
    .I1(_04602_),
    .I2(_04943_),
    .I3(_04944_),
    .S0(_04653_),
    .S1(_04612_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18269_ (.I0(_04942_),
    .I1(_04945_),
    .S(_04583_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18270_ (.A1(net1782),
    .A2(_04946_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18271_ (.A1(_01244_),
    .A2(net1614),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18272_ (.A1(_01245_),
    .A2(net1578),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18273_ (.A1(_01248_),
    .A2(net1587),
    .B(_04948_),
    .C(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18274_ (.A1(net1448),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18275_ (.I(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18276_ (.A1(net1443),
    .A2(_01026_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18277_ (.A1(_04791_),
    .A2(_04790_),
    .B(net1427),
    .C(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18278_ (.A1(net1442),
    .A2(net1405),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18279_ (.A1(net1441),
    .A2(_01026_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18280_ (.A1(_04955_),
    .A2(_04953_),
    .B(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18281_ (.A1(net1439),
    .A2(_04954_),
    .A3(_04957_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18282_ (.A1(_04954_),
    .A2(_04957_),
    .B(net1439),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18283_ (.A1(_04958_),
    .A2(_04959_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18284_ (.I0(_04952_),
    .I1(_04960_),
    .S(_04684_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18285_ (.I0(_04951_),
    .I1(_04961_),
    .S(net1815),
    .Z(_04962_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18286_ (.A1(_10491_),
    .A2(net1507),
    .A3(_04947_),
    .A4(_04962_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18287_ (.A1(net1508),
    .A2(_04940_),
    .B(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1392 (.I(_04853_),
    .Z(net1391));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18289_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .I1(net1374),
    .S(net1497),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18290_ (.I0(_04942_),
    .I1(_04945_),
    .S(net1615),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1395 (.I(net1393),
    .Z(net1394));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18292_ (.A1(_01255_),
    .A2(net1587),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18293_ (.A1(_01251_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01252_),
    .C(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _18294_ (.A1(net1455),
    .A2(_08839_),
    .A3(_04736_),
    .B1(_04737_),
    .B2(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18295_ (.A1(net1441),
    .A2(net1439),
    .A3(_04923_),
    .Z(_04971_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18296_ (.A1(_01027_),
    .A2(_01033_),
    .A3(_01022_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18297_ (.A1(net1439),
    .A2(_01026_),
    .B(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18298_ (.I(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18299_ (.A1(net1397),
    .A2(_04971_),
    .B(_04974_),
    .C(net1440),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18300_ (.A1(net1437),
    .A2(_04975_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1391 (.I(_05101_),
    .Z(net1390));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18302_ (.I0(_00972_),
    .I1(_04976_),
    .S(_04683_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18303_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(_04978_),
    .S(net1718),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18304_ (.I0(_04970_),
    .I1(_04979_),
    .S(net1815),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18305_ (.A1(net1782),
    .A2(_04966_),
    .B(_04980_),
    .C(_10523_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18306_ (.I0(net39),
    .I1(net32),
    .I2(\load_store_unit_i.rdata_q[16] ),
    .I3(net62),
    .S0(net1886),
    .S1(net1887),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18307_ (.A1(\load_store_unit_i.data_sign_ext_q ),
    .A2(_04939_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18308_ (.A1(_04569_),
    .A2(_04983_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2292 (.I(_08399_),
    .Z(net2291));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18310_ (.A1(_03455_),
    .A2(_04693_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2293 (.I(net1456),
    .Z(net2292));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18312_ (.A1(net1833),
    .A2(_04982_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18313_ (.A1(net1507),
    .A2(net1373),
    .B(_04988_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2466 (.I(net2469),
    .Z(net2465));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18315_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .I1(net1370),
    .S(net1498),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18316_ (.I0(net40),
    .I1(net43),
    .I2(\load_store_unit_i.rdata_q[17] ),
    .I3(net63),
    .S0(net1886),
    .S1(net1887),
    .Z(_04991_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18317_ (.A1(_04560_),
    .A2(_04991_),
    .B(_04984_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18318_ (.A1(_04915_),
    .A2(_04918_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18319_ (.A1(_01258_),
    .A2(net1614),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18320_ (.A1(_01259_),
    .A2(net1578),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18321_ (.A1(_01262_),
    .A2(net1587),
    .B(_04994_),
    .C(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18322_ (.A1(_09585_),
    .A2(net1783),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18323_ (.A1(net2288),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_04996_),
    .C(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18324_ (.A1(_04920_),
    .A2(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18325_ (.I0(_04993_),
    .I1(_04999_),
    .S(_04583_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18326_ (.A1(net1440),
    .A2(_04958_),
    .Z(_05001_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18327_ (.A1(net1437),
    .A2(_05001_),
    .B(net1438),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18328_ (.A1(net1424),
    .A2(_05002_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18329_ (.I0(_00974_),
    .I1(_05003_),
    .S(_04683_),
    .Z(_05004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18330_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(_05004_),
    .S(net1718),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18331_ (.A1(net1783),
    .A2(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18332_ (.A1(_08043_),
    .A2(_11087_),
    .B1(_04998_),
    .B2(_04609_),
    .C(_05006_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18333_ (.A1(_05000_),
    .A2(_05007_),
    .B(net1508),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18334_ (.A1(net1508),
    .A2(_04992_),
    .B(net1367),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2301 (.I(_08388_),
    .Z(net2300));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18336_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .I1(net1362),
    .S(net1497),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18337_ (.A1(_01171_),
    .A2(net1587),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18338_ (.A1(_01167_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01168_),
    .C(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18339_ (.A1(net1454),
    .A2(_04660_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18340_ (.A1(_04737_),
    .A2(_05012_),
    .B(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18341_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(_00981_),
    .S(_04684_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18342_ (.I0(_05014_),
    .I1(_05015_),
    .S(net1815),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18343_ (.A1(_04578_),
    .A2(_04581_),
    .B(_04728_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18344_ (.A1(_04578_),
    .A2(_04581_),
    .A3(_04808_),
    .B(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18345_ (.I0(net1691),
    .I1(_01312_),
    .S(_04636_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18346_ (.I0(net2116),
    .I1(net1677),
    .S(_04636_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18347_ (.I0(_05019_),
    .I1(_05020_),
    .S(net1612),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18348_ (.A1(_01319_),
    .A2(net1616),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18349_ (.A1(_01176_),
    .A2(net1616),
    .Z(_05023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18350_ (.A1(_08297_),
    .A2(_08317_),
    .B(_04636_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18351_ (.A1(_01326_),
    .A2(net1616),
    .B(net1703),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _18352_ (.A1(net1703),
    .A2(_05022_),
    .A3(_05023_),
    .B1(_05024_),
    .B2(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18353_ (.I0(_04640_),
    .I1(_04643_),
    .I2(_05021_),
    .I3(_05026_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18354_ (.I0(_04820_),
    .I1(_04822_),
    .I2(_04847_),
    .I3(_05027_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18355_ (.A1(net1615),
    .A2(_05028_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18356_ (.A1(net1615),
    .A2(_05018_),
    .B(_05029_),
    .C(_04609_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18357_ (.A1(_10909_),
    .A2(net1508),
    .A3(_05016_),
    .A4(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18358_ (.A1(net1886),
    .A2(_04860_),
    .A3(net44),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18359_ (.A1(_04557_),
    .A2(net1887),
    .A3(net35),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18360_ (.A1(_05032_),
    .A2(_05033_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18361_ (.A1(\load_store_unit_i.rdata_q[4] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[12] ),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18362_ (.I0(_05034_),
    .I1(_05035_),
    .S(net1833),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18363_ (.A1(net1886),
    .A2(net1887),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18364_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net52),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18365_ (.A1(_05037_),
    .A2(_05038_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18366_ (.A1(net58),
    .A2(_04870_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18367_ (.A1(_04694_),
    .A2(_05036_),
    .A3(_05039_),
    .A4(_05040_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18368_ (.A1(_05031_),
    .A2(_05041_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2294 (.I(net1428),
    .Z(net2293));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18370_ (.A1(_04692_),
    .A2(_04694_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18371_ (.A1(_07968_),
    .A2(_09519_),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_05044_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18372_ (.A1(_09518_),
    .A2(_05045_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2300 (.I(_07808_),
    .Z(net2299));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18374_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net1496),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18375_ (.A1(_04617_),
    .A2(_04894_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18376_ (.I0(_04892_),
    .I1(_05048_),
    .S(_04667_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18377_ (.A1(_01269_),
    .A2(net1587),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18378_ (.A1(_01265_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01266_),
    .C(_05050_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18379_ (.A1(net2171),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_05051_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18380_ (.A1(_01032_),
    .A2(_01034_),
    .A3(_01039_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18381_ (.A1(_04924_),
    .A2(_04971_),
    .B(_04974_),
    .C(_05053_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18382_ (.A1(_01035_),
    .A2(net1438),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18383_ (.A1(net1424),
    .A2(_05055_),
    .B(net1425),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18384_ (.A1(_05054_),
    .A2(_05056_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18385_ (.A1(net1422),
    .A2(_05057_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18386_ (.I0(_00975_),
    .I1(_05058_),
    .S(_04683_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18387_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(_05059_),
    .S(net1718),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18388_ (.I0(_05052_),
    .I1(_05060_),
    .S(net1815),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18389_ (.A1(net1782),
    .A2(_05049_),
    .B(_05061_),
    .C(_10565_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18390_ (.I0(net41),
    .I1(net54),
    .I2(\load_store_unit_i.rdata_q[18] ),
    .I3(net33),
    .S0(net1886),
    .S1(net1887),
    .Z(_05063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18391_ (.A1(net1833),
    .A2(_05063_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18392_ (.A1(net1507),
    .A2(net1369),
    .B(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2299 (.I(net1449),
    .Z(net2298));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2467 (.I(net2468),
    .Z(net2466));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18395_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .I1(net1368),
    .S(net1498),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18396_ (.I0(_04615_),
    .I1(_04839_),
    .S(_04653_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18397_ (.I0(_04848_),
    .I1(_05068_),
    .S(_04583_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18398_ (.A1(_01276_),
    .A2(net1587),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18399_ (.A1(_01272_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01273_),
    .C(_05070_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18400_ (.A1(net1436),
    .A2(_04660_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18401_ (.A1(_04737_),
    .A2(_05071_),
    .B(_05072_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18402_ (.A1(net1439),
    .A2(_01035_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu9t5v0__and4_4 _18403_ (.A1(net1424),
    .A2(_04954_),
    .A3(_04957_),
    .A4(_05074_),
    .Z(_05075_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18404_ (.A1(_01040_),
    .A2(net1438),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18405_ (.A1(_01035_),
    .A2(_01040_),
    .A3(_01032_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18406_ (.A1(_05076_),
    .A2(_05077_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18407_ (.A1(net1425),
    .A2(_05075_),
    .A3(_05078_),
    .Z(_05079_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18408_ (.A1(net1422),
    .A2(_05079_),
    .B(net1423),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18409_ (.A1(net1420),
    .A2(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18410_ (.I0(_00980_),
    .I1(_05081_),
    .S(_04683_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18411_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(_05082_),
    .S(net1718),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18412_ (.I0(_05073_),
    .I1(_05083_),
    .S(net1815),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18413_ (.A1(net1782),
    .A2(_05069_),
    .B(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18414_ (.A1(_09585_),
    .A2(_04693_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18415_ (.I0(net42),
    .I1(net57),
    .I2(\load_store_unit_i.rdata_q[19] ),
    .I3(net34),
    .S0(net1886),
    .S1(net1887),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18416_ (.A1(net1833),
    .A2(_05087_),
    .B(_04984_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18417_ (.A1(_09585_),
    .A2(_10585_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18418_ (.I0(_05088_),
    .I1(_05089_),
    .S(net1507),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18419_ (.A1(_05085_),
    .A2(_05086_),
    .B(_05090_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1390 (.I(_03490_),
    .Z(net1389));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18421_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .I1(net1366),
    .S(_04697_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18422_ (.A1(_01283_),
    .A2(net1587),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18423_ (.A1(_01279_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01280_),
    .C(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18424_ (.A1(_04737_),
    .A2(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18425_ (.A1(net2278),
    .A2(_04660_),
    .B(_05095_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18426_ (.I(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18427_ (.A1(_01046_),
    .A2(net1420),
    .A3(net1419),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18428_ (.A1(_01052_),
    .A2(_01058_),
    .A3(_01045_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18429_ (.A1(net1419),
    .A2(_01051_),
    .B(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18430_ (.A1(_05054_),
    .A2(_05056_),
    .A3(_05098_),
    .B(_05100_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18431_ (.I(_01046_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18432_ (.I(net1423),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18433_ (.A1(_05102_),
    .A2(_05057_),
    .B(_05103_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18434_ (.A1(net1420),
    .A2(_05104_),
    .B(net1421),
    .C(net1419),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18435_ (.A1(net1390),
    .A2(_05105_),
    .B(_04683_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18436_ (.A1(_00981_),
    .A2(_04683_),
    .B(_05106_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18437_ (.I0(_05097_),
    .I1(_05107_),
    .S(net1718),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18438_ (.I0(_05096_),
    .I1(_05108_),
    .S(net1815),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18439_ (.A1(_04912_),
    .A2(_04825_),
    .B(_05109_),
    .C(_10622_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18440_ (.A1(net1615),
    .A2(_04815_),
    .B(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18441_ (.I0(net44),
    .I1(net58),
    .I2(\load_store_unit_i.rdata_q[20] ),
    .I3(net35),
    .S0(net1886),
    .S1(net1887),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18442_ (.A1(net1833),
    .A2(_05112_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18443_ (.A1(net1507),
    .A2(net1361),
    .B(_05113_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2468 (.I(net2465),
    .Z(net2467));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18445_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .I1(net1354),
    .S(_04697_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18446_ (.A1(_01290_),
    .A2(net1587),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18447_ (.A1(_01286_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01287_),
    .C(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _18448_ (.A1(_09015_),
    .A2(net1434),
    .A3(_04736_),
    .B1(_04737_),
    .B2(_05117_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18449_ (.I(net1421),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18450_ (.A1(net1425),
    .A2(net1423),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18451_ (.I(net1420),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18452_ (.A1(_05102_),
    .A2(_05103_),
    .B(_05121_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _18453_ (.A1(_05075_),
    .A2(_05078_),
    .A3(_05120_),
    .B(_05122_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18454_ (.A1(_05119_),
    .A2(_05123_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18455_ (.A1(net1419),
    .A2(_05124_),
    .B(_01057_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18456_ (.A1(net1417),
    .A2(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18457_ (.I0(_00985_),
    .I1(_05126_),
    .S(_04683_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18458_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(_05127_),
    .S(net1718),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18459_ (.I0(_05118_),
    .I1(_05128_),
    .S(net1815),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18460_ (.A1(_04617_),
    .A2(_04765_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18461_ (.A1(_04667_),
    .A2(_04760_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18462_ (.A1(_04667_),
    .A2(_05130_),
    .B(_05131_),
    .C(_04609_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _18463_ (.A1(_10645_),
    .A2(net1508),
    .A3(_05129_),
    .A4(_05132_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18464_ (.I0(net45),
    .I1(net59),
    .I2(\load_store_unit_i.rdata_q[21] ),
    .I3(net36),
    .S0(net1886),
    .S1(net1887),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18465_ (.A1(net1833),
    .A2(_05134_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18466_ (.A1(_04986_),
    .A2(_04984_),
    .A3(_05135_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18467_ (.A1(_05133_),
    .A2(_05136_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2469 (.I(\core_clock_gate_i.en_latch ),
    .Z(net2468));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18469_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .I1(net1360),
    .S(net1497),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18470_ (.I0(_04722_),
    .I1(_04735_),
    .S(_04583_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18471_ (.A1(_01297_),
    .A2(net1587),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18472_ (.A1(_01293_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01294_),
    .C(_05140_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18473_ (.A1(net1432),
    .A2(_04660_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18474_ (.A1(_04737_),
    .A2(_05141_),
    .B(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18475_ (.A1(_01057_),
    .A2(net1390),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18476_ (.A1(net1417),
    .A2(_05144_),
    .B(net1418),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18477_ (.A1(net1415),
    .A2(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18478_ (.I0(_00992_),
    .I1(_05146_),
    .S(_04683_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18479_ (.I0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .I1(_05147_),
    .S(net1718),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18480_ (.I0(_05143_),
    .I1(_05148_),
    .S(net1815),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _18481_ (.A1(net1782),
    .A2(_05139_),
    .B(_10662_),
    .C(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18482_ (.I0(net46),
    .I1(net60),
    .I2(\load_store_unit_i.rdata_q[22] ),
    .I3(net37),
    .S0(net1886),
    .S1(net1887),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18483_ (.A1(_04560_),
    .A2(_05151_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18484_ (.A1(_05150_),
    .A2(net1507),
    .B(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2470 (.I(net2466),
    .Z(net2469));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18486_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .I1(net2471),
    .S(net1498),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18487_ (.I0(_04618_),
    .I1(_04656_),
    .S(net1615),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18488_ (.A1(_01304_),
    .A2(net1587),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18489_ (.A1(_01300_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01301_),
    .C(_05156_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18490_ (.A1(_04442_),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_05157_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18491_ (.A1(net1421),
    .A2(_01057_),
    .A3(net1418),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18492_ (.A1(net1419),
    .A2(_01057_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18493_ (.A1(net1417),
    .A2(_05160_),
    .B(net1418),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18494_ (.A1(_05123_),
    .A2(_05159_),
    .B(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18495_ (.A1(net1415),
    .A2(_05162_),
    .B(net1416),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18496_ (.A1(net1414),
    .A2(_05163_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18497_ (.I0(_00087_),
    .I1(_05164_),
    .S(_04683_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18498_ (.I(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18499_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(_05166_),
    .S(net1718),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18500_ (.I0(_05158_),
    .I1(_05167_),
    .S(net1815),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18501_ (.A1(net1782),
    .A2(_05155_),
    .B(_05168_),
    .C(_10677_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18502_ (.I0(net47),
    .I1(net61),
    .I2(\load_store_unit_i.rdata_q[23] ),
    .I3(net38),
    .S0(net1886),
    .S1(net1887),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18503_ (.A1(_04560_),
    .A2(_05170_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18504_ (.A1(net1507),
    .A2(net1358),
    .B(_05171_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1389 (.I(_04750_),
    .Z(net1388));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18506_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .I1(net1353),
    .S(net1498),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18507_ (.A1(_01057_),
    .A2(_01063_),
    .A3(_01069_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18508_ (.A1(_05101_),
    .A2(_05174_),
    .Z(_05175_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18509_ (.A1(_01064_),
    .A2(_01063_),
    .A3(_01069_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18510_ (.A1(_01070_),
    .A2(_01069_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18511_ (.A1(_05176_),
    .A2(_05177_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18512_ (.A1(net1414),
    .A2(_05175_),
    .A3(_05178_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18513_ (.A1(_01075_),
    .A2(_05179_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18514_ (.A1(_01082_),
    .A2(_05180_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone2471 (.I(_05318_),
    .Z(net2470));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18516_ (.I0(_04682_),
    .I1(_05181_),
    .S(_04683_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18517_ (.I(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18518_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(_05184_),
    .S(net1718),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18519_ (.I0(_04615_),
    .I1(_04623_),
    .S(_04823_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18520_ (.A1(_04805_),
    .A2(_05186_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18521_ (.A1(_01311_),
    .A2(net1587),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18522_ (.A1(_01307_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01308_),
    .C(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18523_ (.A1(_04737_),
    .A2(_05189_),
    .B(net1783),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18524_ (.A1(net2065),
    .A2(_04660_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18525_ (.A1(_10696_),
    .A2(_05187_),
    .A3(_05190_),
    .A4(_05191_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18526_ (.I0(_04641_),
    .I1(_05020_),
    .S(net1703),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18527_ (.I0(_04716_),
    .I1(_05193_),
    .S(net1551),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18528_ (.I0(_04812_),
    .I1(_05194_),
    .S(_04712_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18529_ (.I0(_04602_),
    .I1(_04943_),
    .I2(_05195_),
    .I3(_04944_),
    .S0(_04581_),
    .S1(_04653_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18530_ (.A1(net1615),
    .A2(_05196_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18531_ (.A1(_08187_),
    .A2(_05185_),
    .B1(_05192_),
    .B2(_05197_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18532_ (.I0(_04555_),
    .I1(_04556_),
    .S(net1886),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18533_ (.A1(net1833),
    .A2(_05199_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18534_ (.A1(net1507),
    .A2(net1357),
    .B(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2472 (.I(_05153_),
    .Z(net2471));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18536_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .I1(net1352),
    .S(net1497),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18537_ (.I0(_04699_),
    .I1(_04700_),
    .S(net1886),
    .Z(_05203_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18538_ (.A1(net1833),
    .A2(_05203_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18539_ (.A1(_08043_),
    .A2(_03333_),
    .A3(net1507),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _18540_ (.I(_01088_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18541_ (.A1(_01076_),
    .A2(_01082_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18542_ (.A1(_01075_),
    .A2(_01082_),
    .B(_01081_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18543_ (.A1(net1380),
    .A2(net1403),
    .B(net1402),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18544_ (.A1(net1404),
    .A2(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18545_ (.I0(_04745_),
    .I1(_05210_),
    .S(_04683_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18546_ (.A1(_07579_),
    .A2(net1815),
    .A3(_05211_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18547_ (.A1(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .A2(net1750),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18548_ (.A1(_01318_),
    .A2(net1587),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18549_ (.A1(_01314_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01315_),
    .C(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18550_ (.A1(net1431),
    .A2(_04660_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18551_ (.A1(_04737_),
    .A2(_05215_),
    .B(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18552_ (.I0(_04621_),
    .I1(_04615_),
    .S(_04729_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18553_ (.I0(_04640_),
    .I1(_04649_),
    .I2(_05021_),
    .I3(_04643_),
    .S0(_04607_),
    .S1(_04712_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18554_ (.I0(_04731_),
    .I1(_05218_),
    .I2(_05219_),
    .I3(_04916_),
    .S0(_04581_),
    .S1(_04653_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18555_ (.I0(_04615_),
    .I1(_04708_),
    .S(_04823_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18556_ (.A1(net1783),
    .A2(_05217_),
    .B1(_05220_),
    .B2(net1615),
    .C1(_05221_),
    .C2(_04723_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18557_ (.A1(_05086_),
    .A2(_05212_),
    .A3(_05213_),
    .A4(_05222_),
    .Z(_05223_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18558_ (.A1(_05204_),
    .A2(_05205_),
    .A3(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1388 (.I(_06458_),
    .Z(net1387));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18560_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .I1(net1356),
    .S(net1498),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18561_ (.I0(net1692),
    .I1(_01319_),
    .S(_04636_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18562_ (.I0(_05019_),
    .I1(_05226_),
    .S(net1703),
    .Z(_05227_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18563_ (.I0(_04715_),
    .I1(_04716_),
    .I2(_05193_),
    .I3(_05227_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18564_ (.I0(_04763_),
    .I1(_05228_),
    .S(_04653_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18565_ (.I0(_04890_),
    .I1(_05229_),
    .S(_04612_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18566_ (.I0(_04615_),
    .I1(_04757_),
    .S(_04823_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18567_ (.I0(_05230_),
    .I1(_05231_),
    .S(_04583_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18568_ (.A1(_01325_),
    .A2(net1587),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18569_ (.A1(_01321_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01322_),
    .C(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18570_ (.A1(net2293),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_05234_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18571_ (.I(_01087_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _18572_ (.A1(_05206_),
    .A2(_05208_),
    .B(_05236_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18573_ (.A1(_05206_),
    .A2(_05207_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18574_ (.A1(_05175_),
    .A2(_05178_),
    .A3(_05238_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18575_ (.A1(net1400),
    .A2(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18576_ (.A1(net1413),
    .A2(_05240_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18577_ (.I0(_04771_),
    .I1(_05241_),
    .S(_04683_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18578_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(_05242_),
    .S(net1718),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18579_ (.I0(_05235_),
    .I1(_05243_),
    .S(net1815),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18580_ (.A1(net1782),
    .A2(_05232_),
    .B(_05244_),
    .C(_10733_),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18581_ (.I0(_04753_),
    .I1(_04754_),
    .S(net1886),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18582_ (.A1(net1833),
    .A2(_05246_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18583_ (.A1(net1355),
    .A2(_04986_),
    .B(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 clone2473 (.I(_05153_),
    .Z(net2472));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18585_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .I1(net1351),
    .S(_04697_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18586_ (.I(_04794_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18587_ (.A1(net1415),
    .A2(_01094_),
    .A3(_05238_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18588_ (.A1(_05123_),
    .A2(_05159_),
    .B(_05161_),
    .C(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18589_ (.A1(_01094_),
    .A2(_05237_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18590_ (.A1(_01094_),
    .A2(net1416),
    .A3(_05238_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18591_ (.A1(_05253_),
    .A2(_05254_),
    .Z(_05255_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18592_ (.A1(_01093_),
    .A2(_05252_),
    .A3(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18593_ (.A1(_01100_),
    .A2(_05256_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18594_ (.A1(_04683_),
    .A2(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18595_ (.A1(_04683_),
    .A2(_05250_),
    .B(_05258_),
    .C(net1718),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18596_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(net1718),
    .B(_05259_),
    .C(net1815),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18597_ (.A1(_01328_),
    .A2(net1614),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18598_ (.A1(_01329_),
    .A2(net1578),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18599_ (.A1(_01332_),
    .A2(net1587),
    .B(_05261_),
    .C(_05262_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18600_ (.A1(net1429),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18601_ (.A1(net1815),
    .A2(_05264_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18602_ (.A1(_04583_),
    .A2(_05018_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18603_ (.A1(_04583_),
    .A2(_05028_),
    .B(_05266_),
    .C(net1782),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18604_ (.A1(_10753_),
    .A2(net1507),
    .A3(_05265_),
    .A4(_05267_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18605_ (.I0(_04785_),
    .I1(_04786_),
    .S(net1886),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18606_ (.A1(net1833),
    .A2(_05269_),
    .B(_04984_),
    .C(_04986_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18607_ (.A1(_05260_),
    .A2(_05268_),
    .B(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2477 (.I(net1630),
    .Z(net2476));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18609_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .I1(net1364),
    .S(net1498),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18610_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(_00985_),
    .S(_04684_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18611_ (.A1(_01178_),
    .A2(net1587),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18612_ (.A1(_01174_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01175_),
    .C(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18613_ (.A1(net1499),
    .A2(_04660_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18614_ (.A1(_04737_),
    .A2(_05275_),
    .B(_05276_),
    .C(net1783),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18615_ (.A1(net1783),
    .A2(_05273_),
    .B(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18616_ (.A1(_10939_),
    .A2(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18617_ (.A1(_04723_),
    .A2(_05230_),
    .B1(_05231_),
    .B2(net1615),
    .C(_05279_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18618_ (.A1(net1886),
    .A2(_04860_),
    .A3(net45),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18619_ (.A1(_04557_),
    .A2(net1887),
    .A3(net36),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18620_ (.A1(_05281_),
    .A2(_05282_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18621_ (.A1(\load_store_unit_i.rdata_q[5] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[13] ),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18622_ (.I0(_05283_),
    .I1(_05284_),
    .S(net1833),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18623_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net53),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18624_ (.A1(_05037_),
    .A2(_05286_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18625_ (.A1(net59),
    .A2(_04870_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18626_ (.A1(_04694_),
    .A2(_05285_),
    .A3(_05287_),
    .A4(_05288_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18627_ (.A1(net1507),
    .A2(_05280_),
    .B(_05289_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 clone2474 (.I(_05153_),
    .Z(net2473));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18629_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net1496),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18630_ (.A1(_01339_),
    .A2(net1587),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18631_ (.A1(_01335_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01336_),
    .C(_05292_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18632_ (.A1(net2138),
    .A2(_04660_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18633_ (.A1(_04737_),
    .A2(_05293_),
    .B(_05294_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18634_ (.I0(_04615_),
    .I1(_04820_),
    .S(_04612_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18635_ (.A1(_08272_),
    .A2(_08293_),
    .B(_04636_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18636_ (.A1(net1676),
    .A2(net1616),
    .B(net1703),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18637_ (.A1(_01326_),
    .A2(net1616),
    .B(net1612),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18638_ (.A1(_05297_),
    .A2(_05298_),
    .B1(_05299_),
    .B2(_05024_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18639_ (.I0(_05227_),
    .I1(_05300_),
    .S(net1551),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18640_ (.I0(_04812_),
    .I1(_04813_),
    .I2(_05301_),
    .I3(_05194_),
    .S0(_04600_),
    .S1(_04612_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18641_ (.I0(_04615_),
    .I1(_04839_),
    .I2(_05296_),
    .I3(_05302_),
    .S0(_03396_),
    .S1(_04653_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18642_ (.I(net1412),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18643_ (.A1(_01094_),
    .A2(_01100_),
    .A3(_05238_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18644_ (.A1(_05174_),
    .A2(_05101_),
    .B(_05178_),
    .C(_05305_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18645_ (.A1(_01094_),
    .A2(_01100_),
    .A3(_05237_),
    .Z(_05307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18646_ (.A1(_01100_),
    .A2(_01093_),
    .B(_05307_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18647_ (.A1(_05304_),
    .A2(_05306_),
    .A3(_05308_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18648_ (.A1(_01106_),
    .A2(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18649_ (.I0(_04853_),
    .I1(_05310_),
    .S(_04683_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18650_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(_05311_),
    .S(net1718),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18651_ (.A1(net1815),
    .A2(_05312_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _18652_ (.A1(net1783),
    .A2(_05295_),
    .B1(_05303_),
    .B2(net1782),
    .C(_05313_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _18653_ (.I0(_10770_),
    .I1(_05314_),
    .S(_09585_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18654_ (.I0(_04832_),
    .I1(_04833_),
    .S(net1886),
    .Z(_05316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18655_ (.A1(net1833),
    .A2(_05316_),
    .B(_04984_),
    .C(net1507),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _18656_ (.A1(_05315_),
    .A2(net1507),
    .B(_05317_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clone2495 (.I(_05318_),
    .Z(net2494));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2484 (.I(net1817),
    .Z(net2483));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18659_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .I1(net1350),
    .S(_04697_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18660_ (.A1(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .A2(net1750),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18661_ (.A1(_01093_),
    .A2(_01099_),
    .A3(_01105_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18662_ (.A1(_01100_),
    .A2(_01099_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18663_ (.A1(_01106_),
    .A2(_05323_),
    .B(_01105_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18664_ (.I(_05324_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18665_ (.A1(_05255_),
    .A2(_05252_),
    .A3(_05322_),
    .B(_05325_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _18666_ (.A1(_01112_),
    .A2(_05326_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18667_ (.I0(_04885_),
    .I1(_05327_),
    .S(_04683_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18668_ (.A1(net1750),
    .A2(_05328_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18669_ (.A1(_05321_),
    .A2(_05329_),
    .B(net1815),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18670_ (.I0(_04615_),
    .I1(_04762_),
    .S(_04823_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18671_ (.A1(_01346_),
    .A2(net1587),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18672_ (.A1(_01342_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01343_),
    .C(_05332_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18673_ (.A1(_04737_),
    .A2(_05333_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18674_ (.A1(net1408),
    .A2(_04660_),
    .B1(_05331_),
    .B2(_04805_),
    .C(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18675_ (.A1(_08265_),
    .A2(_08267_),
    .B(_04636_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18676_ (.A1(net1675),
    .A2(net1616),
    .B(net1703),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18677_ (.A1(net1676),
    .A2(net1616),
    .B(net1612),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18678_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_05338_),
    .B2(_05297_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18679_ (.I0(_04643_),
    .I1(_05021_),
    .I2(_05026_),
    .I3(_05339_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18680_ (.I0(_04757_),
    .I1(_04759_),
    .I2(_04758_),
    .I3(_05340_),
    .S0(_04653_),
    .S1(_04612_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18681_ (.A1(net1615),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18682_ (.A1(_05335_),
    .A2(_05342_),
    .B(_04997_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18683_ (.A1(_10787_),
    .A2(net1508),
    .A3(_05343_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18684_ (.I0(net53),
    .I1(net36),
    .I2(net59),
    .I3(net45),
    .S0(net1886),
    .S1(net1887),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18685_ (.A1(net1833),
    .A2(_05345_),
    .B(_04984_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18686_ (.A1(_05330_),
    .A2(_05344_),
    .B1(_05346_),
    .B2(_04694_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2483 (.I(_01264_),
    .Z(net2482));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18688_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .I1(net1363),
    .S(_04697_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18689_ (.I0(_04900_),
    .I1(_04901_),
    .S(net1886),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18690_ (.A1(_04560_),
    .A2(_05349_),
    .B(_04984_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18691_ (.A1(_08050_),
    .A2(_08077_),
    .B(_04636_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18692_ (.A1(_01347_),
    .A2(net1616),
    .B(net1703),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18693_ (.A1(net1675),
    .A2(net1616),
    .B(net1612),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18694_ (.A1(_05351_),
    .A2(_05352_),
    .B1(_05353_),
    .B2(_05336_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18695_ (.I0(_05193_),
    .I1(_05227_),
    .I2(_05300_),
    .I3(_05354_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18696_ (.I0(_04708_),
    .I1(_04714_),
    .I2(_04720_),
    .I3(_05355_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18697_ (.A1(_04578_),
    .A2(_04581_),
    .A3(_04729_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18698_ (.I0(_04621_),
    .I1(_04615_),
    .S(_05357_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18699_ (.A1(_01353_),
    .A2(net1587),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18700_ (.A1(_01349_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01350_),
    .C(_05359_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18701_ (.A1(net2122),
    .A2(_04660_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18702_ (.A1(_04737_),
    .A2(_05360_),
    .B(_05361_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18703_ (.A1(net1615),
    .A2(_05356_),
    .B1(_05358_),
    .B2(_04723_),
    .C(_05362_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18704_ (.A1(net1815),
    .A2(_05363_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18705_ (.A1(net1412),
    .A2(_01105_),
    .A3(_01111_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _18706_ (.A1(_05306_),
    .A2(_05308_),
    .A3(_05365_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18707_ (.A1(_01106_),
    .A2(_01105_),
    .A3(_01111_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18708_ (.A1(_01112_),
    .A2(_01111_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18709_ (.A1(_05367_),
    .A2(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18710_ (.A1(net1411),
    .A2(_05366_),
    .A3(_05369_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18711_ (.A1(_05366_),
    .A2(_05369_),
    .B(net1411),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18712_ (.A1(_05370_),
    .A2(_05371_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18713_ (.I0(_04926_),
    .I1(_05372_),
    .S(_04683_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18714_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(_05373_),
    .S(net1718),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18715_ (.A1(net1815),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18716_ (.A1(_10810_),
    .A2(net1507),
    .A3(_05364_),
    .A4(_05375_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18717_ (.A1(net1508),
    .A2(_05350_),
    .B(_05376_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2481 (.I(_06392_),
    .Z(net2480));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18719_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .I1(net1349),
    .S(net1498),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18720_ (.I0(_04936_),
    .I1(_04937_),
    .S(net1886),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18721_ (.A1(_04560_),
    .A2(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18722_ (.A1(_04986_),
    .A2(_04984_),
    .A3(_05380_),
    .Z(_05381_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18723_ (.A1(_10159_),
    .A2(_10839_),
    .B1(_10840_),
    .B2(net1560),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18724_ (.A1(net1562),
    .A2(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18725_ (.A1(\cs_registers_i.dscratch0_q[31] ),
    .A2(net1556),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _18726_ (.A1(\cs_registers_i.dscratch1_q[31] ),
    .A2(_10188_),
    .B1(_10239_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .C1(net91),
    .C2(net1563),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18727_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_10197_),
    .B(_10245_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _18728_ (.A1(_05383_),
    .A2(_05384_),
    .A3(_05385_),
    .A4(_05386_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18729_ (.A1(_01112_),
    .A2(_01118_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18730_ (.A1(_01118_),
    .A2(_01111_),
    .B(_01117_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18731_ (.A1(_05326_),
    .A2(_05388_),
    .B(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _18732_ (.A1(_01124_),
    .A2(_05390_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18733_ (.I0(_04960_),
    .I1(_05391_),
    .S(_04683_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _18734_ (.A1(net1750),
    .A2(_05392_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18735_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net1750),
    .B(net1783),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18736_ (.I0(_04615_),
    .I1(_04943_),
    .S(_04823_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18737_ (.A1(_09470_),
    .A2(_04636_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _18738_ (.A1(_08082_),
    .A2(_08099_),
    .A3(_04636_),
    .B(net1703),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18739_ (.A1(_01347_),
    .A2(net1616),
    .B(net1612),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18740_ (.A1(_05396_),
    .A2(_05397_),
    .B1(_05398_),
    .B2(_05351_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18741_ (.I0(_05021_),
    .I1(_05026_),
    .I2(_05339_),
    .I3(_05399_),
    .S0(net1551),
    .S1(_04712_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _18742_ (.I0(_04623_),
    .I1(_04635_),
    .I2(_04651_),
    .I3(_05400_),
    .S0(_04612_),
    .S1(_04653_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18743_ (.A1(_04583_),
    .A2(_05401_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18744_ (.A1(net1615),
    .A2(_05395_),
    .B(_05402_),
    .C(net1782),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18745_ (.A1(_00944_),
    .A2(net1587),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18746_ (.A1(_00940_),
    .A2(net1614),
    .B1(net1578),
    .B2(_00941_),
    .C(_05404_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18747_ (.A1(_04737_),
    .A2(_05405_),
    .B(net1783),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18748_ (.A1(net2051),
    .A2(_04660_),
    .B(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18749_ (.A1(_05393_),
    .A2(_05394_),
    .B1(_05403_),
    .B2(_05407_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _18750_ (.A1(_10825_),
    .A2(_05387_),
    .A3(net1508),
    .A4(_05408_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _18751_ (.A1(_05381_),
    .A2(_05409_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2480 (.I(net1768),
    .Z(net2479));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18753_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .I1(net1348),
    .S(_04697_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18754_ (.I0(_05220_),
    .I1(_05221_),
    .S(net1615),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18755_ (.A1(_01185_),
    .A2(net1587),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18756_ (.A1(_01181_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01182_),
    .C(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18757_ (.A1(_04737_),
    .A2(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18758_ (.A1(net1500),
    .A2(_04660_),
    .B(_05415_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18759_ (.I(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18760_ (.I0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .I1(_00992_),
    .S(_04684_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18761_ (.I0(_05417_),
    .I1(_05418_),
    .S(net1815),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18762_ (.A1(net1782),
    .A2(_05412_),
    .B(_05419_),
    .C(_10954_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18763_ (.A1(net1886),
    .A2(_04860_),
    .A3(net46),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18764_ (.A1(_04557_),
    .A2(net1887),
    .A3(net37),
    .Z(_05422_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18765_ (.A1(_05421_),
    .A2(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18766_ (.A1(\load_store_unit_i.rdata_q[6] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[14] ),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18767_ (.I0(_05423_),
    .I1(_05424_),
    .S(_04560_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18768_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net55),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[22] ),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18769_ (.A1(_05037_),
    .A2(_05426_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18770_ (.A1(net60),
    .A2(_04870_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18771_ (.A1(_04694_),
    .A2(_05425_),
    .A3(_05427_),
    .A4(_05428_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18772_ (.A1(net1507),
    .A2(_05420_),
    .B(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2479 (.I(_06391_),
    .Z(net2478));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18774_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net1496),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18775_ (.A1(_04723_),
    .A2(_05196_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18776_ (.A1(_01192_),
    .A2(net1587),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18777_ (.A1(_01188_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01189_),
    .C(_05433_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18778_ (.A1(net1512),
    .A2(_04660_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18779_ (.A1(_04737_),
    .A2(_05434_),
    .B(_05435_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18780_ (.I(_00087_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18781_ (.I0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .I1(_05437_),
    .S(_04684_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18782_ (.I0(_05436_),
    .I1(_05438_),
    .S(net1815),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18783_ (.A1(net1615),
    .A2(_05186_),
    .B(_05439_),
    .C(_10982_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18784_ (.A1(_05432_),
    .A2(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18785_ (.A1(_04860_),
    .A2(_04873_),
    .A3(\load_store_unit_i.rdata_q[15] ),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18786_ (.A1(net1887),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .B(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18787_ (.A1(_04860_),
    .A2(net47),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18788_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(\load_store_unit_i.rdata_q[23] ),
    .B1(net56),
    .B2(\load_store_unit_i.data_type_q[1] ),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _18789_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(_05443_),
    .B1(_05444_),
    .B2(_04560_),
    .C1(_05445_),
    .C2(_04860_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18790_ (.I0(net38),
    .I1(\load_store_unit_i.rdata_q[7] ),
    .S(_04560_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18791_ (.I0(net61),
    .I1(_05447_),
    .S(net1887),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18792_ (.I0(_05446_),
    .I1(_05448_),
    .S(_04557_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18793_ (.I0(_05441_),
    .I1(_05449_),
    .S(net1508),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 clone2478 (.I(_09871_),
    .Z(net2477));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18795_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net1496),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1387 (.I(_06502_),
    .Z(net1386));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18797_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net1496),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1386 (.I(_06502_),
    .Z(net1385));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18799_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net1496),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2494 (.I(_00449_),
    .Z(net2493));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18801_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net1496),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2485 (.I(_00865_),
    .Z(net2484));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18803_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net1496),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2493 (.I(_00449_),
    .Z(net2492));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18805_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net1496),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2492 (.I(_05208_),
    .Z(net2491));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18807_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net1496),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1385 (.I(_06506_),
    .Z(net1384));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1384 (.I(_06506_),
    .Z(net1383));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18810_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net1496),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2496 (.I(_09837_),
    .Z(net2495));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18812_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net1496),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1383 (.I(_06679_),
    .Z(net1382));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18814_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net1496),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18816_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net1496),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1381 (.I(_05163_),
    .Z(net1380));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18818_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net1496),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1380 (.I(_05497_),
    .Z(net1379));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18820_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .S(net1496),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18822_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net1496),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1382 (.I(_04782_),
    .Z(net1381));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18824_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net1496),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1379 (.I(_06489_),
    .Z(net1378));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18826_ (.I0(net1359),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net1496),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18828_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net1496),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1378 (.I(_04898_),
    .Z(net1377));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18831_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net1496),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1377 (.I(_04830_),
    .Z(net1376));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18833_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net1496),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1376 (.I(_04858_),
    .Z(net1375));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18835_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net1496),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1375 (.I(_04964_),
    .Z(net1374));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18837_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net1496),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1373 (.I(_05107_),
    .Z(net1372));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18839_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net1496),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1372 (.I(_04931_),
    .Z(net1371));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18841_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net1496),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1371 (.I(_04989_),
    .Z(net1370));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18843_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net1496),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1370 (.I(_05062_),
    .Z(net1369));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18845_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net1496),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18846_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(_00972_),
    .S(_04684_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18847_ (.A1(_08127_),
    .A2(_03412_),
    .A3(_03422_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18848_ (.A1(_01144_),
    .A2(net1587),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18849_ (.A1(_01141_),
    .A2(net1614),
    .B1(net1578),
    .B2(_01142_),
    .C(_05480_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18850_ (.A1(net1540),
    .A2(_04736_),
    .B1(_04737_),
    .B2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18851_ (.A1(_04723_),
    .A2(_05401_),
    .B1(_05395_),
    .B2(net1615),
    .C(_05482_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18852_ (.A1(_03424_),
    .A2(_03427_),
    .B(_08127_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18853_ (.A1(_03402_),
    .A2(_05479_),
    .B(_05483_),
    .C(_05484_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18854_ (.A1(_09585_),
    .A2(net1783),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18855_ (.A1(net1815),
    .A2(_05478_),
    .B1(_05485_),
    .B2(_05486_),
    .C(_10223_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18856_ (.A1(_04860_),
    .A2(net32),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18857_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net48),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[16] ),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18858_ (.A1(net1886),
    .A2(_04860_),
    .A3(net39),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18859_ (.A1(_04557_),
    .A2(net1887),
    .A3(net62),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18860_ (.A1(_05490_),
    .A2(_05491_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18861_ (.A1(\load_store_unit_i.rdata_q[0] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[8] ),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18862_ (.I0(_05492_),
    .I1(_05493_),
    .S(_04560_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _18863_ (.A1(net1886),
    .A2(_05488_),
    .B1(_05037_),
    .B2(_05489_),
    .C(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18864_ (.A1(_04694_),
    .A2(_05495_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18865_ (.A1(net1508),
    .A2(_05487_),
    .B(_05496_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1368 (.I(_05008_),
    .Z(net1367));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _18867_ (.I(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18868_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(_05499_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _18869_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_09520_),
    .A3(_05044_),
    .A4(_05500_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1367 (.I(_05091_),
    .Z(net1366));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18871_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .I1(net1379),
    .S(net1505),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18872_ (.A1(\load_store_unit_i.rdata_q[1] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[9] ),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18873_ (.A1(net1886),
    .A2(_04860_),
    .A3(net40),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18874_ (.A1(net63),
    .A2(_04862_),
    .B(_05504_),
    .C(_04560_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18875_ (.A1(_04560_),
    .A2(_05503_),
    .B(_05505_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18876_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net49),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[17] ),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _18877_ (.A1(_04860_),
    .A2(_05507_),
    .B(net1886),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18878_ (.I0(net43),
    .I1(_05506_),
    .S(net1887),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _18879_ (.A1(_05506_),
    .A2(_05508_),
    .B1(_05509_),
    .B2(net1886),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18880_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(_00974_),
    .S(_04684_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18881_ (.A1(_08187_),
    .A2(_05511_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18882_ (.A1(_04583_),
    .A2(_05356_),
    .Z(_05513_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18883_ (.A1(net1615),
    .A2(_05358_),
    .B(_05513_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18884_ (.A1(_01147_),
    .A2(net1614),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18885_ (.A1(_01148_),
    .A2(net1578),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18886_ (.A1(_01150_),
    .A2(net1587),
    .B(_05515_),
    .C(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18887_ (.A1(net1539),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_05517_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18888_ (.A1(_04609_),
    .A2(_05514_),
    .B(_05518_),
    .C(net1783),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _18889_ (.A1(_05512_),
    .A2(_05519_),
    .B(_10605_),
    .C(net1508),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18890_ (.A1(net1508),
    .A2(_05510_),
    .B(_05520_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 clone2475 (.I(_09751_),
    .Z(net2474));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18892_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .I1(net1453),
    .S(net1505),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18893_ (.A1(\load_store_unit_i.rdata_q[2] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[10] ),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18894_ (.A1(net1886),
    .A2(_04860_),
    .A3(net41),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18895_ (.A1(_04557_),
    .A2(net1887),
    .A3(net33),
    .Z(_05525_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _18896_ (.A1(net1833),
    .A2(_05524_),
    .A3(_05525_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18897_ (.A1(net1833),
    .A2(_05523_),
    .B(_05526_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18898_ (.A1(_04557_),
    .A2(_04860_),
    .A3(net54),
    .Z(_05528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18899_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net50),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[18] ),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18900_ (.A1(_05037_),
    .A2(_05529_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _18901_ (.A1(_04986_),
    .A2(_05527_),
    .A3(_05528_),
    .A4(_05530_),
    .Z(_05531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18902_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(_00975_),
    .S(_04684_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18903_ (.A1(_08187_),
    .A2(_05532_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18904_ (.A1(_01153_),
    .A2(net1614),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18905_ (.A1(_01154_),
    .A2(net1578),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18906_ (.A1(_01157_),
    .A2(net1587),
    .B(_05534_),
    .C(_05535_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18907_ (.A1(net1521),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _18908_ (.A1(_04762_),
    .A2(_04823_),
    .B(_04583_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18909_ (.A1(net1615),
    .A2(_05341_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _18910_ (.A1(_04609_),
    .A2(_05538_),
    .A3(_05539_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18911_ (.A1(net1783),
    .A2(_05537_),
    .A3(_05540_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18912_ (.A1(_05533_),
    .A2(_05541_),
    .B(_10257_),
    .C(net1507),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _18913_ (.A1(_05531_),
    .A2(_05542_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1365 (.I(_05271_),
    .Z(net1364));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18915_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .I1(_05543_),
    .S(net1505),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18916_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net51),
    .B1(_04874_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18917_ (.A1(net57),
    .A2(_04870_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18918_ (.A1(net1886),
    .A2(_04860_),
    .A3(net42),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _18919_ (.A1(_04557_),
    .A2(net1887),
    .A3(net34),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _18920_ (.A1(_05547_),
    .A2(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _18921_ (.A1(\load_store_unit_i.rdata_q[3] ),
    .A2(_04862_),
    .B1(_04864_),
    .B2(\load_store_unit_i.rdata_q[11] ),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18922_ (.I0(_05549_),
    .I1(_05550_),
    .S(net1833),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18923_ (.A1(_05037_),
    .A2(_05545_),
    .B(_05546_),
    .C(_05551_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18924_ (.I0(_10889_),
    .I1(_05552_),
    .S(net1508),
    .Z(_05553_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18925_ (.A1(_04653_),
    .A2(_05296_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18926_ (.A1(_01160_),
    .A2(net1614),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _18927_ (.A1(_01161_),
    .A2(net1578),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18928_ (.A1(_01164_),
    .A2(net1587),
    .B(_05555_),
    .C(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _18929_ (.A1(net1519),
    .A2(_04660_),
    .B1(_04665_),
    .B2(_05557_),
    .C(net1815),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18930_ (.A1(_04578_),
    .A2(_05302_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18931_ (.A1(_04653_),
    .A2(_04839_),
    .B(_05559_),
    .C(_04805_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _18932_ (.A1(_04583_),
    .A2(_05554_),
    .B(_05558_),
    .C(_05560_),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18933_ (.I0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .I1(_00980_),
    .S(_04684_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18934_ (.A1(_08187_),
    .A2(_05562_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _18935_ (.A1(_09585_),
    .A2(_04986_),
    .A3(_05561_),
    .A4(_05563_),
    .Z(_05564_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _18936_ (.A1(_05553_),
    .A2(_05564_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1364 (.I(_05347_),
    .Z(net1363));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18938_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .I1(_05565_),
    .S(net1506),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1362 (.I(_05111_),
    .Z(net1361));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18940_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .I1(_05042_),
    .S(net1505),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1361 (.I(_05137_),
    .Z(net1360));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18942_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .I1(net1396),
    .S(net1505),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1360 (.I(_05153_),
    .Z(net1359));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18944_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .I1(net1399),
    .S(net1505),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1358 (.I(_05198_),
    .Z(net1357));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18946_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .I1(_05450_),
    .S(net1505),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18947_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .I1(net1392),
    .S(net1506),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18948_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .I1(net1388),
    .S(net1506),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1356 (.I(_05245_),
    .Z(net1355));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18950_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .I1(net1381),
    .S(net1506),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18951_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .I1(net1376),
    .S(net1505),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18952_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .I1(net1375),
    .S(net1506),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18953_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .I1(net1377),
    .S(net1506),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18954_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .I1(net1371),
    .S(net1506),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .I1(net1374),
    .S(net1506),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18956_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .I1(net1370),
    .S(net1506),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18957_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .I1(net1362),
    .S(net1506),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .I1(net1368),
    .S(net1506),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18959_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .I1(net1366),
    .S(net1506),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1355 (.I(_05114_),
    .Z(net1354));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .I1(net1354),
    .S(net1506),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18962_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .I1(net1360),
    .S(net1506),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18963_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .I1(net1359),
    .S(net1506),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18964_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .I1(net1353),
    .S(net1506),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18965_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .I1(net1352),
    .S(net1506),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18966_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .I1(net1356),
    .S(net1506),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18967_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .I1(net1351),
    .S(net1506),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18968_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .I1(net1364),
    .S(net1506),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18969_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .I1(net2494),
    .S(net1506),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18970_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .I1(net1363),
    .S(net1506),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .I1(net1349),
    .S(net1506),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18972_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .I1(net1348),
    .S(net1505),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _18973_ (.A1(_07968_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_05044_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _18974_ (.A1(_05500_),
    .A2(_05573_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1354 (.I(_05172_),
    .Z(net1353));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18976_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .I1(net1379),
    .S(_05574_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18977_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .I1(net1453),
    .S(_05574_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18978_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .I1(_05543_),
    .S(_05574_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18979_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .I1(_05565_),
    .S(net1494),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18980_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .I1(_05042_),
    .S(_05574_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .I1(net1396),
    .S(_05574_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18982_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .I1(net1399),
    .S(_05574_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18983_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .I1(_05450_),
    .S(_05574_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18984_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .I1(net1392),
    .S(net1495),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18985_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .I1(net1388),
    .S(net1494),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1353 (.I(_05201_),
    .Z(net1352));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18987_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .I1(net1381),
    .S(net1494),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18988_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .I1(net1376),
    .S(_05574_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18989_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .I1(net1375),
    .S(net1494),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18990_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .I1(net1377),
    .S(net1494),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18991_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .I1(net1371),
    .S(net1494),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18992_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .I1(net1374),
    .S(net1494),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18993_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .I1(net1370),
    .S(net1494),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18994_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .I1(net1362),
    .S(net1494),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18995_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .I1(net1368),
    .S(net1495),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18996_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .I1(net1366),
    .S(net1495),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1352 (.I(_05248_),
    .Z(net1351));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18998_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .I1(net1354),
    .S(net1495),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18999_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .I1(net1360),
    .S(net1494),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19000_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .I1(net2471),
    .S(net1494),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19001_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .I1(net1353),
    .S(net1494),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19002_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .I1(net1352),
    .S(net1494),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19003_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .I1(net1356),
    .S(net1495),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19004_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .I1(net1351),
    .S(net1495),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19005_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .I1(net1364),
    .S(net1495),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19006_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .I1(net2470),
    .S(net1495),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19007_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .I1(net1363),
    .S(net1495),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19008_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .I1(net1349),
    .S(net1495),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19009_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .I1(net1348),
    .S(_05574_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _19010_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(_09519_),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_05044_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19011_ (.A1(_05500_),
    .A2(_05578_),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place1351 (.I(_05318_),
    .Z(net1350));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19013_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .I1(net1379),
    .S(_05579_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19014_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .I1(net1453),
    .S(_05579_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19015_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .I1(_05543_),
    .S(_05579_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19016_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .I1(_05565_),
    .S(net1493),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19017_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .I1(_05042_),
    .S(_05579_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19018_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .I1(net1396),
    .S(_05579_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19019_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .I1(net1399),
    .S(_05579_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19020_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .I1(_05450_),
    .S(net1493),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19021_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .I1(net1392),
    .S(net1493),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19022_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .I1(net1388),
    .S(_05579_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1350 (.I(_05377_),
    .Z(net1349));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19024_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .I1(net1381),
    .S(net1493),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19025_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .I1(net1376),
    .S(_05579_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19026_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .I1(net1375),
    .S(_05579_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19027_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .I1(net1377),
    .S(_05579_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19028_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .I1(net1371),
    .S(_05579_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19029_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .I1(net1374),
    .S(_05579_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19030_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .I1(net1370),
    .S(net1493),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19031_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .I1(net1362),
    .S(_05579_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19032_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .I1(net1368),
    .S(net1493),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19033_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .I1(net1366),
    .S(net1493),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1359 (.I(_05169_),
    .Z(net1358));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19035_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .I1(net1354),
    .S(net1493),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19036_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .I1(net1360),
    .S(_05579_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19037_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .I1(net2472),
    .S(_05579_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19038_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .I1(net1353),
    .S(net1493),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19039_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .I1(net1352),
    .S(_05579_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19040_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .I1(net1356),
    .S(net1493),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19041_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .I1(net1351),
    .S(net1493),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19042_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .I1(net1364),
    .S(net1493),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19043_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .I1(net2470),
    .S(net1493),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19044_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .I1(net1363),
    .S(net1493),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19045_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .I1(net1349),
    .S(net1493),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19046_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .I1(net1348),
    .S(net1493),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1357 (.I(_05224_),
    .Z(net1356));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19048_ (.A1(_05045_),
    .A2(_05500_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1349 (.I(_05410_),
    .Z(net1348));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19050_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(_05584_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2043 (.I(net146),
    .Z(net2042));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19052_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(net1492),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2028 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Z(net2027));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19054_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(net1492),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2024 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Z(net2023));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19056_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net1492),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19057_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S(net1492),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19058_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S(_05584_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19059_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S(_05584_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19060_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S(net1492),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19061_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S(net1492),
    .Z(_02038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19062_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S(net1492),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2027 (.I(\cs_registers_i.pc_if_i[1] ),
    .Z(net2026));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19064_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S(net1492),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19065_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S(_05584_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19066_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S(net1492),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19067_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S(net1492),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19068_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S(net1492),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19069_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S(net1492),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19070_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(net1492),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19071_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S(net1492),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19072_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S(net1492),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19073_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S(net1492),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2035 (.I(net2033),
    .Z(net2034));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19075_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S(net1492),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19076_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S(net1492),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19077_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S(net1492),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19078_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S(net1492),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19079_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S(net1492),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19080_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S(net1492),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19081_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S(net1492),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19082_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S(net1492),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19083_ (.I0(net2494),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S(net1492),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19084_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S(net1492),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19085_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S(net1492),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19086_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S(net1492),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19087_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A2(_05499_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _19088_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_09520_),
    .A3(_05044_),
    .A4(_05591_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place2022 (.I(\id_stage_i.controller_i.instr_i[12] ),
    .Z(net2021));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19090_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .S(net1504),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19091_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .S(net1504),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19092_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .S(net1504),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19093_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .S(net1504),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19094_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .S(net1504),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19095_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .S(net1504),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19096_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .S(net1504),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19097_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .S(net1504),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19098_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .S(net1504),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19099_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .S(net1504),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place2021 (.I(\id_stage_i.controller_i.instr_i[13] ),
    .Z(net2020));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19101_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .S(net1504),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19102_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .S(net1504),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19103_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .S(net1504),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19104_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .S(net1504),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19105_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .S(net1504),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19106_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .S(net1504),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19107_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .S(net1504),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19108_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .S(net1504),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19109_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .S(net1504),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19110_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .S(net1504),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2046 (.I(net143),
    .Z(net2045));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19112_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .S(net1504),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19113_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .S(net1504),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19114_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .S(net1504),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19115_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .S(net1504),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19116_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .S(net1504),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19117_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .S(net1504),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19118_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .S(net1504),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19119_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .S(net1504),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19120_ (.I0(net2494),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .S(net1504),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19121_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .S(net1504),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19122_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .S(net1504),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19123_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .S(net1504),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19124_ (.A1(_05573_),
    .A2(_05591_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_23_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_23_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19126_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .S(net1491),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19127_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .S(net1491),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19128_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .S(net1491),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19129_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .S(net1491),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19130_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .S(net1491),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19131_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .S(net1491),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19132_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .S(net1491),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19133_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .S(net1491),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19134_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .S(net1491),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19135_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .S(net1491),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1960 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .Z(net1959));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19137_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .S(net1491),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19138_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .S(net1491),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19139_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .S(net1491),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19140_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .S(net1491),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19141_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .S(net1491),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19142_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .S(net1491),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19143_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .S(net1491),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19144_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .S(net1491),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19145_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .S(net1491),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19146_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .S(net1491),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1959 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .Z(net1958));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19148_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .S(net1491),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19149_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .S(net1491),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19150_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .S(net1491),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19151_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .S(net1491),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19152_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .S(net1491),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19153_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .S(net1491),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19154_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .S(net1491),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19155_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .S(net1491),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19156_ (.I0(net2494),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .S(net1491),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19157_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .S(net1491),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19158_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .S(net1491),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19159_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .S(net1491),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19160_ (.A1(_05578_),
    .A2(_05591_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1961 (.I(net1959),
    .Z(net1960));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19162_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .I1(net1379),
    .S(net1490),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19163_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .I1(net1453),
    .S(net1490),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19164_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .I1(_05543_),
    .S(net1490),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19165_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .I1(_05565_),
    .S(net1490),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19166_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .I1(_05042_),
    .S(net1490),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19167_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .I1(net1396),
    .S(net1490),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19168_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .I1(net1399),
    .S(net1490),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19169_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .I1(_05450_),
    .S(net1490),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19170_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .I1(net1392),
    .S(net1490),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19171_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .I1(net1388),
    .S(net1490),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19172_ (.A1(_09518_),
    .A2(_05573_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1975 (.I(net1973),
    .Z(net1974));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19174_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .S(_05602_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1974 (.I(net1972),
    .Z(net1973));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19176_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .I1(net1381),
    .S(net1490),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19177_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .I1(net1376),
    .S(net1490),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19178_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .I1(net1375),
    .S(net1490),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19179_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .I1(net1377),
    .S(net1490),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19180_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .I1(net1371),
    .S(net1490),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19181_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .I1(net1374),
    .S(net1490),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19182_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .I1(net1370),
    .S(net1490),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19183_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .I1(net1362),
    .S(net1490),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19184_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .I1(net1368),
    .S(net1490),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19185_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .I1(net1366),
    .S(net1490),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19186_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .S(_05602_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1973 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net1972));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19188_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .I1(net1354),
    .S(net1490),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19189_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .I1(net1360),
    .S(net1490),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19190_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .I1(net2473),
    .S(net1490),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19191_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .I1(net1353),
    .S(net1490),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19192_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .I1(net1352),
    .S(net1490),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19193_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .I1(net1356),
    .S(net1490),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19194_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .I1(net1351),
    .S(net1490),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19195_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .I1(net1364),
    .S(net1490),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19196_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .I1(net2470),
    .S(net1490),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19197_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .I1(net1363),
    .S(net1490),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19198_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .S(_05602_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19199_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .I1(net1349),
    .S(net1490),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19200_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .I1(net1348),
    .S(net1490),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19201_ (.A1(_05045_),
    .A2(_05591_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1981 (.I(net1976),
    .Z(net1980));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19203_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S(net1488),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19204_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S(net1488),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19205_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S(net1488),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19206_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S(net1488),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19207_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S(net1488),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19208_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S(net1488),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19209_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S(net1488),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19210_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S(net1488),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19211_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .S(net1489),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19212_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S(net1488),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19213_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S(net1488),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1955 (.I(net1944),
    .Z(net1954));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19215_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S(net1488),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19216_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S(net1488),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19217_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S(net1488),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19218_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S(net1488),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19219_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S(net1488),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19220_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S(net1488),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19221_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S(net1488),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19222_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S(net1488),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19223_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .S(_05602_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19224_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S(net1488),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19225_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S(net1488),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1879 (.I(net1877),
    .Z(net1878));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19227_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S(net1488),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19228_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S(net1488),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19229_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S(net1488),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19230_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S(net1488),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19231_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S(net1488),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19232_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S(net1488),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19233_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S(net1488),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19234_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S(net1488),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19235_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .S(_05602_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19236_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S(net1488),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19237_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S(net1488),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19238_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S(net1488),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19239_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S(net1488),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _19240_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A2(_09520_),
    .A3(_04691_),
    .A4(_05044_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1864 (.I(_07657_),
    .Z(net1863));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19242_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .S(net1502),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19243_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .S(net1502),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19244_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .S(net1502),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19245_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .S(net1503),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19246_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .S(net1502),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19247_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .S(net1502),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19248_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .S(_05602_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19249_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .S(net1502),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19250_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .S(net1503),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19251_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .S(net1503),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19252_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .S(net1502),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1927 (.I(net1925),
    .Z(net1926));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19254_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .S(net1502),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19255_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .S(net1502),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19256_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .S(net1502),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19257_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .S(net1503),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19258_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .S(net1502),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19259_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .S(net1503),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19260_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .S(net1489),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19261_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .S(net1503),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19262_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .S(net1502),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19263_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .S(net1503),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19264_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .S(net1503),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1806 (.I(_06492_),
    .Z(net1805));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19266_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .S(net1503),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19267_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .S(net1502),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19268_ (.I0(net2472),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .S(net1502),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19269_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .S(net1503),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19270_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .S(net1502),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19271_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .S(net1503),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19272_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .S(net1489),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19273_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .S(net1503),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19274_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .S(net1503),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19275_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .S(net1503),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19276_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .S(net1503),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19277_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .S(net1503),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19278_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .S(net1503),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19279_ (.A1(_04691_),
    .A2(_05573_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place2009 (.I(net2005),
    .Z(net2008));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19281_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .I1(net1379),
    .S(net1487),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19282_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .I1(net1453),
    .S(net1487),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19283_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .I1(_05543_),
    .S(net1487),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19284_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .I1(_05565_),
    .S(_05614_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19285_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .S(net1489),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19286_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .I1(_05042_),
    .S(net1487),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19287_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .I1(net1396),
    .S(net1487),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19288_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .I1(net1399),
    .S(net1487),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19289_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .I1(_05450_),
    .S(_05614_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19290_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .I1(net1392),
    .S(_05614_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19291_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .I1(net1388),
    .S(net1487),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1750 (.I(_09770_),
    .Z(net1749));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19293_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .I1(net1381),
    .S(net1487),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19294_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .I1(net1376),
    .S(net1487),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19295_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .I1(net1375),
    .S(net1487),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19296_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .I1(net1377),
    .S(net1487),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1661 (.I(_09774_),
    .Z(net1660));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19298_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .S(net1489),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19299_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .I1(net1371),
    .S(net1487),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19300_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .I1(net1374),
    .S(net1487),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19301_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .I1(net1370),
    .S(net1487),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19302_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .I1(net1362),
    .S(net1487),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19303_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .I1(net1368),
    .S(_05614_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19304_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .I1(net1366),
    .S(_05614_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1662 (.I(net1660),
    .Z(net1661));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19306_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .I1(net1354),
    .S(_05614_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19307_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .I1(net1360),
    .S(net1487),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19308_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .I1(net2472),
    .S(net1487),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19309_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .I1(net1353),
    .S(net1487),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19310_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .S(_05602_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19311_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .I1(net1352),
    .S(net1487),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19312_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .I1(net1356),
    .S(_05614_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19313_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .I1(net1351),
    .S(_05614_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19314_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .I1(net1364),
    .S(_05614_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19315_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .I1(net2470),
    .S(_05614_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19316_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .I1(net1363),
    .S(_05614_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19317_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .I1(net1349),
    .S(_05614_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19318_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .I1(net1348),
    .S(_05614_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19319_ (.A1(_04691_),
    .A2(_05578_),
    .Z(_05619_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1593 (.I(_09881_),
    .Z(net1592));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19321_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S(_05619_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19322_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .S(_05619_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19323_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .S(net1489),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19324_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .S(_05619_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19325_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .S(net1486),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19326_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .S(_05619_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19327_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S(_05619_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19328_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S(_05619_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19329_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S(net1486),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19330_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .S(net1486),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19331_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S(_05619_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1592 (.I(_09884_),
    .Z(net1591));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19333_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S(_05619_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19334_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(_05619_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19335_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .S(net1489),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19336_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .S(_05619_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19337_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .S(net1486),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19338_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .S(_05619_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19339_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .S(net1486),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19340_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .S(net1486),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19341_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .S(_05619_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19342_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .S(net1486),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19343_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .S(net1486),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1594 (.I(_09875_),
    .Z(net1593));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19345_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .S(net1486),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19346_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .S(_05619_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19347_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .S(net1489),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19348_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .S(_05619_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19349_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .S(net1486),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19350_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .S(_05619_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19351_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .S(net1486),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19352_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .S(net1486),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19353_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .S(net1486),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19354_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .S(net1486),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19355_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .S(net1486),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19356_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .S(net1486),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19357_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .S(net1486),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19358_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .S(net1489),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19359_ (.A1(_04691_),
    .A2(_05045_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1597 (.I(_09838_),
    .Z(net1596));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19361_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(_05623_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19362_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S(_05623_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19363_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S(_05623_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19364_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S(net1485),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19365_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(_05623_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19366_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(_05623_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19367_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S(_05623_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19368_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(net1485),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19369_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(net1485),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19370_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(_05623_),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19371_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .S(net1489),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1596 (.I(_09857_),
    .Z(net1595));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19373_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(_05623_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19374_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(_05623_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19375_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S(_05623_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19376_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(net1485),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19377_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S(_05623_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19378_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(net1485),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19379_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S(net1485),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19380_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S(_05623_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19381_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S(net1485),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19382_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S(net1485),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19383_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .S(net1489),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1599 (.I(_09824_),
    .Z(net1598));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19385_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S(net1485),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19386_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S(_05623_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19387_ (.I0(net1359),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S(_05623_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19388_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S(net1485),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19389_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S(_05623_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19390_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S(net1485),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19391_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(net1485),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19392_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S(net1485),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19393_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S(net1485),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19394_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S(net1485),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19395_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .S(net1489),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19396_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S(net1485),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19397_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S(net1485),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19398_ (.A1(_07968_),
    .A2(_09519_),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_04695_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19399_ (.A1(_09518_),
    .A2(_05627_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1595 (.I(_09872_),
    .Z(net1594));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19401_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .S(_05628_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19402_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .S(_05628_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19403_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .S(_05628_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19404_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .S(net1484),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19405_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .S(_05628_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19406_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .S(_05628_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19407_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .S(_05628_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19408_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .S(net1484),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19409_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .S(net1489),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19410_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .S(net1484),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19411_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .S(_05628_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1591 (.I(_09893_),
    .Z(net1590));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19413_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .S(_05628_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19414_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .S(_05628_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19415_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .S(_05628_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19416_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .S(net1484),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19417_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .S(_05628_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19418_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .S(net1484),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19419_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .S(net1484),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19420_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .S(_05628_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload43 (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19422_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .S(net1489),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19423_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .S(net1484),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19424_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .S(net1484),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload46 (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19426_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .S(net1484),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19427_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .S(_05628_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19428_ (.I0(net2471),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .S(net1484),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19429_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .S(net1484),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19430_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .S(net1484),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19431_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .S(net1484),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19432_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .S(net1484),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19433_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .S(net1484),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19434_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .S(net1489),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19435_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .S(net1484),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19436_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .S(net1484),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19437_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .S(net1484),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19438_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .S(net1484),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19439_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A2(_09519_),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_04695_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19440_ (.A1(_09518_),
    .A2(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2084 (.I(_00869_),
    .Z(net2083));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19442_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .I1(net1379),
    .S(_05634_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19443_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .I1(net1453),
    .S(_05634_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19444_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .I1(_05543_),
    .S(_05634_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19445_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .I1(_05565_),
    .S(net1482),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19446_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .I1(_05042_),
    .S(net1483),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19447_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .I1(net1396),
    .S(net1483),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19448_ (.I0(net2473),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .S(net1489),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19449_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .I1(net1399),
    .S(_05634_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19450_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .I1(_05450_),
    .S(_05634_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1509 (.I(_04551_),
    .Z(net1508));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19452_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .I1(net1392),
    .S(_05634_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 clone2090 (.I(net2091),
    .Z(net2089));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19454_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .I1(net1388),
    .S(net1483),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1486 (.I(_05623_),
    .Z(net1485));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1485 (.I(_05628_),
    .Z(net1484));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19457_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .I1(net1381),
    .S(net1483),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1483 (.I(_05634_),
    .Z(net1482));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19459_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .I1(net1376),
    .S(_05634_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1478 (.I(_05679_),
    .Z(net1477));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19461_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .I1(net1375),
    .S(net1483),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1476 (.I(_05681_),
    .Z(net1475));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19463_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .I1(net1377),
    .S(net1482),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1474 (.I(_05689_),
    .Z(net1473));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19465_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .I1(net1371),
    .S(net1483),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1471 (.I(_05698_),
    .Z(net1470));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19467_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .I1(net1374),
    .S(net1482),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19468_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .S(net1489),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1470 (.I(_05702_),
    .Z(net1469));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19470_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .I1(net1370),
    .S(net1482),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1468 (.I(_05706_),
    .Z(net1467));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19472_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .I1(net1362),
    .S(net1483),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1466 (.I(_05711_),
    .Z(net1465));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19474_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .I1(net1368),
    .S(net1482),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 rebuffer2476 (.I(net2481),
    .Z(net2475));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19476_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .I1(net1366),
    .S(_05634_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output255 (.I(net254),
    .Z(instr_req_o));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output254 (.I(net253),
    .Z(instr_addr_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19479_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .I1(net1354),
    .S(_05634_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output253 (.I(net252),
    .Z(instr_addr_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19481_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .I1(net1360),
    .S(net1483),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output252 (.I(net251),
    .Z(instr_addr_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19483_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .I1(net2472),
    .S(net1482),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output251 (.I(net250),
    .Z(instr_addr_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19485_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .I1(net1353),
    .S(net1482),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output250 (.I(net249),
    .Z(instr_addr_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19487_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .I1(net1352),
    .S(net1483),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output249 (.I(net248),
    .Z(instr_addr_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19489_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .I1(net1356),
    .S(net1482),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19490_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .S(net1489),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output248 (.I(net247),
    .Z(instr_addr_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19492_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .I1(net1351),
    .S(_05634_),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output247 (.I(net246),
    .Z(instr_addr_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19494_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .I1(net1364),
    .S(net1482),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output246 (.I(net245),
    .Z(instr_addr_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19496_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .I1(net1350),
    .S(_05634_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output245 (.I(net244),
    .Z(instr_addr_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19498_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .I1(net1363),
    .S(net1482),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output244 (.I(net243),
    .Z(instr_addr_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19500_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .I1(net1349),
    .S(net1482),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output243 (.I(net242),
    .Z(instr_addr_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19502_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .I1(net1348),
    .S(_05634_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output242 (.I(net241),
    .Z(instr_addr_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _19504_ (.A1(_07968_),
    .A2(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A3(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A4(_04695_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19505_ (.A1(_09518_),
    .A2(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output241 (.I(net240),
    .Z(instr_addr_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19507_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .I1(net1379),
    .S(_05664_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output240 (.I(net239),
    .Z(instr_addr_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19509_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .I1(net1453),
    .S(_05664_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output239 (.I(net238),
    .Z(instr_addr_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19511_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .I1(_05543_),
    .S(_05664_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output238 (.I(net237),
    .Z(instr_addr_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19513_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .I1(_05565_),
    .S(net1481),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19514_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .S(net1489),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output237 (.I(net236),
    .Z(instr_addr_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19516_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .I1(_05042_),
    .S(net1480),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output236 (.I(net235),
    .Z(instr_addr_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19518_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .I1(net1396),
    .S(net1480),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output235 (.I(net234),
    .Z(instr_addr_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19520_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .I1(net1399),
    .S(_05664_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output234 (.I(net233),
    .Z(instr_addr_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19522_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .I1(_05450_),
    .S(_05664_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19523_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .I1(net1392),
    .S(_05664_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19524_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .I1(net1388),
    .S(net1480),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output233 (.I(net232),
    .Z(instr_addr_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19526_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .I1(net1381),
    .S(net1480),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19527_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .I1(net1376),
    .S(_05664_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19528_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .I1(net1375),
    .S(net1480),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19529_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .I1(net1377),
    .S(net1481),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19530_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .S(net1489),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19531_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .I1(net1371),
    .S(net1480),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19532_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .I1(net1374),
    .S(net1481),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19533_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .I1(net1370),
    .S(net1481),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19534_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .I1(net1362),
    .S(net1480),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19535_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .I1(net1368),
    .S(net1481),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19536_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .I1(net1366),
    .S(_05664_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output232 (.I(net231),
    .Z(instr_addr_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19538_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .I1(net1354),
    .S(_05664_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19539_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .I1(net1360),
    .S(net1481),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19540_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .I1(net2471),
    .S(net1481),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19541_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .I1(net1353),
    .S(net1481),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19542_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .S(net1489),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19543_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .I1(net1352),
    .S(net1480),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19544_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .I1(net1356),
    .S(net1481),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19545_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .I1(net1351),
    .S(_05664_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19546_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .I1(net1364),
    .S(net1481),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19547_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .I1(net1350),
    .S(_05664_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19548_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .I1(net1363),
    .S(net1481),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19549_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .I1(net1349),
    .S(net1481),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19550_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .I1(net1348),
    .S(_05664_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19551_ (.A1(_09518_),
    .A2(_04696_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output231 (.I(net230),
    .Z(instr_addr_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19553_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .I1(net1379),
    .S(_05675_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19554_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .I1(net1453),
    .S(_05675_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19555_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .S(net1489),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19556_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .I1(_05543_),
    .S(_05675_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19557_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .I1(_05565_),
    .S(net1479),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19558_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .I1(_05042_),
    .S(net1478),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19559_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .I1(net1396),
    .S(net1478),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19560_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .I1(net1399),
    .S(_05675_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19561_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .I1(_05450_),
    .S(_05675_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19562_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .I1(net1392),
    .S(_05675_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19563_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .I1(net1388),
    .S(net1478),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output230 (.I(net229),
    .Z(instr_addr_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19565_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .I1(net1381),
    .S(net1478),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19566_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .I1(net1376),
    .S(_05675_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19567_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .S(net1489),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19568_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .I1(net1375),
    .S(net1478),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19569_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .I1(net1377),
    .S(net1479),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19570_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .I1(net1371),
    .S(net1478),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19571_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .I1(net1374),
    .S(net1479),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19572_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .I1(net1370),
    .S(net1479),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19573_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .I1(net1362),
    .S(net1478),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19574_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .I1(net1368),
    .S(net1479),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19575_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .I1(net1366),
    .S(_05675_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output229 (.I(net228),
    .Z(instr_addr_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19577_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .I1(net1354),
    .S(_05675_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19578_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .I1(net1360),
    .S(net1478),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19579_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .S(net1489),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19580_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .I1(net2471),
    .S(net1479),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19581_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .I1(net1353),
    .S(net1479),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19582_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .I1(net1352),
    .S(net1478),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19583_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .I1(net1356),
    .S(net1479),
    .Z(_02470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19584_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .I1(net1351),
    .S(_05675_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19585_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .I1(net1364),
    .S(net1479),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19586_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .I1(net1350),
    .S(_05675_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19587_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .I1(net1363),
    .S(net1479),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19588_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .I1(net1349),
    .S(net1479),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19589_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .I1(net1348),
    .S(net1478),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19590_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .S(net1489),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19591_ (.A1(_05500_),
    .A2(_05627_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output228 (.I(net227),
    .Z(instr_addr_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19593_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .S(_05679_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19594_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .S(_05679_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19595_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .S(_05679_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19596_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .S(net1477),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19597_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .S(_05679_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19598_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .S(net1477),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19599_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .S(_05679_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19600_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .S(net1477),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19601_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .S(net1477),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19602_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .S(_05679_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19603_ (.A1(_09518_),
    .A2(_05578_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output227 (.I(net226),
    .Z(instr_addr_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19605_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .I1(net1379),
    .S(_05681_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output226 (.I(net225),
    .Z(instr_addr_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19607_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .S(_05679_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19608_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .S(_05679_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19609_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .S(_05679_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19610_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .S(net1477),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19611_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .S(_05679_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19612_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .S(_05679_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19613_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .S(net1477),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19614_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .S(_05679_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19615_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .S(net1477),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19616_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .S(net1477),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19617_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .I1(net1453),
    .S(_05681_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output225 (.I(net224),
    .Z(instr_addr_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19619_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .S(net1477),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19620_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .S(_05679_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19621_ (.I0(net2472),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .S(net1477),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19622_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .S(net1477),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19623_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .S(_05679_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19624_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .S(net1477),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19625_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .S(net1477),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19626_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .S(net1477),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19627_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .S(net1477),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19628_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .S(net1477),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19629_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .I1(_05543_),
    .S(_05681_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19630_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .S(net1477),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19631_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .S(net1477),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19632_ (.A1(_05500_),
    .A2(_05633_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output224 (.I(net223),
    .Z(data_we_o));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19634_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .I1(net1379),
    .S(_05685_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19635_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .I1(net1453),
    .S(_05685_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19636_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .I1(_05543_),
    .S(_05685_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19637_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .I1(_05565_),
    .S(net1474),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19638_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .I1(_05042_),
    .S(_05685_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19639_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .I1(net1396),
    .S(net1474),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19640_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .I1(net1399),
    .S(_05685_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19641_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .I1(_05450_),
    .S(net1474),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19642_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .I1(_05565_),
    .S(net1475),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19643_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .I1(net1392),
    .S(net1474),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19644_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .I1(net1388),
    .S(_05685_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output223 (.I(net222),
    .Z(data_wdata_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19646_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .I1(net1381),
    .S(_05685_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19647_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .I1(net1376),
    .S(_05685_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19648_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .I1(net1375),
    .S(_05685_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19649_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .I1(net1377),
    .S(net1474),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19650_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .I1(net1371),
    .S(_05685_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19651_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .I1(net1374),
    .S(_05685_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19652_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .I1(net1370),
    .S(net1474),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19653_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .I1(net1362),
    .S(_05685_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19654_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .I1(_05042_),
    .S(_05681_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19655_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .I1(net1368),
    .S(net1474),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19656_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .I1(net1366),
    .S(net1474),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output222 (.I(net221),
    .Z(data_wdata_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19658_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .I1(net1354),
    .S(net1474),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19659_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .I1(net1360),
    .S(_05685_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19660_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .I1(net2471),
    .S(net1474),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19661_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .I1(net1353),
    .S(net1474),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19662_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .I1(net1352),
    .S(_05685_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19663_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .I1(net1356),
    .S(net1474),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19664_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .I1(net1351),
    .S(net1474),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19665_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .I1(net1364),
    .S(net1474),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19666_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .I1(net1396),
    .S(_05681_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19667_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .I1(net2470),
    .S(net1474),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19668_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .I1(net1363),
    .S(net1474),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19669_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .I1(net1349),
    .S(net1474),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19670_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .I1(net1348),
    .S(net1474),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19671_ (.A1(_05500_),
    .A2(_05663_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output221 (.I(net220),
    .Z(data_wdata_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19673_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .I1(net1379),
    .S(net1473),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19674_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .I1(net1453),
    .S(net1473),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19675_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .I1(_05543_),
    .S(net1473),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19676_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .I1(_05565_),
    .S(net1473),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19677_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .I1(_05042_),
    .S(net1473),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19678_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .I1(net1396),
    .S(net1473),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19679_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .I1(net1399),
    .S(_05681_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19680_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .I1(net1399),
    .S(net1473),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19681_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .I1(_05450_),
    .S(net1473),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19682_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .I1(net1392),
    .S(net1473),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19683_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .I1(net1388),
    .S(net1473),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output220 (.I(net219),
    .Z(data_wdata_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19685_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .I1(net1381),
    .S(net1473),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19686_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .I1(net1376),
    .S(net1473),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19687_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .I1(net1375),
    .S(net1473),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19688_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .I1(net1377),
    .S(net1473),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19689_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .I1(net1371),
    .S(net1473),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19690_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .I1(net1374),
    .S(net1473),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19691_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .I1(_05450_),
    .S(_05681_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19692_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .I1(net1370),
    .S(net1473),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19693_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .I1(net1362),
    .S(net1473),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19694_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .I1(net1368),
    .S(net1473),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19695_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .I1(net1366),
    .S(net1473),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net218),
    .Z(data_wdata_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19697_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .I1(net1354),
    .S(net1473),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19698_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .I1(net1360),
    .S(net1473),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19699_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .I1(net2471),
    .S(net1473),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19700_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .I1(net1353),
    .S(net1473),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19701_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .I1(net1352),
    .S(net1473),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19702_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .I1(net1356),
    .S(net1473),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19703_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .I1(net1392),
    .S(net1475),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19704_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .I1(net1351),
    .S(net1473),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19705_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .I1(net1364),
    .S(net1473),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19706_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .I1(net2494),
    .S(net1473),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19707_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .I1(net1363),
    .S(net1473),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19708_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .I1(net1349),
    .S(net1473),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19709_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .I1(net1348),
    .S(net1473),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19710_ (.A1(_04696_),
    .A2(_05500_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net217),
    .Z(data_wdata_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19712_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(_05693_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19713_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(_05693_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19714_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S(_05693_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19715_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S(net1472),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19716_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .I1(net1388),
    .S(net1475),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19717_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S(_05693_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19718_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S(net1472),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19719_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S(_05693_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19720_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S(net1472),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19721_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(net1472),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19722_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S(_05693_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net216),
    .Z(data_wdata_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19724_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S(_05693_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19725_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(_05693_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19726_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S(_05693_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19727_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S(net1472),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net215),
    .Z(data_wdata_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19729_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .I1(net1381),
    .S(net1475),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19730_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(net1472),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19731_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S(net1472),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19732_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(net1472),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19733_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S(_05693_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19734_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S(net1472),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19735_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S(net1472),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net214),
    .Z(data_wdata_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19737_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S(net1472),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19738_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S(net1472),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19739_ (.I0(net2472),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S(net1472),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19740_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S(net1472),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19741_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .I1(net1376),
    .S(_05681_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19742_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S(net1472),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19743_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S(net1472),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19744_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S(net1472),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19745_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S(net1472),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19746_ (.I0(net2470),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S(net1472),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19747_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(net1472),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19748_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S(net1472),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19749_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S(net1472),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19750_ (.A1(_05591_),
    .A2(_05627_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net213),
    .Z(data_wdata_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19752_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .I1(net1379),
    .S(net1470),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19753_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .I1(net1453),
    .S(net1470),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19754_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .I1(net1375),
    .S(net1475),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19755_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .I1(_05543_),
    .S(net1470),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19756_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .I1(_05565_),
    .S(net1471),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19757_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .I1(_05042_),
    .S(net1470),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19758_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .I1(net1396),
    .S(net1471),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19759_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .I1(net1399),
    .S(net1470),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19760_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .I1(_05450_),
    .S(net1471),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19761_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .I1(net1392),
    .S(net1471),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19762_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .I1(net1388),
    .S(net1470),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net212),
    .Z(data_wdata_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19764_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .I1(net1381),
    .S(net1471),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19765_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .I1(net1376),
    .S(net1470),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19766_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .I1(net1377),
    .S(net1475),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19767_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .I1(net1375),
    .S(net1470),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19768_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .I1(net1377),
    .S(net1471),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19769_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .I1(net1371),
    .S(net1470),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19770_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .I1(net1374),
    .S(net1471),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19771_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .I1(net1370),
    .S(net1471),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19772_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .I1(net1362),
    .S(net1470),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19773_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .I1(net1368),
    .S(net1471),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19774_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .I1(net1366),
    .S(net1471),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net211),
    .Z(data_wdata_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19776_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .I1(net1354),
    .S(net1471),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19777_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .I1(net1360),
    .S(net1470),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19778_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .I1(net1371),
    .S(net1475),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19779_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .I1(net2473),
    .S(net1471),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19780_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .I1(net1353),
    .S(net1471),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19781_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .I1(net1352),
    .S(net1470),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19782_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .I1(net1356),
    .S(net1471),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19783_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .I1(net1351),
    .S(net1471),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19784_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .I1(net1364),
    .S(net1471),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19785_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .I1(net1350),
    .S(net1471),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19786_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .I1(net1363),
    .S(net1471),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19787_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .I1(net1349),
    .S(net1471),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19788_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .I1(net1348),
    .S(net1471),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19789_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .I1(net1374),
    .S(net1475),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19790_ (.A1(_05591_),
    .A2(_05633_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net210),
    .Z(data_wdata_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19792_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .S(net1469),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19793_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .S(net1469),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19794_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .S(net1469),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19795_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .S(net1469),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19796_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .S(net1469),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19797_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .S(net1469),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19798_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .S(net1469),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19799_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .S(_05702_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19800_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .S(_05702_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19801_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .S(net1469),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19802_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .I1(net1370),
    .S(net1476),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net209),
    .Z(data_wdata_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19804_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .S(net1469),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19805_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .S(net1469),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19806_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .S(net1469),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19807_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .S(net1469),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19808_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .S(net1469),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19809_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .S(net1469),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19810_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .S(net1469),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19811_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .S(net1469),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19812_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .S(net1469),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19813_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .S(_05702_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19814_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .I1(net1362),
    .S(net1475),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net208),
    .Z(data_wdata_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19816_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .S(_05702_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19817_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .S(net1469),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19818_ (.I0(net1359),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .S(net1469),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19819_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .S(net1469),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19820_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .S(net1469),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19821_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .S(net1469),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19822_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .S(_05702_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19823_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .S(net1469),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19824_ (.I0(net2494),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .S(_05702_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19825_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .S(net1469),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19826_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .I1(net1368),
    .S(net1476),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19827_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .S(net1469),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19828_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .S(net1469),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19829_ (.A1(_05591_),
    .A2(_05663_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net207),
    .Z(data_wdata_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19831_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .I1(net1379),
    .S(net1467),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19832_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .I1(net1453),
    .S(net1467),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19833_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .I1(_05543_),
    .S(net1467),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19834_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .I1(_05565_),
    .S(net1468),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19835_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .I1(_05042_),
    .S(net1467),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19836_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .I1(net1396),
    .S(net1468),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19837_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .I1(net1399),
    .S(net1467),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19838_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .I1(_05450_),
    .S(net1468),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19839_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .I1(net1366),
    .S(net1476),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19840_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .I1(net1392),
    .S(net1468),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19841_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .I1(net1388),
    .S(net1467),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net206),
    .Z(data_wdata_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19843_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .I1(net1381),
    .S(net1468),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19844_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .I1(net1376),
    .S(net1467),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19845_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .I1(net1375),
    .S(net1467),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19846_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .I1(net1377),
    .S(net1468),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19847_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .I1(net1371),
    .S(net1467),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19848_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .I1(net1374),
    .S(net1467),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19849_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .I1(net1370),
    .S(net1468),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19850_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .I1(net1362),
    .S(net1467),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net205),
    .Z(data_wdata_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19852_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .I1(net1354),
    .S(net1476),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19853_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .I1(net1368),
    .S(net1468),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19854_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .I1(net1366),
    .S(net1468),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net204),
    .Z(data_wdata_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19856_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .I1(net1354),
    .S(net1468),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19857_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .I1(net1360),
    .S(net1467),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19858_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .I1(net1359),
    .S(net1468),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19859_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .I1(net1353),
    .S(net1468),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19860_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .I1(net1352),
    .S(net1467),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19861_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .I1(net1356),
    .S(net1468),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19862_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .I1(net1351),
    .S(net1468),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19863_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .I1(net1364),
    .S(net1468),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19864_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .I1(net1360),
    .S(net1475),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19865_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .I1(net2494),
    .S(net1468),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19866_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .I1(net1363),
    .S(net1468),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19867_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .I1(net1349),
    .S(net1468),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19868_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .I1(net1348),
    .S(net1468),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19869_ (.A1(_04696_),
    .A2(_05591_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net203),
    .Z(data_wdata_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19871_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .I1(net1379),
    .S(net1465),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19872_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .I1(net1453),
    .S(net1465),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19873_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .I1(_05543_),
    .S(net1465),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19874_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .I1(_05565_),
    .S(net1466),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19875_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .I1(_05042_),
    .S(net1465),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19876_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .I1(net1396),
    .S(net1466),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19877_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .I1(net2472),
    .S(net1475),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19878_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .I1(net1399),
    .S(net1465),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19879_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .I1(_05450_),
    .S(_05711_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19880_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .I1(net1392),
    .S(_05711_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19881_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .I1(net1388),
    .S(net1465),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net202),
    .Z(data_wdata_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19883_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .I1(net1381),
    .S(net1466),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19884_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .I1(net1376),
    .S(net1465),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19885_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .I1(net1375),
    .S(net1465),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19886_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .I1(net1377),
    .S(net1466),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19887_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .I1(net1371),
    .S(net1465),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19888_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .I1(net1374),
    .S(net1466),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19889_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .I1(net1353),
    .S(net1476),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19890_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .I1(net1370),
    .S(net1466),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19891_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .I1(net1362),
    .S(net1465),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19892_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .I1(net1368),
    .S(net1466),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19893_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .I1(net1366),
    .S(_05711_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net201),
    .Z(data_wdata_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19895_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .I1(net1354),
    .S(_05711_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19896_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .I1(net1360),
    .S(net1465),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19897_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .I1(net1359),
    .S(net1466),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19898_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .I1(net1353),
    .S(net1466),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19899_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .I1(net1352),
    .S(net1465),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19900_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .I1(net1356),
    .S(net1466),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19901_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .I1(net1352),
    .S(net1475),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19902_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .I1(net1351),
    .S(_05711_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19903_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .I1(net1364),
    .S(net1466),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19904_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .I1(net1350),
    .S(_05711_),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19905_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .I1(net1363),
    .S(net1466),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19906_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .I1(net1349),
    .S(net1466),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19907_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .I1(net1348),
    .S(_05711_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19908_ (.A1(_04691_),
    .A2(_05627_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net200),
    .Z(data_wdata_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19910_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .I1(net1379),
    .S(net1463),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19911_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .I1(net1453),
    .S(net1463),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19912_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .I1(_05543_),
    .S(net1463),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19913_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .I1(_05565_),
    .S(net1464),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19914_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .I1(net1356),
    .S(net1476),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19915_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .I1(_05042_),
    .S(net1463),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19916_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .I1(net1396),
    .S(net1464),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19917_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .I1(net1399),
    .S(net1463),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19918_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .I1(_05450_),
    .S(net1464),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19919_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .I1(net1392),
    .S(net1464),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19920_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .I1(net1388),
    .S(net1463),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net199),
    .Z(data_wdata_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19922_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .I1(net1381),
    .S(net1464),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19923_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .I1(net1376),
    .S(net1463),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19924_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .I1(net1375),
    .S(net1463),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19925_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .I1(net1377),
    .S(net1464),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19926_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .I1(net1351),
    .S(net1476),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19927_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .I1(net1371),
    .S(net1463),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19928_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .I1(net1374),
    .S(net1464),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19929_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .I1(net1370),
    .S(net1464),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19930_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .I1(net1362),
    .S(net1463),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19931_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .I1(net1368),
    .S(net1464),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19932_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .I1(net1366),
    .S(net1464),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net198),
    .Z(data_wdata_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19934_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .I1(net1354),
    .S(net1464),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19935_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .I1(net1360),
    .S(net1463),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19936_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .I1(net1359),
    .S(net1464),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19937_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .I1(net1353),
    .S(net1464),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19938_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .I1(net1364),
    .S(net1476),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19939_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .I1(net1352),
    .S(net1463),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19940_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .I1(net1356),
    .S(net1464),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19941_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .I1(net1351),
    .S(net1464),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19942_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .I1(net1364),
    .S(net1464),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19943_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .I1(net1350),
    .S(net1464),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19944_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .I1(net1363),
    .S(net1464),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19945_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .I1(net1349),
    .S(net1464),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19946_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .I1(net1348),
    .S(net1464),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _19947_ (.A1(_04691_),
    .A2(_05633_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net197),
    .Z(data_wdata_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19949_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .I1(net1379),
    .S(_05719_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19950_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .I1(net1453),
    .S(_05719_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19951_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .I1(net2470),
    .S(net1476),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19952_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .I1(_05543_),
    .S(net1461),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19953_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .I1(_05565_),
    .S(net1461),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19954_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .I1(_05042_),
    .S(_05719_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19955_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .I1(net1396),
    .S(net1461),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19956_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .I1(net1399),
    .S(_05719_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19957_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .I1(_05450_),
    .S(net1462),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19958_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .I1(net1392),
    .S(net1462),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19959_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .I1(net1388),
    .S(net1461),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net196),
    .Z(data_wdata_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19961_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .I1(net1381),
    .S(net1461),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19962_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .I1(net1376),
    .S(_05719_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19963_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .I1(net1363),
    .S(net1476),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19964_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .I1(net1375),
    .S(net1461),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19965_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .I1(net1377),
    .S(net1462),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19966_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .I1(net1371),
    .S(net1461),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19967_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .I1(net1374),
    .S(net1461),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19968_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .I1(net1370),
    .S(net1462),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19969_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .I1(net1362),
    .S(net1461),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19970_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .I1(net1368),
    .S(net1462),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19971_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .I1(net1366),
    .S(net1462),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net195),
    .Z(data_wdata_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19973_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .I1(net1354),
    .S(net1462),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19974_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .I1(net1360),
    .S(net1461),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19975_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .I1(net1349),
    .S(net1476),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19976_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .I1(net2471),
    .S(net1461),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19977_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .I1(net1353),
    .S(net1462),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19978_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .I1(net1352),
    .S(net1461),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19979_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .I1(net1356),
    .S(net1461),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19980_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .I1(net1351),
    .S(net1462),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19981_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .I1(net1364),
    .S(net1461),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19982_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .I1(net2494),
    .S(net1462),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19983_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .I1(net1363),
    .S(net1462),
    .Z(_02826_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19984_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .I1(net1349),
    .S(net1462),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19985_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .I1(net1348),
    .S(_05719_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19986_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .I1(net1348),
    .S(_05681_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _19987_ (.A1(_04691_),
    .A2(_05663_),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net194),
    .Z(data_wdata_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19989_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S(_05723_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19990_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .S(_05723_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19991_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .S(_05723_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19992_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .S(net1460),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19993_ (.I0(_05042_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .S(_05723_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19994_ (.I0(net1396),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .S(net1460),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19995_ (.I0(net1399),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S(_05723_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19996_ (.I0(_05450_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .S(net1460),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19997_ (.I0(net1392),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .S(net1460),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19998_ (.I0(net1388),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S(_05723_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _19999_ (.I0(net1379),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net1496),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net193),
    .Z(data_wdata_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20001_ (.I0(net1381),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .S(net1460),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20002_ (.I0(net1376),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .S(_05723_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20003_ (.I0(net1375),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .S(_05723_),
    .Z(_02843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20004_ (.I0(net1377),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .S(net1460),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20005_ (.I0(net1371),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .S(_05723_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20006_ (.I0(net1374),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .S(_05723_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20007_ (.I0(net1370),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .S(net1460),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20008_ (.I0(net1362),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .S(_05723_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20009_ (.I0(net1368),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .S(net1460),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20010_ (.I0(net1366),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .S(net1460),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20011_ (.I0(net1453),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net1496),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net192),
    .Z(data_wdata_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20013_ (.I0(net1354),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .S(net1460),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20014_ (.I0(net1360),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .S(_05723_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20015_ (.I0(net1359),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .S(net1460),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20016_ (.I0(net1353),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .S(net1460),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20017_ (.I0(net1352),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .S(_05723_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20018_ (.I0(net1356),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .S(net1460),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20019_ (.I0(net1351),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .S(net1460),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20020_ (.I0(net1364),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .S(net1460),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20021_ (.I0(net1350),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .S(net1460),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20022_ (.I0(net1363),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .S(net1460),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20023_ (.I0(_05543_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net1496),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20024_ (.I0(net1349),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .S(net1460),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20025_ (.I0(net1348),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .S(net1460),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20026_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .I1(net1379),
    .S(_04697_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20027_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .I1(net1453),
    .S(_04697_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20028_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .I1(_05543_),
    .S(net1497),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20029_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .I1(_05565_),
    .S(net1498),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20030_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .I1(_05042_),
    .S(_04697_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20031_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .I1(net1396),
    .S(_04697_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20032_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .I1(net1399),
    .S(_04697_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20033_ (.I0(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .I1(_05450_),
    .S(_04697_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20034_ (.I0(_05565_),
    .I1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net1496),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20035_ (.A1(_09497_),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A3(_10074_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net191),
    .Z(data_wdata_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20037_ (.A1(net1932),
    .A2(_00948_),
    .A3(_09526_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20038_ (.I(_00948_),
    .ZN(_05730_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20039_ (.A1(net1903),
    .A2(_00952_),
    .A3(_05730_),
    .A4(_09638_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20040_ (.A1(_05729_),
    .A2(_05731_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20041_ (.A1(_07642_),
    .A2(_09533_),
    .A3(_09621_),
    .A4(_05732_),
    .Z(_05733_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20042_ (.A1(_09528_),
    .A2(_09898_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20043_ (.A1(_05734_),
    .A2(_09646_),
    .B(_09658_),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20044_ (.A1(_09625_),
    .A2(_05733_),
    .B(_05735_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20045_ (.A1(\id_stage_i.controller_i.exc_req_d ),
    .A2(_05736_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20046_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(\cs_registers_i.dcsr_q[2] ),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20047_ (.A1(_03900_),
    .A2(_05738_),
    .B(\cs_registers_i.debug_mode_i ),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20048_ (.I(_05739_),
    .ZN(_05740_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20049_ (.A1(net1395),
    .A2(_05740_),
    .ZN(_05741_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20050_ (.A1(_05727_),
    .A2(_05737_),
    .A3(_05741_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20051_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09942_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20052_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_09498_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20053_ (.A1(_09920_),
    .A2(_05744_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20054_ (.A1(_09919_),
    .A2(net1808),
    .A3(_05743_),
    .A4(_05745_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20055_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20056_ (.A1(_09617_),
    .A2(_05740_),
    .Z(_05748_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20057_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09920_),
    .A3(_05748_),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20058_ (.A1(_09497_),
    .A2(_05747_),
    .B(_05749_),
    .C(_09498_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20059_ (.A1(net1932),
    .A2(_09905_),
    .A3(_03995_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20060_ (.A1(_05740_),
    .A2(_05751_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20061_ (.A1(_09499_),
    .A2(_05752_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20062_ (.A1(_09528_),
    .A2(_09899_),
    .A3(_09902_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20063_ (.A1(_05753_),
    .A2(_05754_),
    .ZN(_05755_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20064_ (.A1(_03901_),
    .A2(_05746_),
    .A3(_05750_),
    .A4(_05755_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20065_ (.A1(_09942_),
    .A2(net1808),
    .A3(_09941_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20066_ (.A1(_03999_),
    .A2(_05736_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20067_ (.I(_05758_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _20068_ (.A1(_09624_),
    .A2(_09636_),
    .A3(_09616_),
    .A4(_05759_),
    .Z(_05760_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20069_ (.A1(_09624_),
    .A2(_09636_),
    .A3(_05759_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20070_ (.A1(_09559_),
    .A2(_09580_),
    .A3(_09583_),
    .ZN(_05762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20071_ (.A1(_09540_),
    .A2(_05758_),
    .B1(_05761_),
    .B2(_05762_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20072_ (.A1(_05760_),
    .A2(_05763_),
    .ZN(_05764_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20073_ (.A1(_05739_),
    .A2(_05757_),
    .B(_09617_),
    .C(_09618_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20074_ (.A1(_09497_),
    .A2(_09920_),
    .B(_05744_),
    .ZN(_05766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20075_ (.A1(_05765_),
    .A2(_05766_),
    .ZN(_05767_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20076_ (.I(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20077_ (.A1(_05727_),
    .A2(_05764_),
    .B(_05768_),
    .ZN(_05769_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20078_ (.A1(net1395),
    .A2(_05769_),
    .ZN(_05770_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20079_ (.A1(_09497_),
    .A2(_09618_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20080_ (.A1(_05748_),
    .A2(_05771_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20081_ (.A1(_05757_),
    .A2(_05770_),
    .A3(_05772_),
    .ZN(_05773_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20082_ (.A1(_05742_),
    .A2(_05756_),
    .B(_05773_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20083_ (.A1(_03436_),
    .A2(net1393),
    .A3(_05757_),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20084_ (.A1(net1395),
    .A2(_05740_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20085_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_05774_),
    .B(_05775_),
    .C(net1809),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20086_ (.A1(_05760_),
    .A2(_05763_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20087_ (.A1(_05757_),
    .A2(_05748_),
    .A3(_05771_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20088_ (.I(_05753_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20089_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09919_),
    .A3(net1808),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20090_ (.A1(_09920_),
    .A2(_05744_),
    .A3(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20091_ (.A1(_05779_),
    .A2(_05754_),
    .B(_05781_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20092_ (.A1(net1809),
    .A2(_05777_),
    .B(_05778_),
    .C(_05782_),
    .ZN(_05783_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20093_ (.A1(_05776_),
    .A2(_05783_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20094_ (.A1(_09910_),
    .A2(_05753_),
    .A3(_05754_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20095_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_09920_),
    .B1(_05740_),
    .B2(_05771_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20096_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_05785_),
    .Z(_05786_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20097_ (.A1(_05744_),
    .A2(_09921_),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20098_ (.A1(_05784_),
    .A2(_05786_),
    .A3(_05787_),
    .Z(_05788_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20099_ (.A1(_05737_),
    .A2(_05775_),
    .B(net1809),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20100_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .A2(_09919_),
    .A3(net1808),
    .A4(_05743_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20101_ (.A1(_09498_),
    .A2(_05790_),
    .B(_09921_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20102_ (.A1(_05788_),
    .A2(_05789_),
    .B(_05791_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20103_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_09910_),
    .A3(_05752_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20104_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_10074_),
    .A3(_05748_),
    .A4(_05792_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20105_ (.A1(_05727_),
    .A2(_05737_),
    .A3(_05775_),
    .B(_05793_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20106_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09919_),
    .B(_09922_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20107_ (.A1(_09942_),
    .A2(net1747),
    .B(_05794_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20108_ (.A1(net2038),
    .A2(_09938_),
    .A3(_09943_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20109_ (.A1(_09939_),
    .A2(_05795_),
    .B(net1746),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20110_ (.A1(_07575_),
    .A2(_09912_),
    .ZN(_05796_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20111_ (.A1(_08127_),
    .A2(_03422_),
    .A3(_03402_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20112_ (.A1(_05797_),
    .A2(_05484_),
    .B(_03404_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _20113_ (.A1(_05796_),
    .A2(_10125_),
    .A3(_03433_),
    .A4(_05798_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20114_ (.A1(_09538_),
    .A2(_09654_),
    .A3(_10125_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20115_ (.A1(_09621_),
    .A2(_03433_),
    .A3(_05800_),
    .B(\id_stage_i.id_fsm_q ),
    .ZN(_05801_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20116_ (.A1(_03403_),
    .A2(_05799_),
    .B(_05801_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net190),
    .Z(data_req_o));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20118_ (.I0(net1798),
    .I1(\alu_adder_result_ex[0] ),
    .S(net1672),
    .Z(_05803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20119_ (.I0(\ex_block_i.alu_i.imd_val_q_i[0] ),
    .I1(_05803_),
    .S(net1548),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20120_ (.I0(net1711),
    .I1(net1451),
    .S(net1672),
    .Z(_05804_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20121_ (.I0(\ex_block_i.alu_i.imd_val_q_i[10] ),
    .I1(_05804_),
    .S(net1548),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20122_ (.I0(net2158),
    .I1(net1457),
    .S(net1672),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20123_ (.I0(\ex_block_i.alu_i.imd_val_q_i[11] ),
    .I1(_05805_),
    .S(net1548),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20124_ (.I0(net2136),
    .I1(net2298),
    .S(net1672),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20125_ (.I0(\ex_block_i.alu_i.imd_val_q_i[12] ),
    .I1(_05806_),
    .S(net1548),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20126_ (.I0(net2157),
    .I1(net1450),
    .S(net1672),
    .Z(_05807_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20127_ (.I0(\ex_block_i.alu_i.imd_val_q_i[13] ),
    .I1(_05807_),
    .S(net1548),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20128_ (.I0(net2192),
    .I1(net2292),
    .S(net1672),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20129_ (.I0(\ex_block_i.alu_i.imd_val_q_i[14] ),
    .I1(_05808_),
    .S(net1548),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20130_ (.I0(net2187),
    .I1(net1448),
    .S(net1672),
    .Z(_05809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20131_ (.I0(\ex_block_i.alu_i.imd_val_q_i[15] ),
    .I1(_05809_),
    .S(net1548),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20132_ (.I0(net2190),
    .I1(net1446),
    .S(net1672),
    .Z(_05810_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20133_ (.I0(\ex_block_i.alu_i.imd_val_q_i[16] ),
    .I1(_05810_),
    .S(net1548),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20134_ (.I0(net1769),
    .I1(net2288),
    .S(net1672),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20135_ (.I0(\ex_block_i.alu_i.imd_val_q_i[17] ),
    .I1(_05811_),
    .S(net1548),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20136_ (.I0(net1768),
    .I1(net1435),
    .S(net1672),
    .Z(_05812_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net189),
    .Z(data_be_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20138_ (.I0(\ex_block_i.alu_i.imd_val_q_i[18] ),
    .I1(_05812_),
    .S(net1548),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net188),
    .Z(data_be_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20140_ (.I0(net1767),
    .I1(net1436),
    .S(net1672),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20141_ (.I0(\ex_block_i.alu_i.imd_val_q_i[19] ),
    .I1(_05815_),
    .S(net1548),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20142_ (.I0(net2185),
    .I1(net1539),
    .S(net1672),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20143_ (.I0(\ex_block_i.alu_i.imd_val_q_i[1] ),
    .I1(_05816_),
    .S(net1548),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20144_ (.I0(net1766),
    .I1(net2278),
    .S(net1672),
    .Z(_05817_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20145_ (.I0(\ex_block_i.alu_i.imd_val_q_i[20] ),
    .I1(_05817_),
    .S(net1548),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20146_ (.I0(net1763),
    .I1(net1410),
    .S(net1672),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20147_ (.I0(\ex_block_i.alu_i.imd_val_q_i[21] ),
    .I1(_05818_),
    .S(net1548),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20148_ (.I0(net1762),
    .I1(net1432),
    .S(net1672),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20149_ (.I0(\ex_block_i.alu_i.imd_val_q_i[22] ),
    .I1(_05819_),
    .S(net1548),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20150_ (.I0(net1761),
    .I1(net169),
    .S(net1672),
    .Z(_05820_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20151_ (.I0(\ex_block_i.alu_i.imd_val_q_i[23] ),
    .I1(_05820_),
    .S(net1548),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20152_ (.I0(net1760),
    .I1(net2204),
    .S(net1672),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20153_ (.I0(\ex_block_i.alu_i.imd_val_q_i[24] ),
    .I1(_05821_),
    .S(net1548),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20154_ (.I0(net1759),
    .I1(net1431),
    .S(net1672),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20155_ (.I0(\ex_block_i.alu_i.imd_val_q_i[25] ),
    .I1(_05822_),
    .S(net1548),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20156_ (.I0(net1758),
    .I1(net1409),
    .S(net1672),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20157_ (.I0(\ex_block_i.alu_i.imd_val_q_i[26] ),
    .I1(_05823_),
    .S(net1548),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20158_ (.I0(net1757),
    .I1(net1429),
    .S(net1672),
    .Z(_05824_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net187),
    .Z(data_be_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20160_ (.I0(\ex_block_i.alu_i.imd_val_q_i[27] ),
    .I1(_05824_),
    .S(net1548),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net186),
    .Z(data_be_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20162_ (.I0(net1756),
    .I1(net2138),
    .S(net1672),
    .Z(_05827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20163_ (.I0(\ex_block_i.alu_i.imd_val_q_i[28] ),
    .I1(_05827_),
    .S(net1548),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20164_ (.I0(net1755),
    .I1(net1408),
    .S(net1672),
    .Z(_05828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20165_ (.I0(\ex_block_i.alu_i.imd_val_q_i[29] ),
    .I1(_05828_),
    .S(net1548),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20166_ (.I0(net1740),
    .I1(net1521),
    .S(net1672),
    .Z(_05829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20167_ (.I0(\ex_block_i.alu_i.imd_val_q_i[2] ),
    .I1(_05829_),
    .S(net1548),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20168_ (.I0(net1753),
    .I1(net2122),
    .S(net1672),
    .Z(_05830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20169_ (.I0(\ex_block_i.alu_i.imd_val_q_i[30] ),
    .I1(_05830_),
    .S(net1548),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20170_ (.A1(net1783),
    .A2(_08174_),
    .A3(net2051),
    .Z(_05831_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20171_ (.A1(net1719),
    .A2(_05831_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20172_ (.I0(\ex_block_i.alu_i.imd_val_q_i[31] ),
    .I1(_05832_),
    .S(net1548),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net1459),
    .Z(data_addr_o[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net1458),
    .Z(data_addr_o[8]));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _20175_ (.A1(net2031),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A3(net1823),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net1512),
    .Z(data_addr_o[7]));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20177_ (.A1(net2019),
    .A2(net1825),
    .A3(_09677_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net1500),
    .Z(data_addr_o[6]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20179_ (.A1(net1806),
    .A2(net1613),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20180_ (.A1(net1718),
    .A2(_04683_),
    .ZN(_05840_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20181_ (.A1(net1784),
    .A2(net1718),
    .A3(_05839_),
    .B1(_05840_),
    .B2(_00972_),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20182_ (.A1(net1549),
    .A2(_04683_),
    .Z(_05842_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20183_ (.A1(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .A2(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20184_ (.I0(\ex_block_i.alu_i.imd_val_q_i[32] ),
    .I1(\alu_adder_result_ex[0] ),
    .S(net1398),
    .Z(_05844_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20185_ (.A1(_00964_),
    .A2(_04486_),
    .Z(_05845_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20186_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .A2(net1613),
    .A3(_05845_),
    .Z(_05846_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20187_ (.A1(net1673),
    .A2(_05844_),
    .B(_05846_),
    .C(net2029),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net1499),
    .Z(data_addr_o[5]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20189_ (.A1(net1750),
    .A2(net1549),
    .Z(_05849_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20190_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05850_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20191_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05851_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20192_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05852_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20193_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05853_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20194_ (.I0(_05850_),
    .I1(_05851_),
    .I2(_05852_),
    .I3(_05853_),
    .S0(_04401_),
    .S1(_04404_),
    .Z(_05854_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20195_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05855_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20196_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05856_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20197_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20198_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .I1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .I2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .I3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .S0(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(_00965_),
    .Z(_05858_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _20199_ (.I0(_05855_),
    .I1(_05856_),
    .I2(_05857_),
    .I3(_05858_),
    .S0(_04401_),
    .S1(_04404_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20200_ (.A1(_04498_),
    .A2(_04407_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20201_ (.I0(_05854_),
    .I1(_05859_),
    .S(_05860_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _20202_ (.A1(net2031),
    .A2(\alu_adder_result_ex[0] ),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C1(_05861_),
    .C2(net2027),
    .ZN(_05862_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20203_ (.A1(_09670_),
    .A2(_05847_),
    .A3(_05849_),
    .A4(_05862_),
    .Z(_05863_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20204_ (.A1(net1549),
    .A2(_05841_),
    .B(_05843_),
    .C(_05863_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20205_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .A2(_04514_),
    .Z(_05864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20206_ (.I0(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .I1(net1539),
    .S(net1398),
    .Z(_05865_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net1454),
    .Z(data_addr_o[4]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20208_ (.I0(_05864_),
    .I1(_05865_),
    .S(net1613),
    .Z(_05867_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20209_ (.A1(net1806),
    .A2(net1613),
    .Z(_05868_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net1519),
    .Z(data_addr_o[3]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20211_ (.A1(net2031),
    .A2(net1539),
    .B1(_05844_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20212_ (.A1(net1786),
    .A2(_05868_),
    .B(_05870_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20213_ (.A1(net2029),
    .A2(_05867_),
    .B(_05871_),
    .ZN(_05872_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net2051),
    .Z(data_addr_o[31]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20215_ (.A1(net1549),
    .A2(_04684_),
    .ZN(_05874_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20216_ (.A1(\ex_block_i.alu_i.imd_val_q_i[33] ),
    .A2(_05842_),
    .B1(_05874_),
    .B2(_00974_),
    .ZN(_05875_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20217_ (.A1(_05849_),
    .A2(_05872_),
    .B(_05875_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net2122),
    .Z(data_addr_o[30]));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20219_ (.A1(_00967_),
    .A2(_04486_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .ZN(_05877_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net1521),
    .Z(data_addr_o[2]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20221_ (.I0(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .I1(net1521),
    .S(net1398),
    .Z(_05879_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20222_ (.A1(net1673),
    .A2(_05879_),
    .B(net2029),
    .ZN(_05880_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net1408),
    .Z(data_addr_o[29]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20224_ (.A1(net2031),
    .A2(net1521),
    .B1(_05865_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05882_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20225_ (.A1(_05877_),
    .A2(_05880_),
    .B(_05882_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20226_ (.A1(net1781),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05884_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20227_ (.A1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A2(_05842_),
    .B(_05883_),
    .C(_05884_),
    .ZN(_05885_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20228_ (.A1(net1549),
    .A2(_04683_),
    .ZN(_05886_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net2138),
    .Z(data_addr_o[28]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20230_ (.A1(net1549),
    .A2(_04684_),
    .Z(_05888_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net1429),
    .Z(data_addr_o[27]));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20232_ (.A1(\ex_block_i.alu_i.imd_val_q_i[34] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_00975_),
    .ZN(_05890_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20233_ (.A1(_05885_),
    .A2(_05890_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20234_ (.I0(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .I1(net1519),
    .S(net1398),
    .Z(_05891_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20235_ (.A1(net1673),
    .A2(_05891_),
    .ZN(_05892_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20236_ (.A1(_00969_),
    .A2(_04486_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20237_ (.A1(net2031),
    .A2(net1519),
    .B1(_05879_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05894_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20238_ (.A1(_08196_),
    .A2(_05892_),
    .A3(_05893_),
    .B(_05894_),
    .ZN(_05895_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20239_ (.A1(net1780),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05896_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20240_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_05842_),
    .B(_05895_),
    .C(_05896_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20241_ (.A1(\ex_block_i.alu_i.imd_val_q_i[35] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_00980_),
    .ZN(_05898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20242_ (.A1(_05897_),
    .A2(_05898_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20243_ (.I0(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .I1(net1454),
    .S(net1398),
    .Z(_05899_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20244_ (.A1(_00964_),
    .A2(_04535_),
    .Z(_05900_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20245_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .A2(net1613),
    .A3(_05900_),
    .Z(_05901_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20246_ (.A1(net1673),
    .A2(_05899_),
    .B(_05901_),
    .C(net2029),
    .ZN(_05902_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20247_ (.A1(net2031),
    .A2(net1454),
    .B1(_05891_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20248_ (.A1(_05902_),
    .A2(_05903_),
    .Z(_05904_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20249_ (.A1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A2(_05842_),
    .B1(_05839_),
    .B2(net1715),
    .C(net1750),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20250_ (.A1(\ex_block_i.alu_i.imd_val_q_i[36] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_00981_),
    .ZN(_05906_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20251_ (.A1(_05904_),
    .A2(_05905_),
    .B(_05906_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20252_ (.I0(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .I1(net1499),
    .S(net1398),
    .Z(_05907_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20253_ (.A1(_00968_),
    .A2(_04535_),
    .Z(_05908_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20254_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .A2(net1613),
    .A3(_05908_),
    .Z(_05909_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20255_ (.A1(net1673),
    .A2(_05907_),
    .B(_05909_),
    .C(net2029),
    .ZN(_05910_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20256_ (.A1(net2031),
    .A2(net1499),
    .B1(_05899_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05911_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20257_ (.A1(_05910_),
    .A2(_05911_),
    .Z(_05912_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20258_ (.A1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A2(_05842_),
    .B1(_05839_),
    .B2(_04468_),
    .C(net1750),
    .ZN(_05913_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20259_ (.A1(\ex_block_i.alu_i.imd_val_q_i[37] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_00985_),
    .ZN(_05914_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20260_ (.A1(_05912_),
    .A2(_05913_),
    .B(_05914_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20261_ (.I0(net1749),
    .I1(net1519),
    .S(net1672),
    .Z(_05915_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20262_ (.I0(\ex_block_i.alu_i.imd_val_q_i[3] ),
    .I1(_05915_),
    .S(net1548),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20263_ (.I0(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .I1(net1500),
    .S(net1398),
    .Z(_05916_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20264_ (.A1(_00967_),
    .A2(_04535_),
    .Z(_05917_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20265_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .A2(net1613),
    .A3(_05917_),
    .Z(_05918_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20266_ (.A1(net1673),
    .A2(_05916_),
    .B(_05918_),
    .C(net2029),
    .ZN(_05919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20267_ (.A1(net2031),
    .A2(net1500),
    .B1(_05907_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05920_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20268_ (.A1(_05919_),
    .A2(_05920_),
    .Z(_05921_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20269_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_05842_),
    .B1(_05839_),
    .B2(_04471_),
    .C(net1750),
    .ZN(_05922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20270_ (.A1(\ex_block_i.alu_i.imd_val_q_i[38] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_00992_),
    .ZN(_05923_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20271_ (.A1(_05921_),
    .A2(_05922_),
    .B(_05923_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20272_ (.I0(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .I1(net1512),
    .S(net1398),
    .Z(_05924_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20273_ (.A1(_00969_),
    .A2(_04535_),
    .Z(_05925_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20274_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .A2(net1613),
    .A3(_05925_),
    .Z(_05926_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20275_ (.A1(net1673),
    .A2(_05924_),
    .B(_05926_),
    .C(net2029),
    .ZN(_05927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20276_ (.A1(net2031),
    .A2(net1512),
    .B1(_05916_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20277_ (.A1(_05927_),
    .A2(_05928_),
    .Z(_05929_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20278_ (.A1(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A2(_05842_),
    .B1(_05839_),
    .B2(_04474_),
    .C(net1750),
    .ZN(_05930_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20279_ (.A1(\ex_block_i.alu_i.imd_val_q_i[39] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_05437_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20280_ (.A1(_05929_),
    .A2(_05930_),
    .B(_05931_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20281_ (.A1(_04681_),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_04682_),
    .ZN(_05932_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20282_ (.I(net1549),
    .ZN(_05933_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20283_ (.A1(_00964_),
    .A2(_04493_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .ZN(_05934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20284_ (.I0(\ex_block_i.alu_i.imd_val_q_i[40] ),
    .I1(net1458),
    .S(net1398),
    .Z(_05935_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20285_ (.A1(net1673),
    .A2(_05935_),
    .ZN(_05936_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20286_ (.A1(net1673),
    .A2(_05934_),
    .B(_05936_),
    .C(_08196_),
    .ZN(_05937_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net1409),
    .Z(data_addr_o[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net1431),
    .Z(data_addr_o[25]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20289_ (.A1(net2031),
    .A2(net1458),
    .B1(_05924_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05940_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20290_ (.A1(net1775),
    .A2(_05868_),
    .B(_05940_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20291_ (.A1(net1718),
    .A2(_05933_),
    .A3(_05937_),
    .A4(_05941_),
    .Z(_05942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20292_ (.A1(_05932_),
    .A2(_05942_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20293_ (.A1(_09670_),
    .A2(_05849_),
    .ZN(_05943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20294_ (.A1(net2031),
    .A2(net1459),
    .B1(_05935_),
    .B2(net2027),
    .C(_05943_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20295_ (.I0(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .I1(net1459),
    .S(net1398),
    .Z(_05945_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20296_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .A2(net1613),
    .A3(_04543_),
    .Z(_05946_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20297_ (.A1(net1673),
    .A2(_05945_),
    .B(_05946_),
    .C(net2029),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20298_ (.A1(net2174),
    .A2(net1750),
    .ZN(_05948_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20299_ (.A1(_05840_),
    .A2(_04745_),
    .B1(_05839_),
    .B2(_05948_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20300_ (.A1(\ex_block_i.alu_i.imd_val_q_i[41] ),
    .A2(_05842_),
    .ZN(_05950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20301_ (.A1(_05944_),
    .A2(_05947_),
    .B1(_05949_),
    .B2(net1549),
    .C(_05950_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20302_ (.I0(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .I1(net1451),
    .S(net1398),
    .Z(_05951_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20303_ (.A1(net1673),
    .A2(_05951_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20304_ (.A1(_00967_),
    .A2(_04493_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20305_ (.A1(net2031),
    .A2(net1451),
    .B1(_05945_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05954_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20306_ (.A1(_08196_),
    .A2(_05952_),
    .A3(_05953_),
    .B(_05954_),
    .ZN(_05955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20307_ (.A1(net1735),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20308_ (.A1(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A2(_05842_),
    .B(_05955_),
    .C(_05956_),
    .ZN(_05957_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20309_ (.A1(\ex_block_i.alu_i.imd_val_q_i[42] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_04771_),
    .ZN(_05958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20310_ (.A1(_05957_),
    .A2(_05958_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20311_ (.I0(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .I1(net1457),
    .S(net1398),
    .Z(_05959_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20312_ (.A1(net1673),
    .A2(_05959_),
    .ZN(_05960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20313_ (.A1(_00969_),
    .A2(_04493_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .ZN(_05961_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20314_ (.A1(net2031),
    .A2(net1457),
    .B1(_05951_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05962_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20315_ (.A1(_08196_),
    .A2(_05960_),
    .A3(_05961_),
    .B(_05962_),
    .ZN(_05963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20316_ (.A1(net1738),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20317_ (.A1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .A2(_05842_),
    .B(_05963_),
    .C(_05964_),
    .ZN(_05965_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20318_ (.A1(\ex_block_i.alu_i.imd_val_q_i[43] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_04794_),
    .ZN(_05966_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20319_ (.A1(_05965_),
    .A2(_05966_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20320_ (.I0(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .I1(net2298),
    .S(net1398),
    .Z(_05967_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20321_ (.A1(net1673),
    .A2(_05967_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20322_ (.A1(_00964_),
    .A2(_04500_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .ZN(_05969_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20323_ (.A1(net2031),
    .A2(net2298),
    .B1(_05959_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05970_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20324_ (.A1(_08196_),
    .A2(_05968_),
    .A3(_05969_),
    .B(_05970_),
    .ZN(_05971_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20325_ (.A1(net1803),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20326_ (.A1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A2(_05842_),
    .B(_05971_),
    .C(_05972_),
    .ZN(_05973_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20327_ (.A1(\ex_block_i.alu_i.imd_val_q_i[44] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(net1391),
    .ZN(_05974_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20328_ (.A1(_05973_),
    .A2(_05974_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20329_ (.I0(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .I1(net1450),
    .S(net1398),
    .Z(_05975_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20330_ (.A1(net1673),
    .A2(_05975_),
    .ZN(_05976_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20331_ (.A1(_00968_),
    .A2(_04500_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .ZN(_05977_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20332_ (.A1(net2031),
    .A2(net1450),
    .B1(_05967_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05978_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20333_ (.A1(_08196_),
    .A2(_05976_),
    .A3(_05977_),
    .B(_05978_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20334_ (.A1(net1734),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05980_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20335_ (.A1(\ex_block_i.alu_i.imd_val_q_i[45] ),
    .A2(_05842_),
    .B(_05979_),
    .C(_05980_),
    .ZN(_05981_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20336_ (.A1(_04880_),
    .A2(_05842_),
    .B1(_05874_),
    .B2(_04885_),
    .C(_05981_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20337_ (.A1(_00967_),
    .A2(_04500_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20338_ (.I0(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .I1(net2292),
    .S(net1398),
    .Z(_05983_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20339_ (.A1(net1673),
    .A2(_05983_),
    .B(net2029),
    .ZN(_05984_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20340_ (.A1(net2031),
    .A2(net2292),
    .B1(_05975_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05985_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20341_ (.A1(_05982_),
    .A2(_05984_),
    .B(_05985_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20342_ (.A1(net1733),
    .A2(_05868_),
    .B(net1718),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20343_ (.A1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A2(_05842_),
    .B(_05986_),
    .C(_05987_),
    .ZN(_05988_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20344_ (.A1(\ex_block_i.alu_i.imd_val_q_i[46] ),
    .A2(_05886_),
    .B1(_05888_),
    .B2(_04926_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20345_ (.A1(_05988_),
    .A2(_05989_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20346_ (.I0(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .I1(net1448),
    .S(net1398),
    .Z(_05990_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20347_ (.A1(_00969_),
    .A2(_04500_),
    .Z(_05991_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20348_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .A2(net1613),
    .A3(_05991_),
    .Z(_05992_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20349_ (.A1(net1673),
    .A2(_05990_),
    .B(_05992_),
    .C(net2029),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20350_ (.A1(net2031),
    .A2(net1448),
    .B1(_05983_),
    .B2(net2027),
    .C(net1806),
    .ZN(_05994_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20351_ (.A1(_05993_),
    .A2(_05994_),
    .Z(_05995_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20352_ (.A1(\ex_block_i.alu_i.imd_val_q_i[47] ),
    .A2(_05842_),
    .B1(_05839_),
    .B2(net1748),
    .C(net1750),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _20353_ (.A1(_04952_),
    .A2(_05842_),
    .B1(_05995_),
    .B2(_05996_),
    .C1(_05874_),
    .C2(_04960_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20354_ (.I(net1794),
    .ZN(_05997_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20355_ (.I0(_05997_),
    .I1(net1454),
    .S(net1672),
    .Z(_05998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20356_ (.I0(\ex_block_i.alu_i.imd_val_q_i[4] ),
    .I1(_05998_),
    .S(net1548),
    .Z(_02923_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net2065),
    .Z(data_addr_o[24]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20358_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(net1446),
    .S(net1398),
    .Z(_06000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20359_ (.A1(_00964_),
    .A2(_04507_),
    .Z(_06001_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net169),
    .Z(data_addr_o[23]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20361_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .A2(net1613),
    .Z(_06003_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20362_ (.A1(net1673),
    .A2(_06000_),
    .B1(_06001_),
    .B2(_06003_),
    .C(net2029),
    .ZN(_06004_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net1432),
    .Z(data_addr_o[22]));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20364_ (.A1(net2031),
    .A2(net1446),
    .B1(_05990_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06006_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20365_ (.A1(net1770),
    .A2(_05868_),
    .B1(_06004_),
    .B2(_06006_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20366_ (.I0(_04978_),
    .I1(_06007_),
    .S(net1750),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20367_ (.I0(\ex_block_i.alu_i.imd_val_q_i[48] ),
    .I1(_06008_),
    .S(net1549),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20368_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(net2288),
    .S(net1398),
    .Z(_06009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20369_ (.A1(_00968_),
    .A2(_04507_),
    .Z(_06010_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20370_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(net1613),
    .Z(_06011_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20371_ (.A1(net1673),
    .A2(_06009_),
    .B1(_06010_),
    .B2(_06011_),
    .C(net2029),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20372_ (.A1(net2031),
    .A2(net2288),
    .B1(_06000_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20373_ (.A1(net1732),
    .A2(_05868_),
    .B1(_06012_),
    .B2(_06013_),
    .ZN(_06014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20374_ (.I0(_05004_),
    .I1(_06014_),
    .S(net1750),
    .Z(_06015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20375_ (.I0(\ex_block_i.alu_i.imd_val_q_i[49] ),
    .I1(_06015_),
    .S(net1549),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20376_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(net1435),
    .S(net1398),
    .Z(_06016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20377_ (.A1(_00967_),
    .A2(_04507_),
    .Z(_06017_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20378_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .A2(net1613),
    .Z(_06018_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20379_ (.A1(net1673),
    .A2(_06016_),
    .B1(_06017_),
    .B2(_06018_),
    .C(net2029),
    .ZN(_06019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20380_ (.A1(net2031),
    .A2(net1435),
    .B1(_06009_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20381_ (.A1(net1731),
    .A2(_05868_),
    .B1(_06019_),
    .B2(_06020_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20382_ (.I0(_05059_),
    .I1(_06021_),
    .S(net1750),
    .Z(_06022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20383_ (.I0(\ex_block_i.alu_i.imd_val_q_i[50] ),
    .I1(_06022_),
    .S(_09687_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20384_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(net1436),
    .S(net1398),
    .Z(_06023_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20385_ (.A1(_00969_),
    .A2(_04507_),
    .Z(_06024_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20386_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .A2(net1613),
    .Z(_06025_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20387_ (.A1(net1673),
    .A2(_06023_),
    .B1(_06024_),
    .B2(_06025_),
    .C(net2029),
    .ZN(_06026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20388_ (.A1(net2031),
    .A2(net1436),
    .B1(_06016_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06027_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20389_ (.A1(net1730),
    .A2(_05868_),
    .B1(_06026_),
    .B2(_06027_),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20390_ (.I0(_05082_),
    .I1(_06028_),
    .S(net1750),
    .Z(_06029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20391_ (.I0(\ex_block_i.alu_i.imd_val_q_i[51] ),
    .I1(_06029_),
    .S(_09687_),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20392_ (.A1(net1750),
    .A2(net1372),
    .ZN(_06030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20393_ (.I0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .I1(net2278),
    .S(net1398),
    .Z(_06031_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20394_ (.A1(_00964_),
    .A2(_04517_),
    .Z(_06032_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20395_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .A2(net1613),
    .Z(_06033_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20396_ (.A1(net1673),
    .A2(_06031_),
    .B1(_06032_),
    .B2(_06033_),
    .C(net2029),
    .ZN(_06034_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20397_ (.A1(net2031),
    .A2(net2278),
    .B1(_06023_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20398_ (.A1(net2161),
    .A2(_05868_),
    .B1(_06034_),
    .B2(_06035_),
    .C(net1718),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20399_ (.A1(_06030_),
    .A2(_06036_),
    .Z(_06037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20400_ (.I0(\ex_block_i.alu_i.imd_val_q_i[52] ),
    .I1(_06037_),
    .S(net1549),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20401_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(net1410),
    .S(net1398),
    .Z(_06038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20402_ (.A1(_00968_),
    .A2(_04517_),
    .Z(_06039_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20403_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .A2(net1613),
    .Z(_06040_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20404_ (.A1(net1673),
    .A2(_06038_),
    .B1(_06039_),
    .B2(_06040_),
    .C(net2029),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20405_ (.A1(net2031),
    .A2(net1410),
    .B1(_06031_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06042_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20406_ (.A1(net1727),
    .A2(_05868_),
    .B1(_06041_),
    .B2(_06042_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20407_ (.I0(_05127_),
    .I1(_06043_),
    .S(net1750),
    .Z(_06044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20408_ (.I0(\ex_block_i.alu_i.imd_val_q_i[53] ),
    .I1(_06044_),
    .S(_09687_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20409_ (.I0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .I1(net1432),
    .S(net1398),
    .Z(_06045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20410_ (.A1(_00967_),
    .A2(_04517_),
    .Z(_06046_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20411_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .A2(net1613),
    .Z(_06047_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20412_ (.A1(net1673),
    .A2(_06045_),
    .B1(_06046_),
    .B2(_06047_),
    .C(net2029),
    .ZN(_06048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20413_ (.A1(net2031),
    .A2(net1432),
    .B1(_06038_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20414_ (.A1(net1726),
    .A2(_05868_),
    .B1(_06048_),
    .B2(_06049_),
    .ZN(_06050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20415_ (.I0(_05147_),
    .I1(_06050_),
    .S(net1750),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20416_ (.I0(\ex_block_i.alu_i.imd_val_q_i[54] ),
    .I1(_06051_),
    .S(_09687_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20417_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(net169),
    .S(net1398),
    .Z(_06052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20418_ (.A1(_00969_),
    .A2(_04517_),
    .Z(_06053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20419_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .A2(net1613),
    .Z(_06054_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20420_ (.A1(net1673),
    .A2(_06052_),
    .B1(_06053_),
    .B2(_06054_),
    .C(net2029),
    .ZN(_06055_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20421_ (.A1(net2031),
    .A2(net169),
    .B1(_06045_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20422_ (.A1(net1725),
    .A2(_05868_),
    .B1(_06055_),
    .B2(_06056_),
    .ZN(_06057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20423_ (.I0(_05166_),
    .I1(_06057_),
    .S(net1750),
    .Z(_06058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20424_ (.I0(\ex_block_i.alu_i.imd_val_q_i[55] ),
    .I1(_06058_),
    .S(_09687_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20425_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(net2065),
    .S(net1398),
    .Z(_06059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20426_ (.A1(_00964_),
    .A2(_04522_),
    .Z(_06060_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20427_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .A2(net1613),
    .Z(_06061_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20428_ (.A1(net1673),
    .A2(_06059_),
    .B1(_06060_),
    .B2(_06061_),
    .C(net2029),
    .ZN(_06062_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20429_ (.A1(net2031),
    .A2(net2065),
    .B1(_06052_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20430_ (.A1(net1723),
    .A2(_05868_),
    .B1(_06062_),
    .B2(_06063_),
    .ZN(_06064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20431_ (.I0(_05184_),
    .I1(_06064_),
    .S(net1750),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20432_ (.I0(\ex_block_i.alu_i.imd_val_q_i[56] ),
    .I1(_06065_),
    .S(_09687_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20433_ (.I0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .I1(net1431),
    .S(net1398),
    .Z(_06066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20434_ (.A1(_00968_),
    .A2(_04522_),
    .Z(_06067_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20435_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .A2(net1613),
    .Z(_06068_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20436_ (.A1(net1673),
    .A2(_06066_),
    .B1(_06067_),
    .B2(_06068_),
    .C(net2029),
    .ZN(_06069_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20437_ (.A1(net2031),
    .A2(net1431),
    .B1(_06059_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06070_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20438_ (.A1(net1722),
    .A2(_05868_),
    .B1(_06069_),
    .B2(_06070_),
    .ZN(_06071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20439_ (.I0(_05211_),
    .I1(_06071_),
    .S(net1750),
    .Z(_06072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20440_ (.I0(\ex_block_i.alu_i.imd_val_q_i[57] ),
    .I1(_06072_),
    .S(_09687_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20441_ (.I0(net1792),
    .I1(net1499),
    .S(net1672),
    .Z(_06073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20442_ (.I0(\ex_block_i.alu_i.imd_val_q_i[5] ),
    .I1(_06073_),
    .S(net1548),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20443_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(net1409),
    .S(net1398),
    .Z(_06074_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20444_ (.A1(_00967_),
    .A2(_04522_),
    .Z(_06075_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20445_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .A2(net1613),
    .Z(_06076_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20446_ (.A1(net1673),
    .A2(_06074_),
    .B1(_06075_),
    .B2(_06076_),
    .C(net2029),
    .ZN(_06077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20447_ (.A1(net2031),
    .A2(net1409),
    .B1(_06066_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20448_ (.A1(net1721),
    .A2(_05868_),
    .B1(_06077_),
    .B2(_06078_),
    .ZN(_06079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20449_ (.I0(_05242_),
    .I1(_06079_),
    .S(net1750),
    .Z(_06080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20450_ (.I0(\ex_block_i.alu_i.imd_val_q_i[58] ),
    .I1(_06080_),
    .S(_09687_),
    .Z(_02935_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20451_ (.A1(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .A2(_05933_),
    .ZN(_06081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20452_ (.I0(\ex_block_i.alu_i.imd_val_q_i[59] ),
    .I1(net1429),
    .S(net1398),
    .Z(_06082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20453_ (.A1(_00969_),
    .A2(_04522_),
    .Z(_06083_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20454_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .A2(net1613),
    .Z(_06084_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20455_ (.A1(net1673),
    .A2(_06082_),
    .B1(_06083_),
    .B2(_06084_),
    .C(net2029),
    .ZN(_06085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20456_ (.A1(net2031),
    .A2(net1429),
    .B1(_06074_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20457_ (.A1(net1720),
    .A2(_05868_),
    .B1(_06085_),
    .B2(_06086_),
    .ZN(_06087_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20458_ (.A1(net1718),
    .A2(_06087_),
    .B(_05259_),
    .C(net1549),
    .ZN(_06088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20459_ (.A1(_06081_),
    .A2(_06088_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20460_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(net2138),
    .S(net1398),
    .Z(_06089_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20461_ (.A1(_00964_),
    .A2(_04527_),
    .Z(_06090_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20462_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .A2(net1613),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20463_ (.A1(net1673),
    .A2(_06089_),
    .B1(_06090_),
    .B2(_06091_),
    .C(net2029),
    .ZN(_06092_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20464_ (.A1(net2031),
    .A2(net2138),
    .B1(_06082_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20465_ (.A1(_09340_),
    .A2(_05868_),
    .B1(_06092_),
    .B2(_06093_),
    .ZN(_06094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20466_ (.I0(_05311_),
    .I1(_06094_),
    .S(net1750),
    .Z(_06095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20467_ (.I0(\ex_block_i.alu_i.imd_val_q_i[60] ),
    .I1(_06095_),
    .S(_09687_),
    .Z(_02937_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20468_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(net1408),
    .S(net1398),
    .Z(_06096_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20469_ (.A1(_00968_),
    .A2(_04527_),
    .Z(_06097_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20470_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .A2(net1613),
    .Z(_06098_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20471_ (.A1(net1673),
    .A2(_06096_),
    .B1(_06097_),
    .B2(_06098_),
    .C(net2029),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20472_ (.A1(net2031),
    .A2(net1408),
    .B1(_06089_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06100_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20473_ (.A1(net1754),
    .A2(_05868_),
    .B1(_06099_),
    .B2(_06100_),
    .C(net1718),
    .ZN(_06101_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20474_ (.A1(_05329_),
    .A2(_06101_),
    .Z(_06102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20475_ (.I0(\ex_block_i.alu_i.imd_val_q_i[61] ),
    .I1(_06102_),
    .S(net1549),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20476_ (.I0(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .I1(net2122),
    .S(net1398),
    .Z(_06103_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20477_ (.A1(net1673),
    .A2(_06103_),
    .ZN(_06104_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20478_ (.A1(_00967_),
    .A2(_04527_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .ZN(_06105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20479_ (.A1(net2031),
    .A2(net2122),
    .B1(_06096_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06106_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20480_ (.A1(net1752),
    .A2(_05868_),
    .Z(_06107_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _20481_ (.A1(_08196_),
    .A2(_06104_),
    .A3(_06105_),
    .B1(_06106_),
    .B2(_06107_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20482_ (.A1(_05849_),
    .A2(_06108_),
    .ZN(_06109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20483_ (.A1(\ex_block_i.alu_i.imd_val_q_i[62] ),
    .A2(_05933_),
    .B1(_09688_),
    .B2(_05373_),
    .ZN(_06110_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20484_ (.A1(_06109_),
    .A2(_06110_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20485_ (.A1(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .A2(net2051),
    .B(net1673),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20486_ (.A1(_00969_),
    .A2(_04527_),
    .B(net1613),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .ZN(_06112_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20487_ (.A1(_08196_),
    .A2(_06111_),
    .A3(_06112_),
    .Z(_06113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20488_ (.A1(net2031),
    .A2(net2051),
    .B1(_06103_),
    .B2(net2027),
    .C(net1806),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20489_ (.A1(_06113_),
    .A2(_06114_),
    .Z(_06115_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20490_ (.A1(_09467_),
    .A2(_05868_),
    .Z(_06116_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20491_ (.A1(net1718),
    .A2(_06115_),
    .A3(_06116_),
    .B(_05393_),
    .ZN(_06117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20492_ (.I0(\ex_block_i.alu_i.imd_val_q_i[63] ),
    .I1(_06117_),
    .S(_09687_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20493_ (.A1(net1806),
    .A2(_09677_),
    .ZN(_06118_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20494_ (.A1(_08194_),
    .A2(_04484_),
    .A3(_04462_),
    .Z(_06119_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20495_ (.A1(_06118_),
    .A2(_06119_),
    .Z(_06120_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20496_ (.A1(_01117_),
    .A2(_05370_),
    .Z(_06121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20497_ (.A1(_01124_),
    .A2(_06121_),
    .B(_01123_),
    .ZN(_06122_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20498_ (.A1(_01131_),
    .A2(_06122_),
    .Z(_06123_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20499_ (.A1(net1718),
    .A2(_06120_),
    .B1(_06123_),
    .B2(_05840_),
    .ZN(_06124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20500_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .I1(_06124_),
    .S(net1549),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20501_ (.A1(_01124_),
    .A2(_05390_),
    .Z(_06125_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20502_ (.A1(_01123_),
    .A2(_06125_),
    .Z(_06126_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20503_ (.A1(_01131_),
    .A2(_06126_),
    .B(_01130_),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20504_ (.A1(_00798_),
    .A2(_00749_),
    .Z(_06128_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20505_ (.A1(_01127_),
    .A2(_00794_),
    .A3(_06128_),
    .ZN(_06129_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20506_ (.A1(_00805_),
    .A2(_00807_),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20507_ (.A1(net1547),
    .A2(_00792_),
    .A3(_06130_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20508_ (.A1(_00800_),
    .A2(_00801_),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20509_ (.A1(net1537),
    .A2(_00793_),
    .ZN(_06133_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20510_ (.A1(_00802_),
    .A2(_00750_),
    .A3(_01125_),
    .ZN(_06134_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20511_ (.A1(_06132_),
    .A2(_06133_),
    .A3(_06134_),
    .ZN(_06135_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20512_ (.A1(_06129_),
    .A2(_06131_),
    .A3(_06135_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20513_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A2(net1716),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20514_ (.A1(net1710),
    .A2(_06137_),
    .Z(_06138_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20515_ (.A1(net1576),
    .A2(_06136_),
    .A3(_06138_),
    .ZN(_06139_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _20516_ (.A1(net1570),
    .A2(_06127_),
    .A3(_06139_),
    .ZN(_06140_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20517_ (.A1(net1718),
    .A2(_06118_),
    .B1(_06140_),
    .B2(_05840_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20518_ (.I0(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .I1(_06141_),
    .S(net1549),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20519_ (.I0(net1790),
    .I1(net1500),
    .S(net1672),
    .Z(_06142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20520_ (.I0(\ex_block_i.alu_i.imd_val_q_i[6] ),
    .I1(_06142_),
    .S(net1548),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20521_ (.I0(net1788),
    .I1(net1512),
    .S(net1672),
    .Z(_06143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20522_ (.I0(\ex_block_i.alu_i.imd_val_q_i[7] ),
    .I1(_06143_),
    .S(net1548),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20523_ (.I0(net1713),
    .I1(net1458),
    .S(net1672),
    .Z(_06144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20524_ (.I0(\ex_block_i.alu_i.imd_val_q_i[8] ),
    .I1(_06144_),
    .S(net1548),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20525_ (.I0(net1709),
    .I1(net1459),
    .S(net1672),
    .Z(_06145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20526_ (.I0(\ex_block_i.alu_i.imd_val_q_i[9] ),
    .I1(_06145_),
    .S(net1548),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20527_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_09901_),
    .B(_09497_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20528_ (.A1(_09938_),
    .A2(_06146_),
    .Z(_06147_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20529_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(net1746),
    .B1(_06147_),
    .B2(\cs_registers_i.csr_mtvec_o[10] ),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20530_ (.I(_06148_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20531_ (.A1(net6),
    .A2(net1618),
    .B1(net1747),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C(_06149_),
    .ZN(_06150_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20532_ (.A1(_08509_),
    .A2(_05727_),
    .B(_10012_),
    .C(_06150_),
    .ZN(_06151_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20533_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .A2(_10012_),
    .Z(_06152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20534_ (.A1(_06151_),
    .A2(_06152_),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20535_ (.A1(\cs_registers_i.csr_mtvec_o[9] ),
    .A2(_06147_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20536_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[9] ),
    .ZN(_06155_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20537_ (.A1(_08455_),
    .A2(_05727_),
    .B(_06154_),
    .C(_06155_),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20538_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_09902_),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .ZN(_06157_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20539_ (.A1(_10074_),
    .A2(_06157_),
    .B(_03901_),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20540_ (.I0(net29),
    .I1(_06156_),
    .S(_06158_),
    .Z(_06159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20541_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .I1(_06159_),
    .S(_10012_),
    .Z(_06160_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20542_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _20543_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[4] ),
    .C1(_04021_),
    .C2(_09945_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20544_ (.I(_06162_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20545_ (.A1(net1809),
    .A2(net1454),
    .B(net1589),
    .C(_06163_),
    .ZN(_06164_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20546_ (.A1(_06161_),
    .A2(net1589),
    .B(_06164_),
    .ZN(_06165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20547_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .ZN(_06166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20548_ (.A1(net1809),
    .A2(net1499),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20549_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(net1747),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20550_ (.A1(_10012_),
    .A2(_04031_),
    .A3(_06167_),
    .A4(_06168_),
    .Z(_06169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20551_ (.A1(_06166_),
    .A2(net1589),
    .B(_06169_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20552_ (.A1(_01375_),
    .A2(_06165_),
    .A3(_06170_),
    .Z(_06171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20553_ (.A1(net1500),
    .A2(net1809),
    .Z(_06172_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20554_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(net1747),
    .Z(_06173_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20555_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(net1746),
    .Z(_06174_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20556_ (.A1(_04037_),
    .A2(_06173_),
    .A3(_06174_),
    .Z(_06175_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20557_ (.A1(_08471_),
    .A2(_08472_),
    .A3(net1809),
    .Z(_06176_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20558_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(_09965_),
    .B1(_06147_),
    .B2(\cs_registers_i.csr_mtvec_o[8] ),
    .ZN(_06177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20559_ (.I(_06177_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20560_ (.A1(net28),
    .A2(net1618),
    .B1(net1747),
    .B2(\cs_registers_i.csr_depc_o[8] ),
    .C(_06178_),
    .ZN(_06179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20561_ (.I(_06179_),
    .ZN(_06180_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _20562_ (.A1(_06172_),
    .A2(_06175_),
    .B1(_06176_),
    .B2(_06180_),
    .C(_09957_),
    .ZN(_06181_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20563_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A3(net1589),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20564_ (.A1(net1512),
    .A2(net1809),
    .ZN(_06183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20565_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[7] ),
    .ZN(_06184_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20566_ (.A1(_06158_),
    .A2(_06183_),
    .A3(_06184_),
    .ZN(_06185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20567_ (.I0(_06185_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .S(net1589),
    .Z(_06186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20568_ (.I(_06186_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20569_ (.A1(_06181_),
    .A2(_06182_),
    .B(_06187_),
    .ZN(_06188_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20570_ (.A1(_06171_),
    .A2(_06188_),
    .Z(_06189_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20571_ (.A1(_06160_),
    .A2(_06189_),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20572_ (.A1(_06153_),
    .A2(_06190_),
    .ZN(_06191_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20573_ (.A1(net1589),
    .A2(_10081_),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net1410),
    .Z(data_addr_o[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net2278),
    .Z(data_addr_o[20]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20576_ (.I0(_06191_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .S(net1542),
    .Z(_02947_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20577_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_09952_),
    .B(_09938_),
    .ZN(_06195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20578_ (.A1(_03901_),
    .A2(_06195_),
    .ZN(_06196_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20579_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_09922_),
    .A3(_09997_),
    .B(_06196_),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20580_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_09965_),
    .ZN(_06198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20581_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(net1747),
    .ZN(_06199_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20582_ (.A1(_06197_),
    .A2(_06198_),
    .A3(_06199_),
    .Z(_06200_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20583_ (.A1(_08496_),
    .A2(_08497_),
    .A3(_05727_),
    .B(_06200_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20584_ (.I0(net7),
    .I1(_06201_),
    .S(_06158_),
    .Z(_06202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20585_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .I1(_06202_),
    .S(_10012_),
    .Z(_06203_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20586_ (.A1(_01373_),
    .A2(_01374_),
    .A3(_06165_),
    .Z(_06204_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20587_ (.A1(_06170_),
    .A2(_06204_),
    .Z(_06205_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20588_ (.A1(_06188_),
    .A2(_06205_),
    .Z(_06206_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20589_ (.A1(_06153_),
    .A2(_06160_),
    .A3(_06206_),
    .Z(_06207_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20590_ (.A1(_06203_),
    .A2(_06207_),
    .Z(_06208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20591_ (.I0(_06208_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .S(net1542),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20592_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20593_ (.A1(\cs_registers_i.csr_mtvec_o[12] ),
    .A2(_06147_),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20594_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[12] ),
    .ZN(_06211_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20595_ (.A1(net8),
    .A2(net1618),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20596_ (.A1(_06210_),
    .A2(_06211_),
    .A3(_06212_),
    .ZN(_06213_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20597_ (.A1(net1809),
    .A2(net1449),
    .B(net1589),
    .C(_06213_),
    .ZN(_06214_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20598_ (.A1(_06209_),
    .A2(net1589),
    .B(_06214_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20599_ (.A1(_06151_),
    .A2(_06152_),
    .A3(_06160_),
    .A4(_06203_),
    .Z(_06216_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20600_ (.A1(_06189_),
    .A2(_06216_),
    .ZN(_06217_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20601_ (.A1(_06215_),
    .A2(_06217_),
    .ZN(_06218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20602_ (.I0(_06218_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .S(net1542),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20603_ (.A1(net9),
    .A2(_06158_),
    .ZN(_06219_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net1436),
    .Z(data_addr_o[19]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20605_ (.A1(\cs_registers_i.csr_mtvec_o[13] ),
    .A2(_06147_),
    .ZN(_06221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20606_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[13] ),
    .ZN(_06222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20607_ (.A1(_06221_),
    .A2(_06222_),
    .ZN(_06223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20608_ (.A1(net1450),
    .A2(net1809),
    .B(net1618),
    .C(_06223_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20609_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .A2(net1589),
    .ZN(_06225_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20610_ (.A1(net1589),
    .A2(_06219_),
    .A3(_06224_),
    .B(_06225_),
    .ZN(_06226_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20611_ (.A1(_06188_),
    .A2(_06205_),
    .A3(_06215_),
    .A4(_06216_),
    .Z(_06227_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20612_ (.A1(_06226_),
    .A2(_06227_),
    .Z(_06228_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net1435),
    .Z(data_addr_o[18]));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20614_ (.I0(_06228_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .S(net1542),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net2288),
    .Z(data_addr_o[17]));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20616_ (.A1(_06188_),
    .A2(_06215_),
    .A3(_06216_),
    .A4(_06226_),
    .Z(_06231_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20617_ (.A1(_06171_),
    .A2(_06231_),
    .Z(_06232_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20618_ (.A1(_01371_),
    .A2(_06232_),
    .Z(_06233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20619_ (.I0(_10081_),
    .I1(_06233_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .Z(_06234_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net1446),
    .Z(data_addr_o[16]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20621_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(net1589),
    .ZN(_06236_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20622_ (.A1(net1456),
    .A2(net1809),
    .Z(_06237_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20623_ (.A1(\cs_registers_i.csr_mtvec_o[14] ),
    .A2(_06147_),
    .ZN(_06238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20624_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20625_ (.A1(_06238_),
    .A2(_06239_),
    .ZN(_06240_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20626_ (.A1(net10),
    .A2(net1618),
    .Z(_06241_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20627_ (.A1(_06241_),
    .A2(_06240_),
    .A3(_06237_),
    .B(net1581),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20628_ (.A1(_06232_),
    .A2(_06242_),
    .Z(_06243_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20629_ (.A1(net1589),
    .A2(_06234_),
    .B1(_06236_),
    .B2(_06243_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20630_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .A2(net1589),
    .ZN(_06244_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20631_ (.A1(\cs_registers_i.csr_mtvec_o[15] ),
    .A2(_06147_),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20632_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[15] ),
    .ZN(_06246_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20633_ (.A1(net1448),
    .A2(net1809),
    .ZN(_06247_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20634_ (.A1(_06158_),
    .A2(_06245_),
    .A3(_06246_),
    .A4(_06247_),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _20635_ (.A1(net11),
    .A2(_06158_),
    .B(_06248_),
    .C(net1581),
    .ZN(_06249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20636_ (.A1(_06249_),
    .A2(_06244_),
    .ZN(_06250_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20637_ (.A1(_06236_),
    .A2(_06242_),
    .ZN(_06251_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20638_ (.A1(_06205_),
    .A2(_06231_),
    .A3(_06251_),
    .Z(_06252_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20639_ (.A1(_06250_),
    .A2(_06252_),
    .Z(_06253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20640_ (.I0(_06253_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .S(_06192_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20641_ (.A1(_09922_),
    .A2(_09997_),
    .Z(_06254_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20642_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_06254_),
    .B(_06196_),
    .ZN(_06255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20643_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_09965_),
    .ZN(_06256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20644_ (.A1(_06255_),
    .A2(_06256_),
    .ZN(_06257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20645_ (.A1(net12),
    .A2(net1618),
    .B1(net1747),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .C(_06257_),
    .ZN(_06258_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20646_ (.A1(net1455),
    .A2(_08839_),
    .A3(_05727_),
    .B(_06258_),
    .ZN(_06259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20647_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .I1(_06259_),
    .S(_10012_),
    .Z(_06260_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20648_ (.A1(_06232_),
    .A2(_06251_),
    .A3(_06250_),
    .Z(_06261_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20649_ (.A1(_06260_),
    .A2(_06261_),
    .Z(_06262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20650_ (.I0(_06262_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .S(_06192_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20651_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(_06147_),
    .Z(_06263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20652_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[17] ),
    .C(_06263_),
    .ZN(_06264_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20653_ (.A1(net1447),
    .A2(net1809),
    .B1(net1618),
    .B2(net13),
    .ZN(_06265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20654_ (.A1(_06264_),
    .A2(_06265_),
    .B(net1589),
    .ZN(_06266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20655_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(net1589),
    .Z(_06267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20656_ (.A1(_06267_),
    .A2(_06266_),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20657_ (.A1(_06251_),
    .A2(_06250_),
    .A3(_06260_),
    .Z(_06269_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20658_ (.A1(_06231_),
    .A2(_06269_),
    .Z(_06270_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20659_ (.A1(_06205_),
    .A2(_06270_),
    .ZN(_06271_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20660_ (.A1(_06268_),
    .A2(_06271_),
    .ZN(_06272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20661_ (.I0(_06272_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .S(_06192_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net1448),
    .Z(data_addr_o[15]));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20663_ (.A1(\cs_registers_i.csr_mtvec_o[18] ),
    .A2(_06147_),
    .Z(_06274_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20664_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[18] ),
    .C(_06274_),
    .ZN(_06275_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20665_ (.I(_06275_),
    .ZN(_06276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20666_ (.A1(net1435),
    .A2(net1809),
    .B1(net1618),
    .B2(net14),
    .C(_06276_),
    .ZN(_06277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20667_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .A2(net1589),
    .ZN(_06278_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20668_ (.A1(net1589),
    .A2(_06277_),
    .B(_06278_),
    .ZN(_06279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20669_ (.A1(_06232_),
    .A2(_06269_),
    .A3(_06268_),
    .Z(_06280_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20670_ (.A1(_06279_),
    .A2(_06280_),
    .Z(_06281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20671_ (.I0(_06281_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .S(_06192_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20672_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .ZN(_06282_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20673_ (.A1(\cs_registers_i.csr_mtvec_o[19] ),
    .A2(_06147_),
    .ZN(_06283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20674_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[19] ),
    .ZN(_06284_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20675_ (.A1(net15),
    .A2(net1618),
    .ZN(_06285_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20676_ (.A1(_06283_),
    .A2(_06284_),
    .A3(_06285_),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20677_ (.A1(net1436),
    .A2(net1809),
    .B(net1589),
    .C(_06286_),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20678_ (.A1(_06282_),
    .A2(net1589),
    .B(_06287_),
    .ZN(_06288_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20679_ (.A1(_06205_),
    .A2(_06279_),
    .Z(_06289_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20680_ (.A1(_06268_),
    .A2(_06270_),
    .A3(_06289_),
    .Z(_06290_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20681_ (.A1(_06288_),
    .A2(_06290_),
    .ZN(_06291_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20682_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(_06192_),
    .ZN(_06292_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20683_ (.A1(_06192_),
    .A2(_06291_),
    .B(_06292_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20684_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .A2(net1589),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20685_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_06254_),
    .Z(_06294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20686_ (.A1(\cs_registers_i.csr_mepc_o[20] ),
    .A2(net1746),
    .B1(_06196_),
    .B2(_06294_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20687_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(net1747),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20688_ (.A1(_06295_),
    .A2(_06296_),
    .ZN(_06297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20689_ (.A1(net1433),
    .A2(net1809),
    .B1(net1618),
    .B2(net16),
    .C(_06297_),
    .ZN(_06298_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20690_ (.A1(net1589),
    .A2(_06298_),
    .Z(_06299_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20691_ (.A1(_06232_),
    .A2(_06269_),
    .ZN(_06300_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20692_ (.A1(_06268_),
    .A2(_06279_),
    .A3(_06288_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20693_ (.A1(_06300_),
    .A2(_06301_),
    .Z(_06302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20694_ (.A1(_06293_),
    .A2(_06299_),
    .B(_06302_),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20695_ (.A1(_06302_),
    .A2(_06299_),
    .Z(_06304_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net2292),
    .Z(data_addr_o[14]));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20697_ (.A1(_10081_),
    .A2(_06302_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .C(net1589),
    .ZN(_06306_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20698_ (.A1(net1542),
    .A2(_06303_),
    .A3(_06304_),
    .B(_06306_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20699_ (.A1(\cs_registers_i.csr_mtvec_o[21] ),
    .A2(_06147_),
    .Z(_06307_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20700_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[21] ),
    .C(_06307_),
    .ZN(_06308_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20701_ (.I(_06308_),
    .ZN(_06309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20702_ (.A1(net17),
    .A2(net1618),
    .B(_06309_),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _20703_ (.A1(_09015_),
    .A2(net1434),
    .A3(_05727_),
    .B(_06310_),
    .ZN(_06311_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_4 _20704_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .I1(_06311_),
    .S(_10012_),
    .Z(_06312_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20705_ (.A1(_06293_),
    .A2(_06299_),
    .Z(_06313_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20706_ (.A1(_06301_),
    .A2(_06313_),
    .ZN(_06314_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20707_ (.A1(_06205_),
    .A2(_06231_),
    .A3(_06269_),
    .A4(_06314_),
    .Z(_06315_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20708_ (.A1(_06312_),
    .A2(_06315_),
    .Z(_06316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20709_ (.I0(_06316_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .S(net1542),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20710_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(net1589),
    .ZN(_06317_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20711_ (.A1(\cs_registers_i.csr_mtvec_o[22] ),
    .A2(_06147_),
    .Z(_06318_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20712_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[22] ),
    .C(_06318_),
    .ZN(_06319_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20713_ (.I(_06319_),
    .ZN(_06320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20714_ (.A1(net1432),
    .A2(net1809),
    .B1(net1618),
    .B2(net18),
    .C(_06320_),
    .ZN(_06321_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20715_ (.A1(net1589),
    .A2(_06321_),
    .Z(_06322_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20716_ (.A1(_06232_),
    .A2(_06269_),
    .A3(_06314_),
    .Z(_06323_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20717_ (.A1(_06312_),
    .A2(_06323_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20718_ (.A1(_06317_),
    .A2(_06322_),
    .B(_06324_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20719_ (.A1(_06324_),
    .A2(_06322_),
    .Z(_06326_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20720_ (.A1(_10081_),
    .A2(_06324_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .C(net1589),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20721_ (.A1(net1542),
    .A2(_06325_),
    .A3(_06326_),
    .B(_06327_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20722_ (.A1(\cs_registers_i.csr_mepc_o[23] ),
    .A2(net1746),
    .B1(_06147_),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20723_ (.I(_06328_),
    .ZN(_06329_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20724_ (.A1(net19),
    .A2(net1618),
    .B1(net1747),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C(_06329_),
    .ZN(_06330_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20725_ (.A1(_09105_),
    .A2(_09106_),
    .A3(_05727_),
    .B(_06330_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20726_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .I1(_06331_),
    .S(_10012_),
    .Z(_06332_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20727_ (.A1(net1589),
    .A2(_06321_),
    .B(_06317_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20728_ (.A1(_06312_),
    .A2(_06315_),
    .A3(_06333_),
    .Z(_06334_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20729_ (.A1(_06332_),
    .A2(_06334_),
    .Z(_06335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20730_ (.I0(_06335_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .S(net1542),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20731_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(net1589),
    .ZN(_06336_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20732_ (.A1(\cs_registers_i.csr_mtvec_o[24] ),
    .A2(_06147_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20733_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .ZN(_06338_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20734_ (.A1(_06337_),
    .A2(_06338_),
    .ZN(_06339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20735_ (.A1(net170),
    .A2(net1809),
    .B1(net1618),
    .B2(net20),
    .C(_06339_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20736_ (.A1(net1589),
    .A2(_06340_),
    .Z(_06341_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20737_ (.A1(_06312_),
    .A2(_06333_),
    .A3(_06332_),
    .Z(_06342_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20738_ (.A1(_06323_),
    .A2(_06342_),
    .ZN(_06343_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20739_ (.A1(_06336_),
    .A2(_06341_),
    .B(_06343_),
    .ZN(_06344_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20740_ (.A1(_06343_),
    .A2(_06341_),
    .Z(_06345_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20741_ (.A1(_10081_),
    .A2(_06343_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .C(net1589),
    .ZN(_06346_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20742_ (.A1(net1542),
    .A2(_06344_),
    .A3(_06345_),
    .B(_06346_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20743_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .A2(net1589),
    .ZN(_06347_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20744_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_06254_),
    .Z(_06348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20745_ (.A1(\cs_registers_i.csr_mepc_o[25] ),
    .A2(_09965_),
    .B1(_06196_),
    .B2(_06348_),
    .ZN(_06349_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20746_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(net1747),
    .ZN(_06350_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20747_ (.A1(_06349_),
    .A2(_06350_),
    .ZN(_06351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20748_ (.A1(net1431),
    .A2(net1809),
    .B1(net1618),
    .B2(net21),
    .C(_06351_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20749_ (.A1(_06352_),
    .A2(net1589),
    .Z(_06353_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20750_ (.A1(net1589),
    .A2(_06340_),
    .B(_06336_),
    .ZN(_06354_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20751_ (.A1(_06342_),
    .A2(_06354_),
    .Z(_06355_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20752_ (.A1(_06315_),
    .A2(_06355_),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20753_ (.A1(_06347_),
    .A2(net2276),
    .B(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20754_ (.A1(_06356_),
    .A2(net2276),
    .Z(_06358_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20755_ (.A1(_10081_),
    .A2(_06356_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .C(net1589),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20756_ (.A1(net1542),
    .A2(_06357_),
    .A3(_06358_),
    .B(_06359_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20757_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(_06147_),
    .Z(_06360_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20758_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .C(_06360_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20759_ (.A1(net22),
    .A2(net1618),
    .ZN(_06362_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20760_ (.A1(net1428),
    .A2(_05727_),
    .B(_06361_),
    .C(_06362_),
    .ZN(_06363_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20761_ (.A1(_06363_),
    .A2(net1581),
    .ZN(_06364_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20762_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(net1589),
    .ZN(_06365_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20763_ (.A1(_06365_),
    .A2(_06364_),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20764_ (.A1(_06347_),
    .A2(_06353_),
    .ZN(_06367_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20765_ (.A1(_06323_),
    .A2(_06355_),
    .A3(_06367_),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20766_ (.A1(_06366_),
    .A2(_06368_),
    .Z(_06369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20767_ (.I0(_06369_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .S(net1542),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20768_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .A2(net1589),
    .ZN(_06370_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20769_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_06254_),
    .Z(_06371_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20770_ (.A1(\cs_registers_i.csr_mepc_o[27] ),
    .A2(_09965_),
    .B1(_06196_),
    .B2(_06371_),
    .ZN(_06372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20771_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(net1747),
    .ZN(_06373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20772_ (.A1(_06372_),
    .A2(_06373_),
    .ZN(_06374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20773_ (.A1(net173),
    .A2(net1809),
    .B1(net1618),
    .B2(net23),
    .C(_06374_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20774_ (.A1(net1589),
    .A2(_06375_),
    .Z(_06376_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20775_ (.A1(_06370_),
    .A2(_06376_),
    .ZN(_06377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20776_ (.I(_06377_),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20777_ (.A1(_10081_),
    .A2(_06370_),
    .B(_06376_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _20778_ (.I(_06313_),
    .ZN(_06380_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20779_ (.A1(_06268_),
    .A2(_06288_),
    .A3(_06380_),
    .Z(_06381_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20780_ (.A1(_06342_),
    .A2(_06354_),
    .A3(_06367_),
    .A4(_06366_),
    .Z(_06382_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20781_ (.A1(_06270_),
    .A2(_06289_),
    .A3(_06381_),
    .A4(_06382_),
    .Z(_06383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20782_ (.I0(_06378_),
    .I1(_06379_),
    .S(_06383_),
    .Z(_06384_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20783_ (.A1(_06192_),
    .A2(_06370_),
    .B(_06384_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20784_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .ZN(_06385_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net1450),
    .Z(data_addr_o[13]));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20786_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_06254_),
    .Z(_06387_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20787_ (.A1(\cs_registers_i.csr_mepc_o[28] ),
    .A2(_09965_),
    .B1(_06196_),
    .B2(_06387_),
    .ZN(_06388_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20788_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(net1747),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20789_ (.A1(_06388_),
    .A2(_06389_),
    .ZN(_06390_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20790_ (.A1(net1809),
    .A2(net1407),
    .B1(net1618),
    .B2(net24),
    .C(_06390_),
    .ZN(_06391_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20791_ (.A1(_06391_),
    .A2(net1589),
    .Z(_06392_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20792_ (.A1(_06385_),
    .A2(_10012_),
    .B(_06392_),
    .ZN(_06393_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20793_ (.A1(_06323_),
    .A2(_06382_),
    .A3(_06377_),
    .Z(_06394_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20794_ (.A1(_06393_),
    .A2(_06394_),
    .Z(_06395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20795_ (.I0(_06395_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .S(_06192_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20796_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(_06147_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20797_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[29] ),
    .ZN(_06397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20798_ (.A1(_06396_),
    .A2(_06397_),
    .ZN(_06398_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20799_ (.A1(net1809),
    .A2(net175),
    .B1(net1618),
    .B2(net25),
    .C(_06398_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20800_ (.A1(_06399_),
    .A2(net1589),
    .Z(_06400_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20801_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .A2(net1589),
    .ZN(_06401_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20802_ (.A1(_06400_),
    .A2(_06401_),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20803_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .ZN(_06403_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20804_ (.A1(_06403_),
    .A2(_06376_),
    .B1(_06392_),
    .B2(_06385_),
    .ZN(_06404_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20805_ (.A1(_06376_),
    .A2(net2478),
    .B(_10012_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20806_ (.A1(_06315_),
    .A2(_06382_),
    .A3(_06404_),
    .A4(_06405_),
    .Z(_06406_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20807_ (.A1(_06402_),
    .A2(_06406_),
    .Z(_06407_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20808_ (.I0(_06407_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .S(_06192_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20809_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .S(net1542),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20810_ (.A1(\cs_registers_i.csr_mtvec_o[30] ),
    .A2(_06147_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20811_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[30] ),
    .ZN(_06409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20812_ (.A1(_06408_),
    .A2(_06409_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20813_ (.A1(net1406),
    .A2(net1809),
    .B1(net1618),
    .B2(net26),
    .C(_06410_),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20814_ (.A1(_06411_),
    .A2(net1589),
    .Z(_06412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20815_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .A2(net1589),
    .ZN(_06413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20816_ (.A1(_06412_),
    .A2(_06413_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20817_ (.A1(_06382_),
    .A2(_06402_),
    .A3(_06404_),
    .A4(_06405_),
    .Z(_06415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20818_ (.A1(_06323_),
    .A2(_06415_),
    .ZN(_06416_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20819_ (.A1(_06414_),
    .A2(_06416_),
    .ZN(_06417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20820_ (.I0(_06417_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .S(net1542),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20821_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_06147_),
    .ZN(_06418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20822_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(net1747),
    .B1(net1746),
    .B2(\cs_registers_i.csr_mepc_o[31] ),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20823_ (.A1(_06418_),
    .A2(_06419_),
    .ZN(_06420_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _20824_ (.A1(net178),
    .A2(net1809),
    .B1(net1618),
    .B2(net27),
    .C(_06420_),
    .ZN(_06421_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _20825_ (.A1(_06421_),
    .A2(net1589),
    .Z(_06422_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20826_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .A2(net1589),
    .ZN(_06423_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _20827_ (.A1(_06422_),
    .A2(_06423_),
    .ZN(_06424_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20828_ (.A1(_06315_),
    .A2(_06414_),
    .A3(_06415_),
    .Z(_06425_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20829_ (.A1(_06424_),
    .A2(_06425_),
    .Z(_06426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20830_ (.I0(_06426_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .S(net1542),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20831_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .S(net1542),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20832_ (.A1(_01375_),
    .A2(_06165_),
    .Z(_06427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20833_ (.I0(_06427_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .S(net1542),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20834_ (.A1(_06170_),
    .A2(_06204_),
    .Z(_06428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20835_ (.I0(_06428_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .S(net1542),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _20836_ (.A1(_06172_),
    .A2(_06175_),
    .B(_09957_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20837_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(net1589),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20838_ (.A1(_06429_),
    .A2(_06430_),
    .ZN(_06431_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20839_ (.A1(_06171_),
    .A2(_06431_),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20840_ (.I0(_06432_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .S(net1542),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20841_ (.A1(_06205_),
    .A2(_06431_),
    .Z(_06433_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20842_ (.A1(_06187_),
    .A2(_06433_),
    .ZN(_06434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20843_ (.I0(_06434_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .S(net1542),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20844_ (.A1(_06176_),
    .A2(_06180_),
    .ZN(_06435_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20845_ (.A1(_06171_),
    .A2(_06186_),
    .A3(_06431_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20846_ (.A1(_06435_),
    .A2(_06436_),
    .B(_06189_),
    .ZN(_06437_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20847_ (.A1(net1589),
    .A2(_06437_),
    .Z(_06438_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20848_ (.A1(_01371_),
    .A2(_06189_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20849_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(_10012_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20850_ (.A1(_10081_),
    .A2(_06436_),
    .B(_06440_),
    .ZN(_06441_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20851_ (.A1(_06438_),
    .A2(_06439_),
    .A3(_06441_),
    .Z(_02975_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20852_ (.A1(_06160_),
    .A2(_06206_),
    .Z(_06442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20853_ (.I0(_06442_),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .S(net1542),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20854_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net133),
    .ZN(_06443_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20855_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_06443_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20856_ (.A1(_10023_),
    .A2(_06444_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net2298),
    .Z(data_addr_o[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net1457),
    .Z(data_addr_o[11]));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20859_ (.A1(net2025),
    .A2(_06444_),
    .ZN(_06448_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20860_ (.A1(net2024),
    .A2(_06448_),
    .Z(_06449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20861_ (.I(net2024),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20862_ (.A1(_10026_),
    .A2(_10033_),
    .Z(_06451_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20863_ (.A1(net2026),
    .A2(_06450_),
    .A3(_06451_),
    .A4(_06448_),
    .Z(_06452_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net1451),
    .Z(data_addr_o[10]));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20865_ (.A1(net2026),
    .A2(_06451_),
    .B(_06444_),
    .C(net2025),
    .ZN(_06454_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20866_ (.A1(_06452_),
    .A2(_06454_),
    .ZN(_06455_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20867_ (.A1(_10027_),
    .A2(_03436_),
    .A3(_06455_),
    .ZN(_06456_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _20868_ (.A1(net1809),
    .A2(_05777_),
    .B(_05767_),
    .C(_06456_),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20869_ (.A1(net1393),
    .A2(_06457_),
    .Z(_06458_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net155),
    .Z(core_sleep_o));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20871_ (.I0(_06445_),
    .I1(_06449_),
    .S(_06458_),
    .Z(_06460_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input155 (.I(test_en_i),
    .Z(net154));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 input154 (.I(rst_ni),
    .Z(net153));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20874_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .ZN(_06463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20875_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .ZN(_06464_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20876_ (.A1(net2024),
    .A2(_10027_),
    .A3(_03436_),
    .A4(_06455_),
    .ZN(_06465_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20877_ (.A1(net1809),
    .A2(_05777_),
    .B(_05767_),
    .C(_06465_),
    .ZN(_06466_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20878_ (.A1(net1394),
    .A2(net1501),
    .Z(_06467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20879_ (.I0(_06463_),
    .I1(_06464_),
    .S(_06467_),
    .Z(_06468_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20880_ (.A1(net1393),
    .A2(_06457_),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input153 (.I(irq_timer_i),
    .Z(net152));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input152 (.I(irq_software_i),
    .Z(net151));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input151 (.I(irq_nm_i),
    .Z(net150));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20884_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_06443_),
    .Z(_06473_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input150 (.I(irq_fast_i[9]),
    .Z(net149));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _20886_ (.A1(_10023_),
    .A2(net2024),
    .A3(net99),
    .A4(net1819),
    .Z(_06475_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20887_ (.A1(_10023_),
    .A2(net2024),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20888_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(net1819),
    .A3(_06476_),
    .Z(_06477_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20889_ (.A1(_03402_),
    .A2(_03423_),
    .B(_03429_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input149 (.I(irq_fast_i[8]),
    .Z(net148));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input148 (.I(irq_fast_i[7]),
    .Z(net147));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _20892_ (.A1(net2025),
    .A2(net2024),
    .A3(net99),
    .A4(net1819),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20893_ (.A1(_06478_),
    .A2(_05769_),
    .A3(_06456_),
    .B(_06481_),
    .ZN(_06482_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20894_ (.A1(_06469_),
    .A2(_06475_),
    .B(_06477_),
    .C(_06482_),
    .ZN(_06483_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20895_ (.A1(_06460_),
    .A2(_06468_),
    .B(_06483_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input147 (.I(irq_fast_i[6]),
    .Z(net146));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20897_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(net2023),
    .Z(_06485_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20898_ (.A1(net2024),
    .A2(_06448_),
    .ZN(_06486_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20899_ (.A1(net2024),
    .A2(_06444_),
    .B(net2023),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20900_ (.I(_06487_),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20901_ (.I0(_06486_),
    .I1(_06488_),
    .S(_06458_),
    .Z(_06489_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input146 (.I(irq_fast_i[5]),
    .Z(net145));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input145 (.I(irq_fast_i[4]),
    .Z(net144));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20904_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .I1(_06485_),
    .S(net1378),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20905_ (.A1(_06450_),
    .A2(net2023),
    .A3(net1819),
    .Z(_06492_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input144 (.I(irq_fast_i[3]),
    .Z(net143));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20907_ (.I0(net99),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(net1805),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input143 (.I(irq_fast_i[2]),
    .Z(net142));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input142 (.I(irq_fast_i[1]),
    .Z(net141));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20910_ (.A1(net1539),
    .A2(net1809),
    .Z(_06496_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _20911_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(net1747),
    .B1(_09965_),
    .B2(\cs_registers_i.csr_mepc_o[1] ),
    .C(_06496_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20912_ (.A1(_03436_),
    .A2(_06455_),
    .Z(_06498_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20913_ (.I(_06498_),
    .ZN(_06499_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20914_ (.A1(net1809),
    .A2(_05777_),
    .B(_05767_),
    .C(_06499_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input141 (.I(irq_fast_i[14]),
    .Z(net140));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20916_ (.A1(net1393),
    .A2(_06500_),
    .ZN(_06502_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input140 (.I(irq_fast_i[13]),
    .Z(net139));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20918_ (.A1(_06451_),
    .A2(net1385),
    .B(net2026),
    .ZN(_06504_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20919_ (.I(_10027_),
    .ZN(_06505_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _20920_ (.A1(net1393),
    .A2(_06500_),
    .Z(_06506_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input139 (.I(irq_fast_i[12]),
    .Z(net138));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input138 (.I(irq_fast_i[11]),
    .Z(net137));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input137 (.I(irq_fast_i[10]),
    .Z(net136));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20924_ (.A1(_06505_),
    .A2(net1384),
    .B(_10012_),
    .ZN(_06510_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20925_ (.A1(_10012_),
    .A2(_06497_),
    .B1(_06504_),
    .B2(_06510_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20926_ (.I(\cs_registers_i.pc_if_i[3] ),
    .ZN(_06511_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20927_ (.A1(_06511_),
    .A2(_00812_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20928_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(\cs_registers_i.pc_if_i[5] ),
    .A3(\cs_registers_i.pc_if_i[6] ),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20929_ (.A1(\cs_registers_i.pc_if_i[7] ),
    .A2(_06513_),
    .Z(_06514_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20930_ (.A1(\cs_registers_i.pc_if_i[8] ),
    .A2(_06514_),
    .Z(_06515_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20931_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_06515_),
    .Z(_06516_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20932_ (.A1(\cs_registers_i.pc_if_i[10] ),
    .A2(_06516_),
    .Z(_06517_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20933_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06512_),
    .A4(_06517_),
    .Z(_06518_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _20934_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(_06518_),
    .Z(_06519_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _20935_ (.I0(_06202_),
    .I1(_06519_),
    .S(net1589),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input136 (.I(irq_fast_i[0]),
    .Z(net135));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20937_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(_06517_),
    .Z(_06521_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20938_ (.I(_01133_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20939_ (.A1(net2026),
    .A2(_01134_),
    .A3(_10034_),
    .ZN(_06523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20940_ (.A1(_06522_),
    .A2(_06523_),
    .B(_06511_),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20941_ (.A1(_06521_),
    .A2(_06524_),
    .Z(_06525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _20942_ (.A1(net1383),
    .A2(_06525_),
    .B(\cs_registers_i.pc_if_i[12] ),
    .C(net1581),
    .ZN(_06526_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20943_ (.A1(\cs_registers_i.pc_if_i[12] ),
    .A2(net1589),
    .A3(net1383),
    .A4(_06525_),
    .Z(_06527_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _20944_ (.A1(_06214_),
    .A2(_06526_),
    .A3(_06527_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input135 (.I(irq_external_i),
    .Z(net134));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20946_ (.A1(\cs_registers_i.pc_if_i[12] ),
    .A2(_06512_),
    .A3(_06521_),
    .Z(_06529_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20947_ (.A1(net1383),
    .A2(_06529_),
    .Z(_06530_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20948_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(net1589),
    .ZN(_06531_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20949_ (.I(\cs_registers_i.pc_if_i[13] ),
    .ZN(_06532_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input134 (.I(instr_rvalid_i),
    .Z(net133));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _20951_ (.A1(_06532_),
    .A2(net1589),
    .A3(net1383),
    .A4(_06529_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20952_ (.A1(net1589),
    .A2(_06219_),
    .A3(_06224_),
    .Z(_06535_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _20953_ (.A1(_06530_),
    .A2(_06531_),
    .B(_06534_),
    .C(_06535_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20954_ (.I(\cs_registers_i.pc_if_i[14] ),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20955_ (.A1(\cs_registers_i.pc_if_i[12] ),
    .A2(_06521_),
    .A3(_06524_),
    .ZN(_06537_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20956_ (.A1(_06532_),
    .A2(_06537_),
    .B(_06242_),
    .ZN(_06538_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20957_ (.A1(net1581),
    .A2(net1383),
    .B(_06538_),
    .ZN(_06539_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20958_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(\cs_registers_i.pc_if_i[14] ),
    .ZN(_06540_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20959_ (.A1(net1386),
    .A2(_06537_),
    .A3(_06540_),
    .B(net1589),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20960_ (.A1(_06536_),
    .A2(_06539_),
    .B1(_06541_),
    .B2(_06242_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20961_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(\cs_registers_i.pc_if_i[14] ),
    .Z(_06542_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20962_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06529_),
    .A4(_06542_),
    .Z(_06543_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20963_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_06543_),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20964_ (.A1(net1581),
    .A2(_06544_),
    .B(_06249_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20965_ (.I(\cs_registers_i.pc_if_i[16] ),
    .ZN(_06545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20966_ (.A1(net1581),
    .A2(_06259_),
    .ZN(_06546_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20967_ (.I(\cs_registers_i.pc_if_i[15] ),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _20968_ (.A1(_06547_),
    .A2(_06537_),
    .A3(_06540_),
    .Z(_06548_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20969_ (.A1(_06546_),
    .A2(_06548_),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20970_ (.A1(net1581),
    .A2(net1383),
    .B(_06549_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input133 (.I(instr_rdata_i[9]),
    .Z(net132));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20972_ (.A1(_06545_),
    .A2(net1386),
    .A3(_06548_),
    .B(net1589),
    .ZN(_06552_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20973_ (.A1(_06545_),
    .A2(_06550_),
    .B1(_06552_),
    .B2(_06546_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20974_ (.I(\cs_registers_i.pc_if_i[17] ),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20975_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_06529_),
    .A3(_06542_),
    .Z(_06554_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20976_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(_06554_),
    .Z(_06555_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _20977_ (.A1(net1581),
    .A2(net1383),
    .B1(_06555_),
    .B2(_06266_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _20978_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(\cs_registers_i.pc_if_i[17] ),
    .A3(_06554_),
    .ZN(_06557_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20979_ (.A1(net1386),
    .A2(_06557_),
    .B(net1589),
    .ZN(_06558_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20980_ (.I(_06266_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20981_ (.A1(_06553_),
    .A2(_06556_),
    .B1(_06558_),
    .B2(_06559_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20982_ (.I(\cs_registers_i.pc_if_i[18] ),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20983_ (.A1(\cs_registers_i.pc_if_i[16] ),
    .A2(\cs_registers_i.pc_if_i[17] ),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20984_ (.A1(net1589),
    .A2(_06277_),
    .Z(_06562_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20985_ (.A1(_06548_),
    .A2(_06561_),
    .B(_06562_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _20986_ (.A1(net1581),
    .A2(net1383),
    .B(_06563_),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20987_ (.A1(_06560_),
    .A2(_06561_),
    .Z(_06565_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20988_ (.A1(net1386),
    .A2(_06548_),
    .A3(_06565_),
    .B(net1589),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _20989_ (.A1(_06560_),
    .A2(_06564_),
    .B1(_06566_),
    .B2(_06562_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _20990_ (.A1(_06560_),
    .A2(_06561_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _20991_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06554_),
    .A4(_06567_),
    .Z(_06568_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _20992_ (.A1(\cs_registers_i.pc_if_i[19] ),
    .A2(_06568_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _20993_ (.A1(net1589),
    .A2(_06569_),
    .B(_06287_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20994_ (.I(\cs_registers_i.pc_if_i[20] ),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _20995_ (.A1(\cs_registers_i.pc_if_i[19] ),
    .A2(_06567_),
    .Z(_06571_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _20996_ (.I(_06571_),
    .ZN(_06572_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _20997_ (.A1(_06548_),
    .A2(_06572_),
    .Z(_06573_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _20998_ (.A1(_06570_),
    .A2(net1386),
    .A3(_06573_),
    .B(net1589),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _20999_ (.A1(_06299_),
    .A2(_06573_),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21000_ (.A1(net1581),
    .A2(net1383),
    .B(_06575_),
    .ZN(_06576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21001_ (.A1(_06299_),
    .A2(_06574_),
    .B1(_06576_),
    .B2(_06570_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21002_ (.I0(_00809_),
    .I1(_00813_),
    .S(net1384),
    .Z(_06577_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21003_ (.A1(_10012_),
    .A2(_06577_),
    .B(_09991_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21004_ (.I(\cs_registers_i.pc_if_i[21] ),
    .ZN(_06578_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21005_ (.A1(\cs_registers_i.pc_if_i[20] ),
    .A2(_06554_),
    .A3(_06571_),
    .Z(_06579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21006_ (.A1(net1581),
    .A2(_06311_),
    .Z(_06580_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21007_ (.A1(net1581),
    .A2(net1383),
    .B1(_06579_),
    .B2(_06580_),
    .ZN(_06581_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21008_ (.A1(net1410),
    .A2(net1809),
    .ZN(_06582_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21009_ (.A1(_06582_),
    .A2(_06310_),
    .Z(_06583_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input132 (.I(instr_rdata_i[8]),
    .Z(net131));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21011_ (.A1(\cs_registers_i.pc_if_i[20] ),
    .A2(\cs_registers_i.pc_if_i[21] ),
    .A3(_06571_),
    .Z(_06585_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21012_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06554_),
    .A4(_06585_),
    .Z(_06586_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21013_ (.I0(_06583_),
    .I1(_06586_),
    .S(net1589),
    .Z(_06587_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21014_ (.A1(_06578_),
    .A2(_06581_),
    .B(_06587_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21015_ (.I(\cs_registers_i.pc_if_i[22] ),
    .ZN(_06588_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input131 (.I(instr_rdata_i[7]),
    .Z(net130));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21017_ (.A1(_06570_),
    .A2(_06578_),
    .A3(_06573_),
    .Z(_06590_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21018_ (.A1(_06322_),
    .A2(_06590_),
    .ZN(_06591_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21019_ (.A1(net1581),
    .A2(net1383),
    .B(_06591_),
    .ZN(_06592_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21020_ (.A1(_06588_),
    .A2(net1386),
    .A3(_06590_),
    .B(net1589),
    .ZN(_06593_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21021_ (.A1(_06588_),
    .A2(_06592_),
    .B1(_06593_),
    .B2(_06322_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21022_ (.I(\cs_registers_i.pc_if_i[23] ),
    .ZN(_06594_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _21023_ (.A1(\cs_registers_i.pc_if_i[20] ),
    .A2(\cs_registers_i.pc_if_i[21] ),
    .A3(_06554_),
    .A4(_06571_),
    .ZN(_06595_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21024_ (.A1(net1581),
    .A2(_06331_),
    .ZN(_06596_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21025_ (.A1(_06588_),
    .A2(_06595_),
    .B(_06596_),
    .ZN(_06597_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21026_ (.A1(net1581),
    .A2(net1383),
    .B(_06597_),
    .ZN(_06598_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21027_ (.A1(\cs_registers_i.pc_if_i[22] ),
    .A2(\cs_registers_i.pc_if_i[23] ),
    .ZN(_06599_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21028_ (.A1(net1386),
    .A2(_06595_),
    .A3(_06599_),
    .B(net1589),
    .ZN(_06600_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21029_ (.A1(_06594_),
    .A2(_06598_),
    .B1(_06600_),
    .B2(_06596_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21030_ (.I(\cs_registers_i.pc_if_i[24] ),
    .ZN(_06601_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21031_ (.A1(_06590_),
    .A2(_06599_),
    .B(_06341_),
    .ZN(_06602_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21032_ (.A1(net1581),
    .A2(net1383),
    .B(_06602_),
    .ZN(_06603_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21033_ (.A1(_06601_),
    .A2(_06599_),
    .Z(_06604_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21034_ (.A1(net1386),
    .A2(_06590_),
    .A3(_06604_),
    .B(net1589),
    .ZN(_06605_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21035_ (.A1(_06601_),
    .A2(_06603_),
    .B1(_06605_),
    .B2(_06341_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21036_ (.I(\cs_registers_i.pc_if_i[25] ),
    .ZN(_06606_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21037_ (.A1(_06595_),
    .A2(_06604_),
    .B(net2276),
    .ZN(_06607_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21038_ (.A1(net1581),
    .A2(net1383),
    .B(_06607_),
    .ZN(_06608_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21039_ (.A1(_06606_),
    .A2(_06604_),
    .Z(_06609_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21040_ (.A1(net1386),
    .A2(_06595_),
    .A3(_06609_),
    .B(net1589),
    .ZN(_06610_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21041_ (.A1(_06606_),
    .A2(_06608_),
    .B1(_06610_),
    .B2(net2276),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21042_ (.I(\cs_registers_i.pc_if_i[26] ),
    .ZN(_06611_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21043_ (.A1(_06590_),
    .A2(_06609_),
    .B(_06364_),
    .ZN(_06612_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21044_ (.A1(net1581),
    .A2(net1383),
    .B(_06612_),
    .ZN(_06613_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21045_ (.A1(_06611_),
    .A2(_06609_),
    .ZN(_06614_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21046_ (.I(_06614_),
    .ZN(_06615_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21047_ (.A1(_06590_),
    .A2(_06615_),
    .Z(_06616_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21048_ (.A1(net1386),
    .A2(_06616_),
    .B(net1589),
    .ZN(_06617_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21049_ (.A1(_06611_),
    .A2(_06613_),
    .B1(_06617_),
    .B2(_06364_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21050_ (.I(\cs_registers_i.pc_if_i[27] ),
    .ZN(_06618_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21051_ (.A1(_06595_),
    .A2(_06615_),
    .Z(_06619_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21052_ (.A1(_06376_),
    .A2(_06619_),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21053_ (.A1(net1581),
    .A2(net1383),
    .B(_06620_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21054_ (.A1(_06618_),
    .A2(net1386),
    .A3(_06619_),
    .B(net1589),
    .ZN(_06622_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21055_ (.A1(_06618_),
    .A2(_06621_),
    .B1(_06622_),
    .B2(_06376_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21056_ (.I(\cs_registers_i.pc_if_i[28] ),
    .ZN(_06623_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21057_ (.A1(_06618_),
    .A2(_06616_),
    .B(net2480),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21058_ (.A1(net1581),
    .A2(net1383),
    .B(_06624_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21059_ (.A1(\cs_registers_i.pc_if_i[27] ),
    .A2(\cs_registers_i.pc_if_i[28] ),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21060_ (.A1(_06615_),
    .A2(_06626_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21061_ (.A1(net1386),
    .A2(_06590_),
    .A3(_06627_),
    .B(net1589),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21062_ (.A1(_06623_),
    .A2(_06625_),
    .B1(_06628_),
    .B2(net2480),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21063_ (.I(\cs_registers_i.pc_if_i[29] ),
    .ZN(_06629_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21064_ (.A1(_06619_),
    .A2(_06626_),
    .B(_06400_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21065_ (.A1(net1581),
    .A2(net1383),
    .B(_06630_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21066_ (.A1(_06629_),
    .A2(_06626_),
    .Z(_06632_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21067_ (.A1(net1386),
    .A2(_06619_),
    .A3(_06632_),
    .B(net1589),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21068_ (.A1(_06629_),
    .A2(_06631_),
    .B1(_06633_),
    .B2(_06400_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21069_ (.I(\cs_registers_i.pc_if_i[30] ),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21070_ (.A1(_06616_),
    .A2(_06632_),
    .B(_06412_),
    .ZN(_06635_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21071_ (.A1(net1581),
    .A2(net1383),
    .B(_06635_),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21072_ (.A1(_06634_),
    .A2(_06632_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21073_ (.A1(_06614_),
    .A2(_06637_),
    .ZN(_06638_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21074_ (.A1(net1386),
    .A2(_06590_),
    .A3(_06638_),
    .B(net1589),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21075_ (.A1(_06634_),
    .A2(_06636_),
    .B1(_06639_),
    .B2(_06412_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21076_ (.A1(_10012_),
    .A2(_10009_),
    .ZN(_06640_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21077_ (.A1(_06511_),
    .A2(_00812_),
    .A3(net1385),
    .B(net1589),
    .ZN(_06641_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21078_ (.A1(_00812_),
    .A2(_06640_),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21079_ (.A1(_10012_),
    .A2(net1384),
    .B(_06642_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21080_ (.A1(_06640_),
    .A2(_06641_),
    .B1(_06643_),
    .B2(_06511_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21081_ (.I(\cs_registers_i.pc_if_i[31] ),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21082_ (.A1(_06634_),
    .A2(_06619_),
    .A3(_06632_),
    .B(_06422_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21083_ (.A1(net1581),
    .A2(net1383),
    .B(_06645_),
    .ZN(_06646_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21084_ (.A1(\cs_registers_i.pc_if_i[31] ),
    .A2(_06637_),
    .ZN(_06647_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21085_ (.A1(net1386),
    .A2(_06619_),
    .A3(_06647_),
    .B(net1589),
    .ZN(_06648_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21086_ (.A1(_06644_),
    .A2(_06646_),
    .B1(_06648_),
    .B2(_06422_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21087_ (.A1(net1384),
    .A2(_06524_),
    .Z(_06649_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21088_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(net1589),
    .Z(_06650_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21089_ (.A1(net1384),
    .A2(_06524_),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(_10012_),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21090_ (.A1(_06649_),
    .A2(_06650_),
    .B(_06651_),
    .C(_06164_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21091_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(net1393),
    .A3(_06500_),
    .A4(_06512_),
    .Z(_06652_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21092_ (.A1(\cs_registers_i.pc_if_i[5] ),
    .A2(_06652_),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21093_ (.A1(net1589),
    .A2(_06653_),
    .B(_06169_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21094_ (.A1(\cs_registers_i.pc_if_i[4] ),
    .A2(\cs_registers_i.pc_if_i[5] ),
    .A3(_06524_),
    .ZN(_06654_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21095_ (.A1(_06429_),
    .A2(_06654_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21096_ (.A1(_10012_),
    .A2(net1384),
    .B(_06655_),
    .ZN(_06656_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21097_ (.I(\cs_registers_i.pc_if_i[6] ),
    .ZN(_06657_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21098_ (.A1(_06429_),
    .A2(net1384),
    .A3(_06513_),
    .A4(_06524_),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21099_ (.A1(_10012_),
    .A2(_06429_),
    .B1(_06656_),
    .B2(_06657_),
    .C(_06658_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21100_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06512_),
    .A4(_06513_),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21101_ (.A1(\cs_registers_i.pc_if_i[7] ),
    .A2(_06659_),
    .Z(_06660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21102_ (.I0(_06185_),
    .I1(_06660_),
    .S(net1589),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21103_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06514_),
    .A4(_06524_),
    .Z(_06661_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21104_ (.A1(\cs_registers_i.pc_if_i[8] ),
    .A2(_06661_),
    .ZN(_06662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21105_ (.A1(_10012_),
    .A2(_06435_),
    .Z(_06663_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21106_ (.A1(net1589),
    .A2(_06662_),
    .B(_06663_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21107_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06512_),
    .A4(_06515_),
    .Z(_06664_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21108_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_06664_),
    .Z(_06665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21109_ (.I0(_06159_),
    .I1(_06665_),
    .S(net1589),
    .Z(_03009_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21110_ (.A1(net1393),
    .A2(_06500_),
    .A3(_06516_),
    .A4(_06524_),
    .Z(_06666_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _21111_ (.A1(\cs_registers_i.pc_if_i[10] ),
    .A2(_06666_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21112_ (.I(_06151_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21113_ (.A1(net1589),
    .A2(_06667_),
    .B(_06668_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21114_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21115_ (.A1(_06450_),
    .A2(net1393),
    .A3(_06457_),
    .Z(_06670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21116_ (.I0(_06469_),
    .I1(_06670_),
    .S(_10023_),
    .Z(_06671_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input130 (.I(instr_rdata_i[6]),
    .Z(net129));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input129 (.I(instr_rdata_i[5]),
    .Z(net128));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21119_ (.I(net101),
    .ZN(_06674_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21120_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21121_ (.I0(_06674_),
    .I1(_06675_),
    .S(net2024),
    .Z(_06676_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21122_ (.A1(net1393),
    .A2(_06457_),
    .B(_10023_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21123_ (.A1(_10023_),
    .A2(net1393),
    .A3(_06457_),
    .Z(_06678_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21124_ (.A1(net1393),
    .A2(net1501),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _21125_ (.A1(net1819),
    .A2(_06677_),
    .A3(_06678_),
    .B(_06679_),
    .ZN(_06680_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input128 (.I(instr_rdata_i[4]),
    .Z(net127));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input127 (.I(instr_rdata_i[3]),
    .Z(net126));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21128_ (.A1(_06669_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06683_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21129_ (.A1(_06669_),
    .A2(_06671_),
    .B1(_06676_),
    .B2(_06680_),
    .C(_06683_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21130_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .ZN(_06684_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input126 (.I(instr_rdata_i[31]),
    .Z(net125));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21132_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(net2024),
    .Z(_06686_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21133_ (.I(_06686_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21134_ (.A1(_06684_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06688_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21135_ (.A1(_06684_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06687_),
    .C(_06688_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21136_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21137_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(net2024),
    .Z(_06690_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21138_ (.I(_06690_),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21139_ (.A1(_06689_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06692_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21140_ (.A1(_06689_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06691_),
    .C(_06692_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21141_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21142_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(net2024),
    .Z(_06694_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21143_ (.I(_06694_),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21144_ (.A1(_06693_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06696_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21145_ (.A1(_06693_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06695_),
    .C(_06696_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21146_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21147_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(net2024),
    .Z(_06698_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21148_ (.I(_06698_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input125 (.I(instr_rdata_i[30]),
    .Z(net124));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21150_ (.A1(_06697_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06701_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21151_ (.A1(_06697_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06699_),
    .C(_06701_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21152_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21153_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(net2024),
    .Z(_06703_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21154_ (.I(_06703_),
    .ZN(_06704_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input124 (.I(instr_rdata_i[2]),
    .Z(net123));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21156_ (.A1(_06702_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06706_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21157_ (.A1(_06702_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06704_),
    .C(_06706_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21158_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21159_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(net2024),
    .Z(_06708_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21160_ (.I(_06708_),
    .ZN(_06709_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21161_ (.A1(_06707_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06710_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21162_ (.A1(_06707_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06709_),
    .C(_06710_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21163_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21164_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21165_ (.I0(_06711_),
    .I1(_06712_),
    .S(_06467_),
    .Z(_06713_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21166_ (.A1(_10023_),
    .A2(net2024),
    .A3(_06712_),
    .A4(_06444_),
    .Z(_06714_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21167_ (.I(net108),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21168_ (.A1(_10023_),
    .A2(_06715_),
    .A3(_06450_),
    .A4(_06444_),
    .Z(_06716_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21169_ (.A1(net2025),
    .A2(_06715_),
    .A3(_06450_),
    .A4(_06444_),
    .Z(_06717_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input123 (.I(instr_rdata_i[29]),
    .Z(net122));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21171_ (.I0(_06716_),
    .I1(_06717_),
    .S(net1387),
    .Z(_06719_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21172_ (.A1(_06460_),
    .A2(_06713_),
    .B(_06714_),
    .C(_06719_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input122 (.I(instr_rdata_i[28]),
    .Z(net121));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input121 (.I(instr_rdata_i[27]),
    .Z(net120));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21175_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06722_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21176_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .A2(net1382),
    .B(_06722_),
    .ZN(_06723_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input120 (.I(instr_rdata_i[26]),
    .Z(net119));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input119 (.I(instr_rdata_i[25]),
    .Z(net118));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21179_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06726_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input118 (.I(instr_rdata_i[24]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21181_ (.A1(net2025),
    .A2(net109),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input117 (.I(instr_rdata_i[23]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input116 (.I(instr_rdata_i[22]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21184_ (.A1(_10023_),
    .A2(net109),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21185_ (.I0(_06728_),
    .I1(_06731_),
    .S(net1387),
    .Z(_06732_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21186_ (.A1(_06460_),
    .A2(_06723_),
    .B(_06726_),
    .C(_06732_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21187_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06733_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21188_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .A2(net1382),
    .B(_06733_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21189_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06735_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21190_ (.A1(net2025),
    .A2(net110),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21191_ (.A1(_10023_),
    .A2(net110),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06737_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21192_ (.I0(_06736_),
    .I1(_06737_),
    .S(net1387),
    .Z(_06738_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21193_ (.A1(_06460_),
    .A2(_06734_),
    .B(_06735_),
    .C(_06738_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21194_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06739_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21195_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .A2(net1382),
    .B(_06739_),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21196_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21197_ (.A1(net2025),
    .A2(net111),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06742_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input115 (.I(instr_rdata_i[21]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21199_ (.A1(_10023_),
    .A2(net111),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06744_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21200_ (.I0(_06742_),
    .I1(_06744_),
    .S(net1387),
    .Z(_06745_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21201_ (.A1(_06460_),
    .A2(_06740_),
    .B(_06741_),
    .C(_06745_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21202_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21203_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(net2024),
    .Z(_06747_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21204_ (.I(_06747_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21205_ (.A1(_06746_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06749_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21206_ (.A1(_06746_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06748_),
    .C(_06749_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21207_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21208_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .A2(net1382),
    .B(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21209_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input114 (.I(instr_rdata_i[20]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21211_ (.A1(net2025),
    .A2(net113),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21212_ (.A1(_10023_),
    .A2(net113),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21213_ (.I0(_06754_),
    .I1(_06755_),
    .S(net1387),
    .Z(_06756_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21214_ (.A1(_06460_),
    .A2(_06751_),
    .B(_06752_),
    .C(_06756_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21215_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06757_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21216_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .A2(net1382),
    .B(_06757_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21217_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21218_ (.A1(net2025),
    .A2(net114),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21219_ (.A1(_10023_),
    .A2(net114),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21220_ (.I0(_06760_),
    .I1(_06761_),
    .S(net1387),
    .Z(_06762_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21221_ (.A1(_06460_),
    .A2(_06758_),
    .B(_06759_),
    .C(_06762_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21222_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06763_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21223_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .A2(net1382),
    .B(_06763_),
    .ZN(_06764_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21224_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21225_ (.A1(net2025),
    .A2(net115),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21226_ (.A1(_10023_),
    .A2(net115),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06767_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21227_ (.I0(_06766_),
    .I1(_06767_),
    .S(net1387),
    .Z(_06768_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21228_ (.A1(_06460_),
    .A2(_06764_),
    .B(_06765_),
    .C(_06768_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21229_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06769_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21230_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .A2(net1382),
    .B(_06769_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21231_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06771_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21232_ (.A1(net2025),
    .A2(net116),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21233_ (.A1(_10023_),
    .A2(net116),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06773_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21234_ (.I0(_06772_),
    .I1(_06773_),
    .S(net1387),
    .Z(_06774_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21235_ (.A1(_06460_),
    .A2(_06770_),
    .B(_06771_),
    .C(_06774_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21236_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06775_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21237_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .A2(net1382),
    .B(_06775_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21238_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21239_ (.A1(net2025),
    .A2(net117),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21240_ (.A1(_10023_),
    .A2(net117),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21241_ (.I0(_06778_),
    .I1(_06779_),
    .S(net1387),
    .Z(_06780_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21242_ (.A1(_06460_),
    .A2(_06776_),
    .B(_06777_),
    .C(_06780_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21243_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06781_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21244_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .A2(net1382),
    .B(_06781_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21245_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06783_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21246_ (.A1(net2025),
    .A2(net118),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06784_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21247_ (.A1(_10023_),
    .A2(net118),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06785_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21248_ (.I0(_06784_),
    .I1(_06785_),
    .S(net1387),
    .Z(_06786_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21249_ (.A1(_06460_),
    .A2(_06782_),
    .B(_06783_),
    .C(_06786_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21250_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06787_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21251_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .A2(net1382),
    .B(_06787_),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21252_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06789_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21253_ (.A1(net2025),
    .A2(net119),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06790_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21254_ (.A1(_10023_),
    .A2(net119),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06791_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21255_ (.I0(_06790_),
    .I1(_06791_),
    .S(net1387),
    .Z(_06792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21256_ (.A1(_06460_),
    .A2(_06788_),
    .B(_06789_),
    .C(_06792_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21257_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06793_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21258_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .A2(net1382),
    .B(_06793_),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21259_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21260_ (.A1(net2025),
    .A2(net120),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21261_ (.A1(_10023_),
    .A2(net120),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21262_ (.I0(_06796_),
    .I1(_06797_),
    .S(net1387),
    .Z(_06798_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21263_ (.A1(_06460_),
    .A2(_06794_),
    .B(_06795_),
    .C(_06798_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21264_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06799_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21265_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .A2(net1382),
    .B(_06799_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21266_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06801_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21267_ (.A1(net2025),
    .A2(net121),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21268_ (.A1(_10023_),
    .A2(net121),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21269_ (.I0(_06802_),
    .I1(_06803_),
    .S(net1387),
    .Z(_06804_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21270_ (.A1(_06460_),
    .A2(_06800_),
    .B(_06801_),
    .C(_06804_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21271_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06805_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21272_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .A2(net1382),
    .B(_06805_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21273_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06807_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21274_ (.A1(net2025),
    .A2(net122),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21275_ (.A1(_10023_),
    .A2(net122),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21276_ (.I0(_06808_),
    .I1(_06809_),
    .S(net1387),
    .Z(_06810_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21277_ (.A1(_06460_),
    .A2(_06806_),
    .B(_06807_),
    .C(_06810_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21278_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .ZN(_06811_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21279_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(net2024),
    .Z(_06812_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21280_ (.I(_06812_),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21281_ (.A1(_06811_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06814_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21282_ (.A1(_06811_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06813_),
    .C(_06814_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21283_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21284_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .A2(net1382),
    .B(_06815_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21285_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21286_ (.A1(net2025),
    .A2(net124),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06818_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21287_ (.A1(_10023_),
    .A2(net124),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21288_ (.I0(_06818_),
    .I1(_06819_),
    .S(net1387),
    .Z(_06820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21289_ (.A1(_06460_),
    .A2(_06816_),
    .B(_06817_),
    .C(_06820_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21290_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .A2(net1394),
    .A3(net1501),
    .Z(_06821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21291_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .A2(net1382),
    .B(_06821_),
    .ZN(_06822_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21292_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .A2(net1819),
    .A3(_06476_),
    .ZN(_06823_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21293_ (.A1(net2025),
    .A2(net125),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21294_ (.A1(_10023_),
    .A2(net125),
    .A3(net2024),
    .A4(net1819),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21295_ (.I0(_06824_),
    .I1(_06825_),
    .S(net1387),
    .Z(_06826_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21296_ (.A1(_06460_),
    .A2(_06822_),
    .B(_06823_),
    .C(_06826_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21297_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(net2023),
    .Z(_06827_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21298_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .I1(_06827_),
    .S(net1378),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21299_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(net2023),
    .Z(_06828_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21300_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .I1(_06828_),
    .S(net1378),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21301_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(net2023),
    .Z(_06829_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21302_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .I1(_06829_),
    .S(net1378),
    .Z(_03038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21303_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(net2023),
    .Z(_06830_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21304_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .I1(_06830_),
    .S(net1378),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21305_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(net2023),
    .Z(_06831_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21306_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .I1(_06831_),
    .S(net1378),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21307_ (.I0(net128),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(net2023),
    .Z(_06832_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21308_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .I1(_06832_),
    .S(net1378),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21309_ (.I0(net129),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(net2023),
    .Z(_06833_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21310_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .I1(_06833_),
    .S(net1378),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21311_ (.I0(net130),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(net2023),
    .Z(_06834_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21312_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .I1(_06834_),
    .S(net1378),
    .Z(_03043_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21313_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .ZN(_06835_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21314_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(net2024),
    .Z(_06836_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21315_ (.I(_06836_),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21316_ (.A1(_06835_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06838_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21317_ (.A1(_06835_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06837_),
    .C(_06838_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input113 (.I(instr_rdata_i[1]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21319_ (.I0(net131),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(net2023),
    .Z(_06840_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21320_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .I1(_06840_),
    .S(net1378),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21321_ (.I0(net132),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(net2023),
    .Z(_06841_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input112 (.I(instr_rdata_i[19]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21323_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .I1(_06841_),
    .S(net1378),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21324_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(net2023),
    .Z(_06843_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21325_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .I1(_06843_),
    .S(net1378),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21326_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(net2023),
    .Z(_06844_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21327_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .I1(_06844_),
    .S(net1378),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21328_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(net2023),
    .Z(_06845_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21329_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .I1(_06845_),
    .S(net1378),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21330_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(net2023),
    .Z(_06846_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21331_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .I1(_06846_),
    .S(net1378),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21332_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(net2023),
    .Z(_06847_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21333_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .I1(_06847_),
    .S(net1378),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21334_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(net2023),
    .Z(_06848_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21335_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .I1(_06848_),
    .S(net1378),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21336_ (.I0(net108),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(net2023),
    .Z(_06849_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21337_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .I1(_06849_),
    .S(net1378),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21338_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(net2023),
    .Z(_06850_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21339_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .I1(_06850_),
    .S(net1378),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21340_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21341_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(net2024),
    .Z(_06852_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21342_ (.I(_06852_),
    .ZN(_06853_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21343_ (.A1(_06851_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06854_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21344_ (.A1(_06851_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06853_),
    .C(_06854_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input111 (.I(instr_rdata_i[18]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21346_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(net2023),
    .Z(_06856_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21347_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .I1(_06856_),
    .S(net1378),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21348_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(net2023),
    .Z(_06857_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input110 (.I(instr_rdata_i[17]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21350_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .I1(_06857_),
    .S(net1378),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21351_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(net2023),
    .Z(_06859_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21352_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .I1(_06859_),
    .S(net1378),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21353_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(net2023),
    .Z(_06860_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21354_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .I1(_06860_),
    .S(net1378),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21355_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(net2023),
    .Z(_06861_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21356_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .I1(_06861_),
    .S(net1378),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21357_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(net2023),
    .Z(_06862_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21358_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .I1(_06862_),
    .S(net1378),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21359_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(net2023),
    .Z(_06863_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21360_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .I1(_06863_),
    .S(net1378),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21361_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(net2023),
    .Z(_06864_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21362_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .I1(_06864_),
    .S(net1378),
    .Z(_03063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21363_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(net2023),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21364_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .I1(_06865_),
    .S(net1378),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21365_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(net2023),
    .Z(_06866_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21366_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .I1(_06866_),
    .S(net1378),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21367_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21368_ (.I0(net128),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(net2024),
    .Z(_06868_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21369_ (.I(_06868_),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21370_ (.A1(_06867_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21371_ (.A1(_06867_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06869_),
    .C(_06870_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21372_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(net2023),
    .Z(_06871_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21373_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .I1(_06871_),
    .S(net1378),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21374_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(net2023),
    .Z(_06872_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21375_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .I1(_06872_),
    .S(net1378),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21376_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(net2023),
    .Z(_06873_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21377_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .I1(_06873_),
    .S(net1378),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21378_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(net2023),
    .Z(_06874_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21379_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .I1(_06874_),
    .S(net1378),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21380_ (.I0(net101),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(net1805),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21381_ (.I0(net112),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(net1805),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21382_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(net1805),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21383_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(net1805),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21384_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(net1805),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21385_ (.I0(net128),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(net1805),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21386_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21387_ (.I0(net129),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(net2024),
    .Z(_06876_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21388_ (.I(_06876_),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21389_ (.A1(_06875_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21390_ (.A1(_06875_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06877_),
    .C(_06878_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21391_ (.I0(net129),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(net1805),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21392_ (.I0(net130),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(net1805),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21393_ (.I0(net131),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(net1805),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(instr_rdata_i[16]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21395_ (.I0(net132),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(net1805),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21396_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(net1805),
    .Z(_03082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21397_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(net1805),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21398_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(net1805),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21399_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(net1805),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21400_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(net1805),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21401_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(net1805),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21402_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21403_ (.I0(net130),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(net2024),
    .Z(_06881_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21404_ (.I(_06881_),
    .ZN(_06882_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21405_ (.A1(_06880_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06883_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21406_ (.A1(_06880_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06882_),
    .C(_06883_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21407_ (.I0(net108),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(net1805),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21408_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(net1805),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21409_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(net1805),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(instr_rdata_i[15]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21411_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(net1805),
    .Z(_03092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21412_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(net1805),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21413_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(net1805),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21414_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(net1805),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21415_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(net1805),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21416_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(net1805),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21417_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(net1805),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21418_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21419_ (.I0(net131),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(net2024),
    .Z(_06886_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21420_ (.I(_06886_),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21421_ (.A1(_06885_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06888_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21422_ (.A1(_06885_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06887_),
    .C(_06888_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21423_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(net1805),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21424_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(net1805),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21425_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(net1805),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21426_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(net1805),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21427_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(net1805),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21428_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(net1805),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21429_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21430_ (.I0(net132),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(net2024),
    .Z(_06890_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21431_ (.I(_06890_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21432_ (.A1(_06889_),
    .A2(net1819),
    .A3(_06679_),
    .Z(_06892_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21433_ (.A1(_06889_),
    .A2(_06671_),
    .B1(_06680_),
    .B2(_06891_),
    .C(_06892_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21434_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .I1(_06153_),
    .S(net1834),
    .Z(net224));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21435_ (.A1(net100),
    .A2(_10081_),
    .Z(_06893_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(instr_rdata_i[14]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21437_ (.I0(net224),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .S(_06893_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21438_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .I1(_06203_),
    .S(net1834),
    .Z(net225));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21439_ (.I0(net225),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .S(_06893_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21440_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .I1(_06215_),
    .S(net1834),
    .Z(net226));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21441_ (.I0(net226),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .S(_06893_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21442_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .I1(_06226_),
    .S(net1834),
    .Z(net227));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21443_ (.I0(net227),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .S(_06893_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21444_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .I1(_06251_),
    .S(net1834),
    .Z(net228));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21445_ (.I0(net228),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .S(_06893_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21446_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .I1(_06250_),
    .S(net1834),
    .Z(net229));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21447_ (.I0(net229),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .S(_06893_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21448_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .I1(_06260_),
    .S(net1834),
    .Z(net230));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21449_ (.I0(net230),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .S(_06893_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(instr_rdata_i[13]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21451_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .I1(_06268_),
    .S(net1834),
    .Z(net231));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21452_ (.I0(net231),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .S(_06893_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21453_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .I1(_06279_),
    .S(net1834),
    .Z(net232));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21454_ (.I0(net232),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .S(_06893_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21455_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .I1(_06288_),
    .S(net1834),
    .Z(net233));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21456_ (.I0(net233),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .S(_06893_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21457_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .I1(_06380_),
    .S(net1834),
    .Z(net234));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(instr_rdata_i[12]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21459_ (.I0(net234),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .S(_06893_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21460_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .I1(_06312_),
    .S(net1834),
    .Z(net235));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21461_ (.I0(net235),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .S(net1541),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21462_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .I1(_06333_),
    .S(net1834),
    .Z(net236));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21463_ (.I0(net236),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .S(_06893_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21464_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .I1(_06332_),
    .S(net1834),
    .Z(net237));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21465_ (.I0(net237),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .S(_06893_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21466_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .I1(_06354_),
    .S(net1834),
    .Z(net238));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21467_ (.I0(net238),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .S(_06893_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21468_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .I1(_06367_),
    .S(net1834),
    .Z(net239));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21469_ (.I0(net239),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .S(_06893_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21470_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .I1(_06366_),
    .S(net1834),
    .Z(net240));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21471_ (.I0(net240),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .S(_06893_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(instr_rdata_i[11]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21473_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .I1(_06377_),
    .S(net1834),
    .Z(net241));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21474_ (.I0(net241),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .S(_06893_),
    .Z(_03124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21475_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .I1(_06393_),
    .S(net1834),
    .Z(net242));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21476_ (.I0(net242),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .S(_06893_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21477_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .I1(_06402_),
    .S(net1834),
    .Z(net243));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21478_ (.I0(net243),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .S(_06893_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21479_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .I1(_01372_),
    .S(net1834),
    .Z(net244));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input103 (.I(instr_rdata_i[10]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21481_ (.I0(net244),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .S(net1541),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21482_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .I1(_06414_),
    .S(net1834),
    .Z(net245));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21483_ (.I0(net245),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .S(_06893_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21484_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .I1(_06424_),
    .S(net1834),
    .Z(net246));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21485_ (.I0(net246),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .S(_06893_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21486_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .I1(_01374_),
    .S(net1834),
    .Z(net247));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21487_ (.I0(net247),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .S(net1541),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21488_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .I1(_06165_),
    .S(net1834),
    .Z(net248));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21489_ (.I0(net248),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .S(net1541),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21490_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .I1(_06170_),
    .S(net1834),
    .Z(net249));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21491_ (.I0(net249),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .S(net1541),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21492_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .I1(_06431_),
    .S(net1834),
    .Z(net250));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21493_ (.I0(net250),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .S(net1541),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21494_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .I1(_06186_),
    .S(net1834),
    .Z(net251));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21495_ (.I0(net251),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .S(_06893_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21496_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .ZN(_06899_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21497_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_06440_),
    .A3(_06663_),
    .B(_06899_),
    .ZN(net252));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21498_ (.I0(net252),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .S(_06893_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21499_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .I1(_06160_),
    .S(net1834),
    .Z(net253));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21500_ (.I0(net253),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .S(net1541),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21501_ (.A1(net64),
    .A2(_09655_),
    .Z(_06900_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21502_ (.I0(_10129_),
    .I1(_06900_),
    .S(net2087),
    .Z(_06901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21503_ (.A1(net2086),
    .A2(\load_store_unit_i.lsu_err_q ),
    .ZN(_06902_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21504_ (.I0(_06901_),
    .I1(_06902_),
    .S(net2098),
    .Z(_06903_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21505_ (.A1(net31),
    .A2(_06903_),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21506_ (.A1(_07550_),
    .A2(_06900_),
    .Z(_06905_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21507_ (.I0(_06904_),
    .I1(_06905_),
    .S(net2081),
    .Z(_06906_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input102 (.I(instr_rdata_i[0]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input101 (.I(instr_gnt_i),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21510_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .I1(\alu_adder_result_ex[0] ),
    .S(net1513),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21511_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .I1(net1451),
    .S(net1513),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21512_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .I1(net1457),
    .S(net1513),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21513_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .I1(net2298),
    .S(net1513),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21514_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .I1(net1450),
    .S(net1513),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21515_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .I1(net2292),
    .S(net1513),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21516_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .I1(net1448),
    .S(net1513),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21517_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .I1(net1446),
    .S(net1513),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21518_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .I1(net2288),
    .S(net1513),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21519_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .I1(net1435),
    .S(net1513),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input100 (.I(instr_err_i),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21521_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .I1(net1436),
    .S(net1513),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21522_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .I1(net1539),
    .S(net1513),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21523_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .I1(net2278),
    .S(net1513),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21524_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .I1(net1410),
    .S(net1513),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21525_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .I1(net1432),
    .S(net1513),
    .Z(_03234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21526_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .I1(net169),
    .S(net1513),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21527_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .I1(net2204),
    .S(net1513),
    .Z(_03236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21528_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .I1(net1431),
    .S(net1513),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21529_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .I1(net1409),
    .S(net1513),
    .Z(_03238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21530_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .I1(net1429),
    .S(net1513),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input99 (.I(hart_id_i[9]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21532_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .I1(net2138),
    .S(net1513),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21533_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .I1(net2169),
    .S(net1513),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21534_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .I1(net176),
    .S(net1513),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21535_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .I1(net2122),
    .S(net1513),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21536_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .I1(net2051),
    .S(net1513),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21537_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .I1(net1519),
    .S(net1513),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21538_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .I1(net1454),
    .S(net1513),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21539_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .I1(net1499),
    .S(net1513),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21540_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .I1(net1500),
    .S(net1513),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21541_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .I1(net1512),
    .S(net1513),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21542_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .I1(net1458),
    .S(net1513),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21543_ (.I0(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .I1(net1459),
    .S(net1513),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21544_ (.A1(_07557_),
    .A2(_07579_),
    .A3(net2149),
    .A4(_07711_),
    .Z(_06911_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21545_ (.I0(_06911_),
    .I1(\load_store_unit_i.data_sign_ext_q ),
    .S(_10132_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21546_ (.A1(_07616_),
    .A2(_10124_),
    .A3(_09538_),
    .Z(net223));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21547_ (.I0(net223),
    .I1(\load_store_unit_i.data_we_q ),
    .S(_10132_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input98 (.I(hart_id_i[8]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21549_ (.A1(net2022),
    .A2(_01360_),
    .Z(_06913_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21550_ (.A1(_08000_),
    .A2(_10125_),
    .ZN(_06914_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21551_ (.I0(_06913_),
    .I1(net1520),
    .S(_06914_),
    .Z(_06915_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21552_ (.A1(net2098),
    .A2(_06915_),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21553_ (.I(net31),
    .ZN(_06917_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21554_ (.A1(_07552_),
    .A2(net64),
    .Z(_06918_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21555_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_06917_),
    .A3(_06918_),
    .ZN(_06919_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21556_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_06916_),
    .B(_06919_),
    .ZN(_06920_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21557_ (.A1(net2098),
    .A2(_10129_),
    .B(net31),
    .ZN(_06921_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21558_ (.A1(net31),
    .A2(_06918_),
    .B(net2087),
    .ZN(_06922_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21559_ (.A1(_06921_),
    .A2(_06922_),
    .B(net2081),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21560_ (.I0(\load_store_unit_i.handle_misaligned_q ),
    .I1(_06920_),
    .S(_06923_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21561_ (.I0(net64),
    .I1(_10129_),
    .S(_07652_),
    .Z(_06924_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21562_ (.A1(net2098),
    .A2(_06924_),
    .Z(_06925_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21563_ (.A1(_07553_),
    .A2(_06917_),
    .A3(_06925_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21564_ (.A1(_10129_),
    .A2(_06916_),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .ZN(_06926_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21565_ (.A1(net31),
    .A2(_06926_),
    .Z(_06927_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21566_ (.A1(_10129_),
    .A2(_06915_),
    .B(net2098),
    .ZN(_06928_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21567_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_06917_),
    .A3(_06928_),
    .Z(_06929_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21568_ (.A1(_06927_),
    .A2(_06929_),
    .B(net2081),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21569_ (.I0(_07553_),
    .I1(_10131_),
    .S(net2087),
    .Z(_06930_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21570_ (.A1(net2098),
    .A2(net64),
    .A3(_06930_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21571_ (.A1(_07652_),
    .A2(net64),
    .Z(_06931_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21572_ (.I0(_06924_),
    .I1(_06931_),
    .S(net2081),
    .Z(_06932_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21573_ (.A1(_07552_),
    .A2(_06932_),
    .Z(_06933_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _21574_ (.A1(net2081),
    .A2(net2086),
    .Z(_06934_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21575_ (.A1(_06918_),
    .A2(_06934_),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21576_ (.A1(_09656_),
    .A2(_06933_),
    .B1(_06935_),
    .B2(_09655_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21577_ (.I0(\alu_adder_result_ex[0] ),
    .I1(net1887),
    .S(_10132_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21578_ (.I0(net1539),
    .I1(net1886),
    .S(_10132_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21579_ (.A1(\load_store_unit_i.data_we_q ),
    .A2(_06935_),
    .Z(_06936_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input97 (.I(hart_id_i[7]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21581_ (.I0(net62),
    .I1(\load_store_unit_i.rdata_q[0] ),
    .S(net1745),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21582_ (.I0(net41),
    .I1(\load_store_unit_i.rdata_q[10] ),
    .S(net1745),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21583_ (.I0(net42),
    .I1(\load_store_unit_i.rdata_q[11] ),
    .S(net1745),
    .Z(_03263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21584_ (.I0(net44),
    .I1(\load_store_unit_i.rdata_q[12] ),
    .S(net1745),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21585_ (.I0(net45),
    .I1(\load_store_unit_i.rdata_q[13] ),
    .S(net1745),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21586_ (.I0(net46),
    .I1(\load_store_unit_i.rdata_q[14] ),
    .S(net1745),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21587_ (.I0(net47),
    .I1(\load_store_unit_i.rdata_q[15] ),
    .S(net1745),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21588_ (.I0(net48),
    .I1(\load_store_unit_i.rdata_q[16] ),
    .S(net1745),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21589_ (.I0(net49),
    .I1(\load_store_unit_i.rdata_q[17] ),
    .S(net1745),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21590_ (.I0(net50),
    .I1(\load_store_unit_i.rdata_q[18] ),
    .S(net1745),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input96 (.I(hart_id_i[6]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21592_ (.I0(net51),
    .I1(\load_store_unit_i.rdata_q[19] ),
    .S(net1745),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21593_ (.I0(net63),
    .I1(\load_store_unit_i.rdata_q[1] ),
    .S(net1745),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21594_ (.I0(net52),
    .I1(\load_store_unit_i.rdata_q[20] ),
    .S(net1745),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21595_ (.I0(net53),
    .I1(\load_store_unit_i.rdata_q[21] ),
    .S(net1745),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21596_ (.I0(net55),
    .I1(\load_store_unit_i.rdata_q[22] ),
    .S(net1745),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21597_ (.I0(net56),
    .I1(\load_store_unit_i.rdata_q[23] ),
    .S(net1745),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21598_ (.I0(net33),
    .I1(\load_store_unit_i.rdata_q[2] ),
    .S(net1745),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21599_ (.I0(net34),
    .I1(\load_store_unit_i.rdata_q[3] ),
    .S(net1745),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21600_ (.I0(net35),
    .I1(\load_store_unit_i.rdata_q[4] ),
    .S(net1745),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21601_ (.I0(net36),
    .I1(\load_store_unit_i.rdata_q[5] ),
    .S(net1745),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21602_ (.I0(net37),
    .I1(\load_store_unit_i.rdata_q[6] ),
    .S(net1745),
    .Z(_03281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21603_ (.I0(net38),
    .I1(\load_store_unit_i.rdata_q[7] ),
    .S(net1745),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21604_ (.I0(net39),
    .I1(\load_store_unit_i.rdata_q[8] ),
    .S(net1745),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21605_ (.I0(net40),
    .I1(\load_store_unit_i.rdata_q[9] ),
    .S(net1745),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21606_ (.A1(\cs_registers_i.priv_mode_id_o[0] ),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_q[0] ),
    .ZN(_06939_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21607_ (.A1(net1746),
    .A2(net1588),
    .ZN(_06940_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _21608_ (.A1(_07773_),
    .A2(net1702),
    .A3(_09635_),
    .A4(_09568_),
    .ZN(_06941_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21609_ (.A1(_10371_),
    .A2(_10193_),
    .A3(_06941_),
    .Z(_06942_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21610_ (.A1(_06940_),
    .A2(_06942_),
    .Z(_06943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21611_ (.A1(_03471_),
    .A2(_10404_),
    .B(net1588),
    .C(net1746),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21612_ (.A1(_06943_),
    .A2(_06944_),
    .Z(_06945_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21613_ (.A1(\cs_registers_i.mstatus_q[2] ),
    .A2(_04146_),
    .B(_06945_),
    .ZN(_06946_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21614_ (.A1(_06939_),
    .A2(_06946_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21615_ (.A1(\cs_registers_i.priv_mode_id_o[1] ),
    .A2(net1588),
    .B1(net1707),
    .B2(\cs_registers_i.mstack_q[1] ),
    .ZN(_06947_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21616_ (.A1(_04146_),
    .A2(_06944_),
    .Z(_06948_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21617_ (.A1(\cs_registers_i.mstatus_q[3] ),
    .A2(_06948_),
    .B(_06945_),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21618_ (.A1(_06947_),
    .A2(_06949_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21619_ (.A1(_09939_),
    .A2(\cs_registers_i.mstack_q[2] ),
    .Z(_06950_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21620_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(net1588),
    .B1(_06950_),
    .B2(net1746),
    .C(_06943_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21621_ (.I(_04146_),
    .ZN(_06952_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21622_ (.A1(_10984_),
    .A2(_06952_),
    .B(_06940_),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21623_ (.I(\cs_registers_i.mstatus_q[4] ),
    .ZN(_06954_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21624_ (.A1(_06954_),
    .A2(_06952_),
    .A3(_06940_),
    .Z(_06955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21625_ (.A1(_06951_),
    .A2(_06953_),
    .B(_06955_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21626_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_06943_),
    .Z(_06956_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21627_ (.A1(\cs_registers_i.mstatus_q[4] ),
    .A2(net1746),
    .Z(_06957_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21628_ (.A1(_10891_),
    .A2(_04015_),
    .A3(_04146_),
    .Z(_06958_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21629_ (.A1(_06956_),
    .A2(_06957_),
    .A3(_06958_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21630_ (.I(\cs_registers_i.pc_if_i[1] ),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input95 (.I(hart_id_i[5]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21632_ (.I0(_06674_),
    .I1(_06669_),
    .S(net2025),
    .Z(_06961_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21633_ (.I0(_06715_),
    .I1(_06711_),
    .S(net2025),
    .Z(_06962_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21634_ (.A1(net2026),
    .A2(_06962_),
    .Z(_06963_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21635_ (.A1(_06959_),
    .A2(_06961_),
    .B(_06963_),
    .ZN(_06964_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input94 (.I(hart_id_i[4]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21637_ (.A1(net2025),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B(_10024_),
    .ZN(_06966_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21638_ (.I0(net109),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(net2025),
    .Z(_06967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21639_ (.A1(net2026),
    .A2(_06967_),
    .ZN(_06968_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21640_ (.A1(net2026),
    .A2(_06966_),
    .B(_06968_),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input93 (.I(hart_id_i[3]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21642_ (.I0(net125),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(net2025),
    .Z(_06971_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21643_ (.I0(net107),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .S(net2025),
    .Z(_06972_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21644_ (.I0(_06971_),
    .I1(_06972_),
    .S(_06959_),
    .Z(_06973_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input92 (.I(hart_id_i[31]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input91 (.I(hart_id_i[30]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21647_ (.I0(net121),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(net2025),
    .Z(_06976_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21648_ (.I0(net104),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .S(net2025),
    .Z(_06977_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21649_ (.A1(_06959_),
    .A2(_06977_),
    .Z(_06978_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21650_ (.A1(net2026),
    .A2(_06976_),
    .B(_06978_),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21651_ (.I0(net131),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .S(net2025),
    .Z(_06980_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21652_ (.I0(net117),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(net2025),
    .Z(_06981_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21653_ (.I0(_06980_),
    .I1(_06981_),
    .S(net2026),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input90 (.I(hart_id_i[2]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21655_ (.I0(net132),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .S(net2025),
    .Z(_06984_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21656_ (.I0(net118),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(net2025),
    .Z(_06985_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21657_ (.I0(_06984_),
    .I1(_06985_),
    .S(net2026),
    .Z(_06986_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input89 (.I(hart_id_i[29]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21659_ (.I0(net130),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .S(net2025),
    .Z(_06988_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21660_ (.I0(net116),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(net2025),
    .Z(_06989_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21661_ (.I0(_06988_),
    .I1(_06989_),
    .S(net2026),
    .Z(_06990_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21662_ (.I0(net119),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(net2025),
    .Z(_06991_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21663_ (.I0(net102),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .S(net2025),
    .Z(_06992_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21664_ (.I0(_06991_),
    .I1(_06992_),
    .S(_06959_),
    .Z(_06993_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21665_ (.I0(net120),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(net2025),
    .Z(_06994_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21666_ (.I0(net103),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .S(net2025),
    .Z(_06995_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21667_ (.I0(_06994_),
    .I1(_06995_),
    .S(_06959_),
    .Z(_06996_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21668_ (.A1(_06993_),
    .A2(_06996_),
    .Z(_06997_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21669_ (.A1(_06982_),
    .A2(_06986_),
    .A3(_06990_),
    .A4(_06997_),
    .Z(_06998_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21670_ (.I0(net124),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(net2025),
    .Z(_06999_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21671_ (.I0(net106),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .S(net2025),
    .Z(_07000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21672_ (.I0(_06999_),
    .I1(_07000_),
    .S(_06959_),
    .Z(_07001_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input88 (.I(hart_id_i[28]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21674_ (.I0(_06979_),
    .I1(_06998_),
    .S(_07001_),
    .Z(_07003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21675_ (.I0(_06976_),
    .I1(_06977_),
    .S(_06959_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input87 (.I(hart_id_i[27]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input86 (.I(hart_id_i[26]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21678_ (.A1(_06959_),
    .A2(_06972_),
    .Z(_07007_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21679_ (.A1(net2026),
    .A2(_06971_),
    .B(_07007_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input85 (.I(hart_id_i[25]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21681_ (.I0(net111),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(net2025),
    .Z(_07010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21682_ (.I0(net126),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .S(net2025),
    .Z(_07011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21683_ (.I0(_07010_),
    .I1(_07011_),
    .S(_06959_),
    .Z(_07012_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input84 (.I(hart_id_i[24]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21685_ (.I0(net115),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(net2025),
    .Z(_07014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21686_ (.I0(net129),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .S(net2025),
    .Z(_07015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21687_ (.I0(_07014_),
    .I1(_07015_),
    .S(_06959_),
    .Z(_07016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21688_ (.I0(net114),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(net2025),
    .Z(_07017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21689_ (.I0(net128),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .S(net2025),
    .Z(_07018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21690_ (.I0(_07017_),
    .I1(_07018_),
    .S(_06959_),
    .Z(_07019_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21691_ (.A1(_07016_),
    .A2(_07019_),
    .Z(_07020_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21692_ (.I0(net113),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(net2025),
    .Z(_07021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21693_ (.I0(net127),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .S(net2025),
    .Z(_07022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21694_ (.I0(_07021_),
    .I1(_07022_),
    .S(_06959_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input83 (.I(hart_id_i[23]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21696_ (.I0(net110),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(net2025),
    .Z(_07025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21697_ (.I0(net123),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .S(net2025),
    .Z(_07026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21698_ (.I0(_07025_),
    .I1(_07026_),
    .S(_06959_),
    .Z(_07027_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _21699_ (.A1(_07012_),
    .A2(_07020_),
    .A3(_07023_),
    .A4(_07027_),
    .ZN(_07028_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21700_ (.A1(_06959_),
    .A2(_07000_),
    .Z(_07029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21701_ (.A1(net2026),
    .A2(_06999_),
    .B(_07029_),
    .ZN(_07030_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21702_ (.A1(_07028_),
    .A2(net1804),
    .ZN(_07031_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21703_ (.A1(_07004_),
    .A2(_07008_),
    .A3(_06998_),
    .A4(_07031_),
    .Z(_07032_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21704_ (.A1(_06973_),
    .A2(_07003_),
    .B(_07032_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input82 (.I(hart_id_i[22]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21706_ (.I(_06967_),
    .ZN(_07035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21707_ (.I0(_06966_),
    .I1(_07035_),
    .S(net2026),
    .Z(_07036_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input81 (.I(hart_id_i[21]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21709_ (.A1(_07004_),
    .A2(_07020_),
    .A3(_06998_),
    .B(_07008_),
    .ZN(_07038_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21710_ (.A1(net1804),
    .A2(_07036_),
    .A3(_07038_),
    .Z(_07039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21711_ (.I0(net122),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(net2025),
    .Z(_07040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21712_ (.I0(net105),
    .I1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .S(net2025),
    .Z(_07041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21713_ (.I0(_07040_),
    .I1(_07041_),
    .S(_06959_),
    .Z(_07042_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input80 (.I(hart_id_i[20]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input79 (.I(hart_id_i[1]),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21716_ (.A1(net1743),
    .A2(_07033_),
    .B(_07039_),
    .C(_07042_),
    .ZN(_07045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21717_ (.A1(_07008_),
    .A2(_07001_),
    .Z(_07046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21718_ (.A1(_07042_),
    .A2(_07046_),
    .Z(_07047_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21719_ (.A1(_06979_),
    .A2(_07028_),
    .A3(_07047_),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input78 (.I(hart_id_i[19]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21721_ (.A1(_06959_),
    .A2(_07041_),
    .Z(_07050_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21722_ (.A1(net2026),
    .A2(_07040_),
    .B(_07050_),
    .ZN(_07051_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21723_ (.A1(_07051_),
    .A2(net1804),
    .Z(_07052_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21724_ (.A1(_06973_),
    .A2(_07052_),
    .Z(_07053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21725_ (.A1(_06959_),
    .A2(_06992_),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21726_ (.A1(net2026),
    .A2(_06991_),
    .B(_07054_),
    .ZN(_07055_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input77 (.I(hart_id_i[18]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input76 (.I(hart_id_i[17]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21729_ (.A1(_07055_),
    .A2(_06996_),
    .ZN(_07058_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21730_ (.A1(_07004_),
    .A2(_07053_),
    .A3(_07058_),
    .Z(_07059_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21731_ (.A1(net1744),
    .A2(_07036_),
    .Z(_07060_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21732_ (.A1(_07048_),
    .A2(_07059_),
    .B(_07060_),
    .ZN(_07061_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21733_ (.A1(net1744),
    .A2(_07045_),
    .B(_07061_),
    .ZN(_07062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21734_ (.I0(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .I1(_07062_),
    .S(net1384),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21735_ (.A1(net99),
    .A2(_10033_),
    .ZN(_07063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21736_ (.A1(_06450_),
    .A2(_07063_),
    .ZN(_07064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21737_ (.A1(net2026),
    .A2(_07064_),
    .B(_10026_),
    .ZN(_07065_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21738_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(_06451_),
    .ZN(_07066_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21739_ (.A1(net2026),
    .A2(_06463_),
    .Z(_07067_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21740_ (.A1(net2024),
    .A2(_07066_),
    .A3(_07067_),
    .Z(_07068_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21741_ (.A1(_07065_),
    .A2(_07068_),
    .ZN(_07069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21742_ (.I0(\id_stage_i.controller_i.instr_fetch_err_i ),
    .I1(_07069_),
    .S(net1384),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21743_ (.A1(net2025),
    .A2(net99),
    .Z(_07070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21744_ (.I0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .I1(_07070_),
    .S(_06450_),
    .Z(_07071_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21745_ (.A1(_07067_),
    .A2(_07071_),
    .Z(_07072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21746_ (.I0(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .I1(_07072_),
    .S(net1384),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21747_ (.A1(net1744),
    .A2(net1743),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21748_ (.I0(\id_stage_i.controller_i.instr_is_compressed_i ),
    .I1(_07073_),
    .S(net1384),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input75 (.I(hart_id_i[16]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21750_ (.I0(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .I1(net1744),
    .S(net1384),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21751_ (.I0(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .I1(_06993_),
    .S(net1384),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21752_ (.I0(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .I1(_06996_),
    .S(net1384),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21753_ (.I0(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .I1(_07004_),
    .S(net1384),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21754_ (.I0(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .I1(_07042_),
    .S(net1384),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input74 (.I(hart_id_i[15]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21756_ (.I0(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .I1(_07001_),
    .S(net1384),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21757_ (.I0(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .I1(_06973_),
    .S(net1384),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21758_ (.I0(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .I1(net1743),
    .S(net1384),
    .Z(_03148_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input73 (.I(hart_id_i[14]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21760_ (.I0(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .I1(_07027_),
    .S(net1384),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21761_ (.I0(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .I1(_07012_),
    .S(net1384),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input72 (.I(hart_id_i[13]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21763_ (.I0(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .I1(_07023_),
    .S(net1384),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input71 (.I(hart_id_i[12]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21765_ (.I0(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .I1(_07019_),
    .S(net1384),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input70 (.I(hart_id_i[11]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21767_ (.I0(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .I1(_07016_),
    .S(net1384),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input69 (.I(hart_id_i[10]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21769_ (.I0(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .I1(_06990_),
    .S(net1384),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21770_ (.I0(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .I1(_06982_),
    .S(net1384),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21771_ (.I0(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .I1(_06986_),
    .S(net1384),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input68 (.I(hart_id_i[0]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21773_ (.A1(_06973_),
    .A2(net1804),
    .Z(_07082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21774_ (.A1(_07036_),
    .A2(_07082_),
    .B(_07042_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21775_ (.A1(net1744),
    .A2(_07083_),
    .Z(_07084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21776_ (.I0(\id_stage_i.controller_i.instr_i[0] ),
    .I1(_07084_),
    .S(net1384),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21777_ (.A1(_07042_),
    .A2(net1804),
    .Z(_07085_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21778_ (.A1(_06973_),
    .A2(_07052_),
    .A3(net1744),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21779_ (.A1(_07051_),
    .A2(_07008_),
    .Z(_07087_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input67 (.I(fetch_enable_i),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21781_ (.I0(_06961_),
    .I1(_06962_),
    .S(net2026),
    .Z(_07089_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(debug_req_i),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(data_rvalid_i),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21784_ (.A1(_06993_),
    .A2(_07087_),
    .B(_07089_),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21785_ (.A1(_07055_),
    .A2(_07085_),
    .B(_07086_),
    .C(_07092_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21786_ (.A1(_07028_),
    .A2(_07053_),
    .Z(_07094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21787_ (.A1(_07089_),
    .A2(_07094_),
    .B(_07055_),
    .ZN(_07095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21788_ (.I0(_07093_),
    .I1(_07095_),
    .S(net1743),
    .Z(_07096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21789_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .I1(_07096_),
    .S(net1384),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21790_ (.A1(net1804),
    .A2(_07087_),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21791_ (.A1(_07060_),
    .A2(_07097_),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21792_ (.A1(_07001_),
    .A2(_07098_),
    .B(_06996_),
    .ZN(_07099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21793_ (.A1(_06993_),
    .A2(_06996_),
    .Z(_07100_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21794_ (.A1(_07004_),
    .A2(_07100_),
    .Z(_07101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21795_ (.A1(_07053_),
    .A2(_07101_),
    .Z(_07102_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(data_rdata_i[9]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21797_ (.A1(_07036_),
    .A2(_07102_),
    .ZN(_07104_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21798_ (.A1(_07099_),
    .A2(_07104_),
    .Z(_07105_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(data_rdata_i[8]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21800_ (.I0(_07087_),
    .I1(_07094_),
    .S(net1743),
    .Z(_07107_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21801_ (.A1(_07089_),
    .A2(_07105_),
    .B1(_07107_),
    .B2(_07099_),
    .ZN(_07108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21802_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .I1(_07108_),
    .S(net1384),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(data_rdata_i[7]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _21804_ (.A1(_06986_),
    .A2(_06990_),
    .A3(_06997_),
    .ZN(_07110_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21805_ (.A1(_06982_),
    .A2(_07110_),
    .Z(_07111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21806_ (.I(_07111_),
    .ZN(_07112_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21807_ (.A1(_07047_),
    .A2(_07112_),
    .Z(_07113_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21808_ (.A1(_06993_),
    .A2(_06996_),
    .ZN(_07114_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21809_ (.A1(_07016_),
    .A2(_07019_),
    .B(_07114_),
    .ZN(_07115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21810_ (.A1(_07051_),
    .A2(_06973_),
    .ZN(_07116_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21811_ (.A1(_06979_),
    .A2(_07087_),
    .B1(_07115_),
    .B2(_07116_),
    .ZN(_07117_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(data_rdata_i[6]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21813_ (.A1(_07042_),
    .A2(_06973_),
    .A3(_07001_),
    .Z(_07119_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21814_ (.A1(_07027_),
    .A2(_07113_),
    .B1(_07117_),
    .B2(net1804),
    .C(_07119_),
    .ZN(_07120_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21815_ (.A1(net1804),
    .A2(_07087_),
    .Z(_07121_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21816_ (.A1(_07089_),
    .A2(net1743),
    .Z(_07122_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21817_ (.A1(_07051_),
    .A2(_07089_),
    .Z(_07123_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21818_ (.A1(_07042_),
    .A2(_07082_),
    .Z(_07124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21819_ (.A1(_07089_),
    .A2(_07036_),
    .Z(_07125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21820_ (.A1(_07124_),
    .A2(_07125_),
    .ZN(_07126_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21821_ (.A1(_07036_),
    .A2(_07123_),
    .B(_07126_),
    .ZN(_07127_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(data_rdata_i[5]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21823_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07127_),
    .B2(_07004_),
    .ZN(_07129_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21824_ (.A1(_07098_),
    .A2(_07120_),
    .B(_07129_),
    .ZN(_07130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21825_ (.I0(net2021),
    .I1(_07130_),
    .S(net1384),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21826_ (.A1(net1744),
    .A2(_07036_),
    .ZN(_07131_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21827_ (.I0(_07016_),
    .I1(_07042_),
    .S(_07004_),
    .Z(_07132_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21828_ (.A1(_07055_),
    .A2(_07132_),
    .Z(_07133_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21829_ (.A1(_07053_),
    .A2(_06996_),
    .A3(_07133_),
    .Z(_07134_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21830_ (.A1(_07012_),
    .A2(_07113_),
    .B(_07134_),
    .ZN(_07135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21831_ (.A1(_07004_),
    .A2(net1804),
    .B(net1743),
    .ZN(_07136_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(data_rdata_i[4]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__oai222_2 _21833_ (.A1(_07052_),
    .A2(net1744),
    .B1(_07131_),
    .B2(_07135_),
    .C1(_07136_),
    .C2(_07051_),
    .ZN(_07138_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(data_rdata_i[3]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21835_ (.I0(\id_stage_i.controller_i.instr_i[13] ),
    .I1(_07138_),
    .S(net1384),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21836_ (.A1(_06979_),
    .A2(_07020_),
    .ZN(_07140_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21837_ (.A1(_07100_),
    .A2(_07140_),
    .ZN(_07141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _21838_ (.A1(_07004_),
    .A2(_07085_),
    .B1(_07113_),
    .B2(_07023_),
    .C1(_07141_),
    .C2(_07053_),
    .ZN(_07142_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21839_ (.A1(net1744),
    .A2(net1743),
    .Z(_07143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21840_ (.A1(_07042_),
    .A2(_07089_),
    .B(_07143_),
    .ZN(_07144_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _21841_ (.A1(_07098_),
    .A2(_07142_),
    .B1(_07144_),
    .B2(net1804),
    .ZN(_07145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21842_ (.I0(\id_stage_i.controller_i.instr_i[14] ),
    .I1(_07145_),
    .S(net1384),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21843_ (.A1(_07042_),
    .A2(_07100_),
    .B(_07004_),
    .ZN(_07146_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21844_ (.A1(_06973_),
    .A2(_07146_),
    .B(_07001_),
    .ZN(_07147_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21845_ (.A1(_06990_),
    .A2(_07147_),
    .Z(_07148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21846_ (.A1(_06979_),
    .A2(_07085_),
    .B(_07046_),
    .ZN(_07149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21847_ (.A1(_07019_),
    .A2(_07113_),
    .B1(_07148_),
    .B2(_07149_),
    .ZN(_07150_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21848_ (.A1(_06990_),
    .A2(_07097_),
    .ZN(_07151_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21849_ (.A1(_07131_),
    .A2(_07150_),
    .A3(_07151_),
    .Z(_07152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21850_ (.A1(_07042_),
    .A2(_07152_),
    .Z(_07153_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21851_ (.A1(_07143_),
    .A2(_07153_),
    .Z(_07154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21852_ (.A1(_07001_),
    .A2(_06990_),
    .B(_07082_),
    .C(net1743),
    .ZN(_07155_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21853_ (.A1(_07004_),
    .A2(_07028_),
    .B(_07053_),
    .ZN(_07156_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21854_ (.A1(_07097_),
    .A2(_07156_),
    .ZN(_07157_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21855_ (.A1(_07089_),
    .A2(net1743),
    .ZN(_07158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21856_ (.A1(_06990_),
    .A2(_07157_),
    .B(_07158_),
    .ZN(_07159_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21857_ (.A1(_07155_),
    .A2(_07159_),
    .B(_07051_),
    .ZN(_07160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21858_ (.A1(_07131_),
    .A2(_07160_),
    .ZN(_07161_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21859_ (.A1(_07008_),
    .A2(_07154_),
    .B1(_07161_),
    .B2(_07152_),
    .ZN(_07162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21860_ (.I0(net2017),
    .I1(_07162_),
    .S(net1384),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21861_ (.I0(_06962_),
    .I1(_06676_),
    .S(net2026),
    .Z(_07163_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21862_ (.A1(_07004_),
    .A2(_07028_),
    .A3(_07008_),
    .Z(_07164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21863_ (.A1(_06982_),
    .A2(_07164_),
    .ZN(_07165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21864_ (.A1(_07042_),
    .A2(_07163_),
    .B1(_07165_),
    .B2(_07052_),
    .ZN(_07166_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21865_ (.A1(net1743),
    .A2(_07166_),
    .B(net1744),
    .ZN(_07167_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21866_ (.I(_07163_),
    .ZN(_07168_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21867_ (.A1(_07004_),
    .A2(_07085_),
    .B1(_07102_),
    .B2(_07168_),
    .C(_07121_),
    .ZN(_07169_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21868_ (.A1(_07016_),
    .A2(_07111_),
    .B(_07047_),
    .ZN(_07170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21869_ (.A1(_07169_),
    .A2(_07170_),
    .ZN(_07171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21870_ (.A1(_06973_),
    .A2(_07001_),
    .ZN(_07172_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _21871_ (.A1(_07001_),
    .A2(_07116_),
    .A3(_07101_),
    .B(_07172_),
    .ZN(_07173_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21872_ (.A1(_07171_),
    .A2(_07173_),
    .Z(_07174_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21873_ (.A1(_07097_),
    .A2(_07171_),
    .B1(_07174_),
    .B2(_06982_),
    .C(net1743),
    .ZN(_07175_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21874_ (.A1(_07167_),
    .A2(_07175_),
    .Z(_07176_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21875_ (.A1(_07051_),
    .A2(_07001_),
    .ZN(_07177_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21876_ (.A1(_07124_),
    .A2(_07163_),
    .ZN(_07178_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21877_ (.A1(_06982_),
    .A2(_07177_),
    .B(_07125_),
    .C(_07178_),
    .ZN(_07179_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21878_ (.A1(_07143_),
    .A2(_07163_),
    .B1(_07176_),
    .B2(_07179_),
    .ZN(_07180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21879_ (.I0(net1965),
    .I1(_07180_),
    .S(net1384),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21880_ (.I0(_06967_),
    .I1(_06747_),
    .S(net2026),
    .Z(_07181_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21881_ (.A1(_06986_),
    .A2(_07157_),
    .B1(_07181_),
    .B2(_07042_),
    .ZN(_07182_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21882_ (.A1(_07051_),
    .A2(_07001_),
    .Z(_07183_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21883_ (.A1(net1744),
    .A2(_07097_),
    .Z(_07184_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21884_ (.A1(net1744),
    .A2(_07183_),
    .B1(_07184_),
    .B2(_06986_),
    .C(_07036_),
    .ZN(_07185_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21885_ (.A1(_07085_),
    .A2(_07113_),
    .Z(_07186_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21886_ (.A1(_07004_),
    .A2(_07186_),
    .ZN(_07187_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21887_ (.A1(_06986_),
    .A2(_07173_),
    .ZN(_07188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21888_ (.A1(_07102_),
    .A2(_07181_),
    .ZN(_07189_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21889_ (.A1(_07184_),
    .A2(_07187_),
    .A3(_07188_),
    .A4(_07189_),
    .Z(_07190_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21890_ (.A1(_07073_),
    .A2(_07126_),
    .ZN(_07191_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21891_ (.A1(_07191_),
    .A2(_07181_),
    .ZN(_07192_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21892_ (.A1(_07158_),
    .A2(_07182_),
    .B1(_07185_),
    .B2(_07190_),
    .C(_07192_),
    .ZN(_07193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21893_ (.I0(net1962),
    .I1(_07193_),
    .S(net1384),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21894_ (.A1(_06993_),
    .A2(net1743),
    .A3(_07123_),
    .A4(_07157_),
    .Z(_07194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21895_ (.I0(_07025_),
    .I1(_06812_),
    .S(net2026),
    .Z(_07195_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21896_ (.A1(_07004_),
    .A2(_07100_),
    .ZN(_07196_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21897_ (.A1(_07051_),
    .A2(_06973_),
    .Z(_07197_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21898_ (.A1(_07196_),
    .A2(_07195_),
    .B(_07197_),
    .ZN(_07198_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21899_ (.A1(_07097_),
    .A2(_07172_),
    .A3(_07187_),
    .A4(_07198_),
    .Z(_07199_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21900_ (.A1(_07055_),
    .A2(_07121_),
    .B(_07199_),
    .ZN(_07200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21901_ (.I0(_07195_),
    .I1(_07200_),
    .S(_07036_),
    .Z(_07201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21902_ (.A1(_06973_),
    .A2(_07195_),
    .B(_07183_),
    .ZN(_07202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21903_ (.A1(_07042_),
    .A2(_07195_),
    .ZN(_07203_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21904_ (.A1(net1743),
    .A2(_07202_),
    .B(_07203_),
    .ZN(_07204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21905_ (.I0(_07201_),
    .I1(_07204_),
    .S(_07089_),
    .Z(_07205_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21906_ (.A1(_07194_),
    .A2(_07205_),
    .Z(_07206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21907_ (.I0(net1960),
    .I1(_07206_),
    .S(net1384),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21908_ (.I0(_07010_),
    .I1(_06836_),
    .S(net2026),
    .Z(_07207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21909_ (.A1(_06996_),
    .A2(_07121_),
    .B1(_07102_),
    .B2(_07207_),
    .ZN(_07208_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21910_ (.A1(_07187_),
    .A2(_07208_),
    .B(_07131_),
    .ZN(_07209_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21911_ (.A1(_07127_),
    .A2(_07207_),
    .Z(_07210_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21912_ (.A1(_07052_),
    .A2(_06996_),
    .A3(_07122_),
    .A4(_07164_),
    .Z(_07211_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21913_ (.A1(_07209_),
    .A2(_07210_),
    .A3(_07211_),
    .Z(_07212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21914_ (.I0(net1958),
    .I1(_07212_),
    .S(net1384),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21915_ (.A1(net1744),
    .A2(_07124_),
    .Z(_07213_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21916_ (.A1(_07089_),
    .A2(_07102_),
    .B(_07213_),
    .C(_07036_),
    .ZN(_07214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21917_ (.I0(\id_stage_i.controller_i.instr_i[1] ),
    .I1(_07214_),
    .S(net1384),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21918_ (.A1(net1743),
    .A2(_07123_),
    .ZN(_07215_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21919_ (.A1(_07008_),
    .A2(net1804),
    .Z(_07216_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21920_ (.A1(_06979_),
    .A2(_06998_),
    .ZN(_07217_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21921_ (.A1(_07028_),
    .A2(net1804),
    .A3(_07217_),
    .Z(_07218_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21922_ (.A1(_07027_),
    .A2(_07218_),
    .B(_07051_),
    .ZN(_07219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21923_ (.A1(_07027_),
    .A2(_07001_),
    .ZN(_07220_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21924_ (.A1(_07219_),
    .A2(_07220_),
    .ZN(_07221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21925_ (.A1(_07027_),
    .A2(_07216_),
    .B1(_07221_),
    .B2(_06973_),
    .ZN(_07222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21926_ (.I0(_07021_),
    .I1(_06852_),
    .S(net2026),
    .Z(_07223_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21927_ (.A1(_07082_),
    .A2(_07196_),
    .B(_07046_),
    .ZN(_07224_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21928_ (.A1(_07042_),
    .A2(_07224_),
    .ZN(_07225_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _21929_ (.A1(_07004_),
    .A2(_07186_),
    .B1(_07223_),
    .B2(_07102_),
    .C1(_07225_),
    .C2(_07027_),
    .ZN(_07226_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21930_ (.A1(_06973_),
    .A2(_07001_),
    .Z(_07227_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21931_ (.I0(_07216_),
    .I1(_07227_),
    .S(_07089_),
    .Z(_07228_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _21932_ (.A1(_07027_),
    .A2(_07051_),
    .A3(_07036_),
    .A4(_07228_),
    .Z(_07229_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21933_ (.A1(_07127_),
    .A2(_07223_),
    .B(_07229_),
    .ZN(_07230_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _21934_ (.A1(_07215_),
    .A2(_07222_),
    .B1(_07226_),
    .B2(_07098_),
    .C(_07230_),
    .ZN(_07231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21935_ (.I0(net2104),
    .I1(_07231_),
    .S(net1384),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21936_ (.I0(_07017_),
    .I1(_06868_),
    .S(net2026),
    .Z(_07232_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21937_ (.A1(_07004_),
    .A2(_07113_),
    .Z(_07233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21938_ (.A1(_07012_),
    .A2(_07225_),
    .B1(_07232_),
    .B2(_07102_),
    .C(_07233_),
    .ZN(_07234_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21939_ (.A1(_07051_),
    .A2(_07089_),
    .ZN(_07235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21940_ (.A1(net1804),
    .A2(net1743),
    .B(_07227_),
    .ZN(_07236_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _21941_ (.A1(_07001_),
    .A2(_07197_),
    .A3(_07131_),
    .Z(_07237_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21942_ (.A1(_07235_),
    .A2(_07236_),
    .B(_07237_),
    .ZN(_07238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21943_ (.A1(_07127_),
    .A2(_07232_),
    .B1(_07238_),
    .B2(_07012_),
    .ZN(_07239_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21944_ (.A1(_07098_),
    .A2(_07234_),
    .B(_07239_),
    .ZN(_07240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21945_ (.I0(net2078),
    .I1(_07240_),
    .S(net1384),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21946_ (.I0(_07014_),
    .I1(_06876_),
    .S(net2026),
    .Z(_07241_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21947_ (.A1(_07023_),
    .A2(_07225_),
    .B1(_07241_),
    .B2(_07102_),
    .C(_07233_),
    .ZN(_07242_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21948_ (.A1(_07215_),
    .A2(_07237_),
    .ZN(_07243_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21949_ (.A1(_07023_),
    .A2(_07001_),
    .Z(_07244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21950_ (.I0(_07016_),
    .I1(_07244_),
    .S(_06973_),
    .Z(_07245_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21951_ (.A1(_07051_),
    .A2(_07125_),
    .A3(_07245_),
    .Z(_07246_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21952_ (.A1(_07127_),
    .A2(_07241_),
    .B1(_07243_),
    .B2(_07023_),
    .C(_07246_),
    .ZN(_07247_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21953_ (.A1(_07098_),
    .A2(_07242_),
    .B(_07247_),
    .ZN(_07248_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(data_rdata_i[31]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21955_ (.I0(net1903),
    .I1(_07248_),
    .S(net1384),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21956_ (.I0(_06989_),
    .I1(_06881_),
    .S(net2026),
    .Z(_07250_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21957_ (.A1(_06979_),
    .A2(_07250_),
    .Z(_07251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21958_ (.I0(_07019_),
    .I1(_07251_),
    .S(_07100_),
    .Z(_07252_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21959_ (.A1(_07019_),
    .A2(_07046_),
    .B1(_07082_),
    .B2(_07252_),
    .ZN(_07253_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21960_ (.A1(_07042_),
    .A2(_07253_),
    .ZN(_07254_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21961_ (.A1(_07233_),
    .A2(_07254_),
    .ZN(_07255_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21962_ (.A1(net1743),
    .A2(_07216_),
    .B(_07123_),
    .ZN(_07256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21963_ (.A1(_07237_),
    .A2(_07256_),
    .ZN(_07257_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21964_ (.A1(_07008_),
    .A2(_07055_),
    .B(_07177_),
    .ZN(_07258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _21965_ (.A1(_07019_),
    .A2(_07257_),
    .B1(_07258_),
    .B2(_07125_),
    .C1(_07250_),
    .C2(_07127_),
    .ZN(_07259_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21966_ (.A1(_07098_),
    .A2(_07255_),
    .B(_07259_),
    .ZN(_07260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21967_ (.I0(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .I1(_07260_),
    .S(net1384),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21968_ (.A1(_07047_),
    .A2(_07111_),
    .B(_07087_),
    .ZN(_07261_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21969_ (.A1(_07131_),
    .A2(_07261_),
    .B(_07215_),
    .ZN(_07262_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21970_ (.A1(_07016_),
    .A2(_07262_),
    .Z(_07263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21971_ (.I0(_07087_),
    .I1(_07085_),
    .S(net1744),
    .Z(_07264_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21972_ (.A1(_06996_),
    .A2(_07036_),
    .A3(_07264_),
    .Z(_07265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21973_ (.I0(_06981_),
    .I1(_06886_),
    .S(net2026),
    .Z(_07266_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _21974_ (.A1(_07127_),
    .A2(_07266_),
    .Z(_07267_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21975_ (.A1(_07053_),
    .A2(_07100_),
    .A3(_07266_),
    .Z(_07268_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21976_ (.A1(_07113_),
    .A2(_07268_),
    .B(_07004_),
    .ZN(_07269_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _21977_ (.A1(_07016_),
    .A2(_07053_),
    .A3(_07114_),
    .ZN(_07270_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _21978_ (.A1(_07269_),
    .A2(_07270_),
    .B(_07098_),
    .ZN(_07271_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _21979_ (.A1(_07263_),
    .A2(_07265_),
    .A3(_07267_),
    .A4(_07271_),
    .Z(_07272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21980_ (.I0(net1899),
    .I1(_07272_),
    .S(net1384),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21981_ (.A1(_07004_),
    .A2(_07053_),
    .A3(_06996_),
    .Z(_07273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21982_ (.I0(_06985_),
    .I1(_06890_),
    .S(net2026),
    .Z(_07274_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _21983_ (.A1(_07055_),
    .A2(_07274_),
    .Z(_07275_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21984_ (.A1(_07047_),
    .A2(_07111_),
    .ZN(_07276_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _21985_ (.A1(_07085_),
    .A2(_07227_),
    .ZN(_07277_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21986_ (.A1(_07276_),
    .A2(_07277_),
    .ZN(_07278_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21987_ (.A1(_07042_),
    .A2(_07111_),
    .ZN(_07279_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21988_ (.A1(_07004_),
    .A2(_07046_),
    .A3(_07279_),
    .Z(_07280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _21989_ (.A1(_07273_),
    .A2(_07275_),
    .B1(_07278_),
    .B2(_07027_),
    .C(_07280_),
    .ZN(_07281_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21990_ (.A1(_07004_),
    .A2(_07060_),
    .ZN(_07282_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _21991_ (.I(_07282_),
    .ZN(_07283_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _21992_ (.A1(_07191_),
    .A2(_07274_),
    .B1(_07283_),
    .B2(_07121_),
    .ZN(_07284_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _21993_ (.A1(_07042_),
    .A2(net1743),
    .A3(_07274_),
    .Z(_07285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21994_ (.A1(_07008_),
    .A2(_07036_),
    .ZN(_07286_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _21995_ (.A1(net1804),
    .A2(_07286_),
    .B(_06979_),
    .C(_07042_),
    .ZN(_07287_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21996_ (.A1(_07285_),
    .A2(_07287_),
    .B(_07089_),
    .ZN(_07288_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _21997_ (.A1(_07098_),
    .A2(_07281_),
    .B(_07284_),
    .C(_07288_),
    .ZN(_07289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _21998_ (.I0(net1898),
    .I1(_07289_),
    .S(net1384),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _21999_ (.A1(_07008_),
    .A2(_07279_),
    .ZN(_07290_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22000_ (.A1(_07019_),
    .A2(_07001_),
    .A3(_07290_),
    .Z(_07291_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22001_ (.A1(_07042_),
    .A2(net1804),
    .A3(_06990_),
    .Z(_07292_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22002_ (.A1(_07291_),
    .A2(_07292_),
    .ZN(_07293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22003_ (.I0(_06991_),
    .I1(_06686_),
    .S(net2026),
    .Z(_07294_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22004_ (.A1(_07055_),
    .A2(_07294_),
    .B(_06996_),
    .C(net1804),
    .ZN(_07295_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22005_ (.A1(_06973_),
    .A2(_07295_),
    .ZN(_07296_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22006_ (.A1(_07046_),
    .A2(_07112_),
    .B1(_07296_),
    .B2(_07051_),
    .ZN(_07297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22007_ (.I0(_07027_),
    .I1(_06990_),
    .S(_06973_),
    .Z(_07298_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22008_ (.A1(_07042_),
    .A2(_07294_),
    .B1(_07298_),
    .B2(_07183_),
    .ZN(_07299_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22009_ (.A1(_07158_),
    .A2(_07299_),
    .ZN(_07300_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22010_ (.A1(_07008_),
    .A2(_06990_),
    .Z(_07301_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22011_ (.I0(_07019_),
    .I1(_07301_),
    .S(net1804),
    .Z(_07302_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22012_ (.A1(_07051_),
    .A2(_07125_),
    .A3(_07302_),
    .Z(_07303_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22013_ (.A1(_07191_),
    .A2(_07294_),
    .B(_07300_),
    .C(_07303_),
    .ZN(_07304_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22014_ (.A1(_07098_),
    .A2(_07293_),
    .B1(_07297_),
    .B2(_07282_),
    .C(_07304_),
    .ZN(_07305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22015_ (.I0(net1897),
    .I1(_07305_),
    .S(net1384),
    .Z(_03175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22016_ (.I0(_06994_),
    .I1(_06690_),
    .S(net2026),
    .Z(_07306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22017_ (.I0(_07012_),
    .I1(_06982_),
    .S(_06973_),
    .Z(_07307_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22018_ (.A1(_07001_),
    .A2(_07307_),
    .Z(_07308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22019_ (.I0(_07306_),
    .I1(_07308_),
    .S(_07123_),
    .Z(_07309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22020_ (.A1(_06982_),
    .A2(_07121_),
    .B1(_07124_),
    .B2(_07306_),
    .ZN(_07310_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22021_ (.A1(_07085_),
    .A2(_07227_),
    .Z(_07311_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22022_ (.A1(_07012_),
    .A2(_07047_),
    .A3(_07111_),
    .Z(_07312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22023_ (.A1(_07016_),
    .A2(_07311_),
    .B(_07312_),
    .ZN(_07313_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22024_ (.A1(_07087_),
    .A2(_07113_),
    .B(_07004_),
    .ZN(_07314_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22025_ (.A1(_07055_),
    .A2(_07306_),
    .B(_07273_),
    .ZN(_07315_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _22026_ (.A1(net1744),
    .A2(_07313_),
    .A3(_07314_),
    .A4(_07315_),
    .Z(_07316_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22027_ (.A1(_07089_),
    .A2(_07310_),
    .B(_07316_),
    .ZN(_07317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22028_ (.I0(_07309_),
    .I1(_07317_),
    .S(_07036_),
    .Z(_07318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22029_ (.I0(net1896),
    .I1(_07318_),
    .S(net1384),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22030_ (.A1(_07098_),
    .A2(_07282_),
    .Z(_07319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22031_ (.I0(_06976_),
    .I1(_06694_),
    .S(net2026),
    .Z(_07320_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22032_ (.A1(_07055_),
    .A2(_07320_),
    .Z(_07321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22033_ (.I0(_07023_),
    .I1(_07004_),
    .S(_07279_),
    .Z(_07322_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22034_ (.A1(_07042_),
    .A2(_06986_),
    .B(_07087_),
    .ZN(_07323_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22035_ (.A1(_06979_),
    .A2(_07172_),
    .B1(_07323_),
    .B2(_07001_),
    .ZN(_07324_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22036_ (.A1(_07273_),
    .A2(_07321_),
    .B1(_07322_),
    .B2(_07046_),
    .C(_07324_),
    .ZN(_07325_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22037_ (.A1(_06986_),
    .A2(_07121_),
    .B1(_07124_),
    .B2(_07320_),
    .ZN(_07326_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22038_ (.I(_07125_),
    .ZN(_07327_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22039_ (.A1(net1743),
    .A2(_07235_),
    .A3(_07320_),
    .ZN(_07328_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22040_ (.A1(_07319_),
    .A2(_07325_),
    .B1(_07326_),
    .B2(_07327_),
    .C(_07328_),
    .ZN(_07329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22041_ (.I0(net1895),
    .I1(_07329_),
    .S(net1384),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22042_ (.I0(_07040_),
    .I1(_06698_),
    .S(net2026),
    .Z(_07330_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22043_ (.A1(_07055_),
    .A2(_07330_),
    .Z(_07331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22044_ (.A1(_07042_),
    .A2(_07055_),
    .B(_07197_),
    .C(_07001_),
    .ZN(_07332_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22045_ (.A1(_07004_),
    .A2(_07001_),
    .B1(_07273_),
    .B2(_07331_),
    .C(_07332_),
    .ZN(_07333_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22046_ (.A1(_06993_),
    .A2(_07121_),
    .A3(_07125_),
    .Z(_07334_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22047_ (.A1(_07127_),
    .A2(_07330_),
    .B(_07334_),
    .ZN(_07335_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22048_ (.A1(_07319_),
    .A2(_07333_),
    .B(_07335_),
    .ZN(_07336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22049_ (.I0(net1894),
    .I1(_07336_),
    .S(net1384),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22050_ (.A1(_07027_),
    .A2(_07102_),
    .B(_07186_),
    .ZN(_07337_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22051_ (.A1(_07158_),
    .A2(_07217_),
    .ZN(_07338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22052_ (.A1(_07027_),
    .A2(_07127_),
    .B1(_07338_),
    .B2(_07094_),
    .ZN(_07339_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22053_ (.A1(_07098_),
    .A2(_07337_),
    .B(_07339_),
    .ZN(_07340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22054_ (.I0(net2145),
    .I1(_07340_),
    .S(net1384),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22055_ (.I0(_06999_),
    .I1(_06703_),
    .S(net2026),
    .Z(_07341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22056_ (.A1(_07020_),
    .A2(_06996_),
    .B(_07055_),
    .ZN(_07342_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22057_ (.A1(_07196_),
    .A2(_07341_),
    .B1(_07342_),
    .B2(_07004_),
    .C(_06997_),
    .ZN(_07343_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22058_ (.A1(_07051_),
    .A2(_06982_),
    .ZN(_07344_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22059_ (.A1(_07197_),
    .A2(_07343_),
    .B(_07344_),
    .ZN(_07345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22060_ (.I0(_07004_),
    .I1(_07345_),
    .S(net1804),
    .Z(_07346_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22061_ (.I(_07319_),
    .ZN(_07347_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22062_ (.A1(_07127_),
    .A2(_07341_),
    .B1(_07346_),
    .B2(_07347_),
    .C(net1385),
    .ZN(_07348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22063_ (.A1(_07947_),
    .A2(net1385),
    .B(_07348_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22064_ (.I0(_06971_),
    .I1(_06708_),
    .S(net2026),
    .Z(_07349_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22065_ (.A1(_07055_),
    .A2(_07349_),
    .B(_06996_),
    .ZN(_07350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22066_ (.A1(_07053_),
    .A2(_07350_),
    .B(_07282_),
    .ZN(_07351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22067_ (.A1(_07127_),
    .A2(_07349_),
    .B(_07351_),
    .C(net1385),
    .ZN(_07352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22068_ (.A1(_08546_),
    .A2(net1385),
    .B(_07352_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22069_ (.A1(_07060_),
    .A2(_07102_),
    .Z(_07353_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22070_ (.A1(_07127_),
    .A2(_07353_),
    .Z(_07354_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22071_ (.A1(_07060_),
    .A2(_07085_),
    .B1(_07354_),
    .B2(_07012_),
    .C(net1385),
    .ZN(_07355_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22072_ (.A1(_07560_),
    .A2(net1385),
    .B(_07355_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22073_ (.A1(_06973_),
    .A2(_07036_),
    .B(_07042_),
    .ZN(_07356_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22074_ (.A1(_07028_),
    .A2(net1743),
    .Z(_07357_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22075_ (.A1(_07197_),
    .A2(_07357_),
    .ZN(_07358_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22076_ (.A1(_07023_),
    .A2(_07356_),
    .B1(_07358_),
    .B2(_07217_),
    .C(_07177_),
    .ZN(_07359_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22077_ (.A1(_06973_),
    .A2(_07101_),
    .B(net1743),
    .ZN(_07360_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22078_ (.A1(net1743),
    .A2(_07277_),
    .B1(_07360_),
    .B2(_07023_),
    .C(net1744),
    .ZN(_07361_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22079_ (.A1(net1744),
    .A2(_07359_),
    .B(_07361_),
    .ZN(_07362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22080_ (.I0(net2189),
    .I1(_07362_),
    .S(net1384),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22081_ (.I(_07113_),
    .ZN(_07363_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22082_ (.A1(_06979_),
    .A2(_07019_),
    .B(_06973_),
    .C(_07100_),
    .ZN(_07364_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22083_ (.A1(_07363_),
    .A2(_07277_),
    .A3(_07364_),
    .Z(_07365_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22084_ (.A1(_07042_),
    .A2(_07089_),
    .B1(_07036_),
    .B2(net1804),
    .ZN(_07366_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22085_ (.A1(_06973_),
    .A2(_07235_),
    .B1(_07366_),
    .B2(_07019_),
    .C(_07131_),
    .ZN(_07367_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22086_ (.A1(_07098_),
    .A2(_07365_),
    .B(_07367_),
    .ZN(_07368_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22087_ (.A1(_07019_),
    .A2(_07073_),
    .B(_07368_),
    .C(net1384),
    .ZN(_07369_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22088_ (.A1(_07581_),
    .A2(net1384),
    .B(_07369_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22089_ (.A1(_07016_),
    .A2(_07102_),
    .B(_07311_),
    .ZN(_07370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22090_ (.A1(_07016_),
    .A2(_07042_),
    .B(_07094_),
    .ZN(_07371_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _22091_ (.A1(_07131_),
    .A2(_07370_),
    .B1(_07371_),
    .B2(_07036_),
    .ZN(_07372_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22092_ (.A1(_07016_),
    .A2(_07191_),
    .B1(_07372_),
    .B2(_07073_),
    .C(net1385),
    .ZN(_07373_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22093_ (.A1(_07566_),
    .A2(net1385),
    .B(_07373_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22094_ (.A1(_07227_),
    .A2(_07283_),
    .ZN(_07374_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22095_ (.A1(_07060_),
    .A2(_07085_),
    .B(_06990_),
    .ZN(_07375_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22096_ (.A1(_06973_),
    .A2(_07375_),
    .Z(_07376_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22097_ (.A1(_07052_),
    .A2(_07131_),
    .B(_06990_),
    .ZN(_07377_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22098_ (.A1(_07374_),
    .A2(_07376_),
    .A3(_07377_),
    .Z(_07378_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22099_ (.A1(_07001_),
    .A2(_07357_),
    .B(_06973_),
    .ZN(_07379_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22100_ (.A1(_07286_),
    .A2(_07379_),
    .B(_07235_),
    .ZN(_07380_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22101_ (.A1(_07027_),
    .A2(_07036_),
    .A3(_07087_),
    .Z(_07381_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _22102_ (.A1(_07004_),
    .A2(net1743),
    .A3(_06998_),
    .A4(_07094_),
    .Z(_07382_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22103_ (.A1(_07381_),
    .A2(_07382_),
    .B(_07089_),
    .ZN(_07383_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22104_ (.A1(_07378_),
    .A2(_07380_),
    .B(_07383_),
    .ZN(_07384_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(data_rdata_i[30]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22106_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .I1(_07384_),
    .S(net1384),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22107_ (.I0(_07087_),
    .I1(_07227_),
    .S(net1744),
    .Z(_07386_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22108_ (.A1(_07012_),
    .A2(_07036_),
    .A3(_07386_),
    .ZN(_07387_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22109_ (.I0(_07124_),
    .I1(_07277_),
    .S(net1744),
    .Z(_07388_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22110_ (.A1(_07235_),
    .A2(_07379_),
    .B1(_07388_),
    .B2(net1743),
    .C(_06982_),
    .ZN(_07389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22111_ (.A1(_07387_),
    .A2(_07389_),
    .ZN(_07390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22112_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .I1(_07390_),
    .S(net1384),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22113_ (.A1(_07023_),
    .A2(_07008_),
    .B1(_07227_),
    .B2(_07016_),
    .ZN(_07391_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22114_ (.A1(_07042_),
    .A2(_07327_),
    .A3(_07391_),
    .Z(_07392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22115_ (.A1(_07052_),
    .A2(_06986_),
    .B(_07244_),
    .ZN(_07393_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22116_ (.A1(_07008_),
    .A2(_07131_),
    .A3(_07393_),
    .Z(_07394_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22117_ (.A1(_06973_),
    .A2(_07123_),
    .A3(_07357_),
    .Z(_07395_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22118_ (.A1(_07042_),
    .A2(_07060_),
    .B(_07395_),
    .ZN(_07396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22119_ (.I0(_07008_),
    .I1(_07124_),
    .S(_07089_),
    .Z(_07397_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22120_ (.A1(_07001_),
    .A2(_07396_),
    .B1(_07397_),
    .B2(net1743),
    .C(_06986_),
    .ZN(_07398_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22121_ (.A1(_07392_),
    .A2(_07394_),
    .A3(_07398_),
    .ZN(_07399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22122_ (.I0(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .I1(_07399_),
    .S(net1384),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22123_ (.I0(\cs_registers_i.pc_id_i[10] ),
    .I1(\cs_registers_i.pc_if_i[10] ),
    .S(net1383),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22124_ (.I0(\cs_registers_i.pc_id_i[11] ),
    .I1(\cs_registers_i.pc_if_i[11] ),
    .S(net1383),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22125_ (.I0(\cs_registers_i.pc_id_i[12] ),
    .I1(\cs_registers_i.pc_if_i[12] ),
    .S(net1383),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22126_ (.I0(\cs_registers_i.pc_id_i[13] ),
    .I1(\cs_registers_i.pc_if_i[13] ),
    .S(net1383),
    .Z(_03192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22127_ (.I0(\cs_registers_i.pc_id_i[14] ),
    .I1(\cs_registers_i.pc_if_i[14] ),
    .S(net1383),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22128_ (.I0(\cs_registers_i.pc_id_i[15] ),
    .I1(\cs_registers_i.pc_if_i[15] ),
    .S(net1383),
    .Z(_03194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22129_ (.I0(\cs_registers_i.pc_id_i[16] ),
    .I1(\cs_registers_i.pc_if_i[16] ),
    .S(net1383),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(data_rdata_i[2]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22131_ (.I0(\cs_registers_i.pc_id_i[17] ),
    .I1(\cs_registers_i.pc_if_i[17] ),
    .S(net1383),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22132_ (.I0(\cs_registers_i.pc_id_i[18] ),
    .I1(\cs_registers_i.pc_if_i[18] ),
    .S(net1383),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22133_ (.I0(\cs_registers_i.pc_id_i[19] ),
    .I1(\cs_registers_i.pc_if_i[19] ),
    .S(net1383),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22134_ (.I0(\cs_registers_i.pc_id_i[1] ),
    .I1(net2026),
    .S(net1384),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22135_ (.I0(\cs_registers_i.pc_id_i[20] ),
    .I1(\cs_registers_i.pc_if_i[20] ),
    .S(net1383),
    .Z(_03200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22136_ (.I0(\cs_registers_i.pc_id_i[21] ),
    .I1(\cs_registers_i.pc_if_i[21] ),
    .S(net1383),
    .Z(_03201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22137_ (.I0(\cs_registers_i.pc_id_i[22] ),
    .I1(\cs_registers_i.pc_if_i[22] ),
    .S(net1383),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22138_ (.I0(\cs_registers_i.pc_id_i[23] ),
    .I1(\cs_registers_i.pc_if_i[23] ),
    .S(net1383),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22139_ (.I0(\cs_registers_i.pc_id_i[24] ),
    .I1(\cs_registers_i.pc_if_i[24] ),
    .S(net1383),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22140_ (.I0(\cs_registers_i.pc_id_i[25] ),
    .I1(\cs_registers_i.pc_if_i[25] ),
    .S(net1383),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(data_rdata_i[29]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22142_ (.I0(\cs_registers_i.pc_id_i[26] ),
    .I1(\cs_registers_i.pc_if_i[26] ),
    .S(net1383),
    .Z(_03206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22143_ (.I0(\cs_registers_i.pc_id_i[27] ),
    .I1(\cs_registers_i.pc_if_i[27] ),
    .S(net1383),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22144_ (.I0(\cs_registers_i.pc_id_i[28] ),
    .I1(\cs_registers_i.pc_if_i[28] ),
    .S(net1383),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22145_ (.I0(\cs_registers_i.pc_id_i[29] ),
    .I1(\cs_registers_i.pc_if_i[29] ),
    .S(net1383),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22146_ (.I0(\cs_registers_i.pc_id_i[2] ),
    .I1(\cs_registers_i.pc_if_i[2] ),
    .S(net1383),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22147_ (.I0(\cs_registers_i.pc_id_i[30] ),
    .I1(\cs_registers_i.pc_if_i[30] ),
    .S(net1383),
    .Z(_03211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22148_ (.I0(\cs_registers_i.pc_id_i[31] ),
    .I1(\cs_registers_i.pc_if_i[31] ),
    .S(net1383),
    .Z(_03212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22149_ (.I0(\cs_registers_i.pc_id_i[3] ),
    .I1(\cs_registers_i.pc_if_i[3] ),
    .S(net1383),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22150_ (.I0(\cs_registers_i.pc_id_i[4] ),
    .I1(\cs_registers_i.pc_if_i[4] ),
    .S(net1383),
    .Z(_03214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22151_ (.I0(\cs_registers_i.pc_id_i[5] ),
    .I1(\cs_registers_i.pc_if_i[5] ),
    .S(net1383),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22152_ (.I0(\cs_registers_i.pc_id_i[6] ),
    .I1(\cs_registers_i.pc_if_i[6] ),
    .S(net1383),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22153_ (.I0(\cs_registers_i.pc_id_i[7] ),
    .I1(\cs_registers_i.pc_if_i[7] ),
    .S(net1383),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22154_ (.I0(\cs_registers_i.pc_id_i[8] ),
    .I1(\cs_registers_i.pc_if_i[8] ),
    .S(net1383),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22155_ (.I0(\cs_registers_i.pc_id_i[9] ),
    .I1(\cs_registers_i.pc_if_i[9] ),
    .S(net1383),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22156_ (.A1(net1834),
    .A2(_10080_),
    .ZN(net254));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _22157_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .ZN(_07402_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22158_ (.A1(_09653_),
    .A2(_07402_),
    .ZN(_07403_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22159_ (.A1(_05781_),
    .A2(net254),
    .A3(_07403_),
    .Z(core_busy_d));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22160_ (.A1(clknet_1_0__leaf_clk_i),
    .A2(net2467),
    .Z(clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22161_ (.I(_01356_),
    .ZN(_07404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22162_ (.I0(_01366_),
    .I1(_07404_),
    .S(net2022),
    .Z(_07405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22163_ (.I0(_07405_),
    .I1(_01357_),
    .S(_06914_),
    .Z(net186));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(data_rdata_i[28]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22165_ (.A1(_01366_),
    .A2(net1522),
    .B(net1885),
    .ZN(_07407_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(data_rdata_i[27]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(data_rdata_i[26]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22168_ (.A1(net1533),
    .A2(net1534),
    .B(\load_store_unit_i.handle_misaligned_q ),
    .C(_06914_),
    .ZN(_07410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22169_ (.A1(_01364_),
    .A2(_10133_),
    .ZN(_07411_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _22170_ (.A1(_10133_),
    .A2(_07407_),
    .B(_07410_),
    .C(_07411_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22171_ (.A1(_01361_),
    .A2(_10133_),
    .Z(_07412_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22172_ (.A1(net2022),
    .A2(_01359_),
    .B(_06914_),
    .ZN(_07413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22173_ (.A1(_01358_),
    .A2(_06914_),
    .B(_07413_),
    .C(\load_store_unit_i.handle_misaligned_q ),
    .ZN(_07414_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22174_ (.A1(net1534),
    .A2(\load_store_unit_i.handle_misaligned_q ),
    .A3(_06914_),
    .Z(_07415_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _22175_ (.A1(_07412_),
    .A2(_07414_),
    .A3(_07415_),
    .Z(net188));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22176_ (.A1(net2022),
    .A2(_06914_),
    .Z(_07416_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _22177_ (.A1(net2022),
    .A2(net1533),
    .B(net1534),
    .C(_06914_),
    .ZN(_07417_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22178_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_07416_),
    .B(_07417_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22179_ (.I(_10129_),
    .ZN(_07418_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22180_ (.A1(_07550_),
    .A2(_07418_),
    .B(net2081),
    .ZN(net190));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(data_rdata_i[25]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(data_rdata_i[24]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22183_ (.A1(net1534),
    .A2(net1713),
    .B1(net2190),
    .B2(net1533),
    .C1(net1522),
    .C2(net1760),
    .ZN(_07421_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22184_ (.I(_07421_),
    .ZN(_07422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22185_ (.I0(net1798),
    .I1(_07422_),
    .S(net1520),
    .Z(net191));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(data_rdata_i[23]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(data_rdata_i[22]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22188_ (.A1(net1522),
    .A2(net1740),
    .B1(net2479),
    .B2(net1534),
    .C1(net1758),
    .C2(net1533),
    .ZN(_07425_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22189_ (.I(_07425_),
    .ZN(_07426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22190_ (.I0(net1711),
    .I1(_07426_),
    .S(net1520),
    .Z(net192));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22191_ (.A1(net1522),
    .A2(net1749),
    .B1(net1767),
    .B2(net1534),
    .C1(net1757),
    .C2(net1533),
    .ZN(_07427_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22192_ (.I(_07427_),
    .ZN(_07428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22193_ (.I0(net2158),
    .I1(_07428_),
    .S(net1520),
    .Z(net193));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22194_ (.I(net1522),
    .ZN(_07429_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(data_rdata_i[21]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22196_ (.A1(net1534),
    .A2(net1766),
    .B1(net1756),
    .B2(net1533),
    .ZN(_07431_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22197_ (.A1(_07429_),
    .A2(net1794),
    .B(_07431_),
    .ZN(_07432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22198_ (.I0(net2136),
    .I1(_07432_),
    .S(net1520),
    .Z(net194));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22199_ (.A1(net1522),
    .A2(net1792),
    .B1(net1763),
    .B2(net1534),
    .C1(net1755),
    .C2(net1533),
    .ZN(_07433_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22200_ (.I(_07433_),
    .ZN(_07434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22201_ (.I0(net2157),
    .I1(_07434_),
    .S(net1520),
    .Z(net195));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22202_ (.A1(net1522),
    .A2(net1790),
    .B1(net1762),
    .B2(net1534),
    .C1(net1753),
    .C2(net1533),
    .ZN(_07435_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22203_ (.I(_07435_),
    .ZN(_07436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22204_ (.I0(net2192),
    .I1(_07436_),
    .S(net1520),
    .Z(net196));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22205_ (.A1(net1522),
    .A2(net1788),
    .B1(net1761),
    .B2(net1534),
    .C1(net1719),
    .C2(net1533),
    .ZN(_07437_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22206_ (.I(_07437_),
    .ZN(_07438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22207_ (.I0(net2187),
    .I1(_07438_),
    .S(net1520),
    .Z(net197));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(data_rdata_i[20]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22209_ (.A1(net1533),
    .A2(net1798),
    .B1(net1760),
    .B2(net1534),
    .C1(net1713),
    .C2(net1522),
    .ZN(_07440_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22210_ (.I(_07440_),
    .ZN(_07441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22211_ (.I0(net2190),
    .I1(_07441_),
    .S(net1520),
    .Z(net198));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22212_ (.A1(net1533),
    .A2(net2185),
    .B1(net1759),
    .B2(net1534),
    .C1(net1709),
    .C2(net1522),
    .ZN(_07442_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22213_ (.I(_07442_),
    .ZN(_07443_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(data_rdata_i[1]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22215_ (.I0(net1769),
    .I1(_07443_),
    .S(net1520),
    .Z(net199));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22216_ (.A1(net1533),
    .A2(net1740),
    .B1(net1758),
    .B2(net1534),
    .C1(net1711),
    .C2(net1522),
    .ZN(_07445_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22217_ (.I(_07445_),
    .ZN(_07446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22218_ (.I0(net2479),
    .I1(_07446_),
    .S(net1520),
    .Z(net200));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22219_ (.A1(net1533),
    .A2(net1749),
    .B1(net1757),
    .B2(net1534),
    .C1(net2158),
    .C2(net1522),
    .ZN(_07447_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22220_ (.I(_07447_),
    .ZN(_07448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22221_ (.I0(net1767),
    .I1(_07448_),
    .S(net1520),
    .Z(net201));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22222_ (.A1(net1534),
    .A2(net1709),
    .B1(net1769),
    .B2(net1533),
    .C1(net1522),
    .C2(net1759),
    .ZN(_07449_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22223_ (.I(_07449_),
    .ZN(_07450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22224_ (.I0(net2185),
    .I1(_07450_),
    .S(net1520),
    .Z(net202));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22225_ (.A1(net1533),
    .A2(_05997_),
    .B1(net1756),
    .B2(net1534),
    .C1(net2136),
    .C2(net1522),
    .ZN(_07451_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22226_ (.A1(_01366_),
    .A2(net1729),
    .Z(_07452_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22227_ (.A1(net1520),
    .A2(_07451_),
    .B(_07452_),
    .ZN(net203));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22228_ (.A1(net1533),
    .A2(net1792),
    .B1(net1755),
    .B2(net1534),
    .C1(net2157),
    .C2(net1522),
    .ZN(_07453_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22229_ (.I(_07453_),
    .ZN(_07454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22230_ (.I0(net1763),
    .I1(_07454_),
    .S(net1520),
    .Z(net204));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22231_ (.A1(net1533),
    .A2(net1790),
    .B1(net1753),
    .B2(net1534),
    .C1(net2192),
    .C2(net1522),
    .ZN(_07455_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22232_ (.I(_07455_),
    .ZN(_07456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22233_ (.I0(net1762),
    .I1(_07456_),
    .S(net1520),
    .Z(net205));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22234_ (.A1(net1533),
    .A2(net1788),
    .B1(net1719),
    .B2(net1534),
    .C1(net2187),
    .C2(net1522),
    .ZN(_07457_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22235_ (.I(_07457_),
    .ZN(_07458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22236_ (.I0(net1761),
    .I1(_07458_),
    .S(net1520),
    .Z(net206));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22237_ (.A1(net1534),
    .A2(net1798),
    .B1(net1713),
    .B2(net1533),
    .C1(net1522),
    .C2(net2190),
    .ZN(_07459_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22238_ (.I(_07459_),
    .ZN(_07460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22239_ (.I0(net1760),
    .I1(_07460_),
    .S(net1520),
    .Z(net207));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22240_ (.A1(net1534),
    .A2(net2185),
    .B1(net1709),
    .B2(net1533),
    .C1(net1522),
    .C2(net1769),
    .ZN(_07461_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22241_ (.I(_07461_),
    .ZN(_07462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22242_ (.I0(net1759),
    .I1(_07462_),
    .S(net1520),
    .Z(net208));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22243_ (.A1(net1534),
    .A2(net1740),
    .B1(net1711),
    .B2(net1533),
    .C1(net1522),
    .C2(net2479),
    .ZN(_07463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22244_ (.I(_07463_),
    .ZN(_07464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22245_ (.I0(net1758),
    .I1(_07464_),
    .S(net1520),
    .Z(net209));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22246_ (.A1(net1534),
    .A2(net1749),
    .B1(net2158),
    .B2(net1533),
    .C1(net1522),
    .C2(net1767),
    .ZN(_07465_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22247_ (.I(_07465_),
    .ZN(_07466_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(data_rdata_i[19]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22249_ (.I0(net1757),
    .I1(_07466_),
    .S(net1520),
    .Z(net210));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22250_ (.A1(net1534),
    .A2(_05997_),
    .B1(net2136),
    .B2(net1533),
    .ZN(_07468_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22251_ (.A1(_07429_),
    .A2(net1729),
    .B(_07468_),
    .ZN(_07469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22252_ (.I0(net1756),
    .I1(_07469_),
    .S(net1520),
    .Z(net211));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22253_ (.A1(net1534),
    .A2(net1792),
    .B1(net2157),
    .B2(net1533),
    .C1(net1522),
    .C2(net1763),
    .ZN(_07470_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22254_ (.I(_07470_),
    .ZN(_07471_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22255_ (.I0(net1755),
    .I1(_07471_),
    .S(net1520),
    .Z(net212));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22256_ (.A1(net1534),
    .A2(net1711),
    .B1(net2479),
    .B2(net1533),
    .C1(net1522),
    .C2(net1758),
    .ZN(_07472_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22257_ (.I(_07472_),
    .ZN(_07473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22258_ (.I0(net1740),
    .I1(_07473_),
    .S(net1520),
    .Z(net213));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22259_ (.A1(net1534),
    .A2(net1790),
    .B1(net2192),
    .B2(net1533),
    .C1(net1522),
    .C2(net1762),
    .ZN(_07474_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22260_ (.I(_07474_),
    .ZN(_07475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22261_ (.I0(net1753),
    .I1(_07475_),
    .S(net1520),
    .Z(net214));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22262_ (.A1(net1534),
    .A2(net1788),
    .B1(net2187),
    .B2(net1533),
    .C1(net1522),
    .C2(net1761),
    .ZN(_07476_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22263_ (.I(_07476_),
    .ZN(_07477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22264_ (.I0(net1719),
    .I1(_07477_),
    .S(net1520),
    .Z(net215));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22265_ (.A1(net1534),
    .A2(net2158),
    .B1(net1767),
    .B2(net1533),
    .C1(net1522),
    .C2(net1757),
    .ZN(_07478_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22266_ (.I(_07478_),
    .ZN(_07479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22267_ (.I0(net1749),
    .I1(_07479_),
    .S(net1520),
    .Z(net216));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22268_ (.A1(net1534),
    .A2(net2136),
    .B1(net1766),
    .B2(net1533),
    .C1(net1522),
    .C2(net1756),
    .ZN(_07480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22269_ (.I0(net1794),
    .I1(_07480_),
    .S(net1520),
    .Z(_07481_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22270_ (.I(_07481_),
    .ZN(net217));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22271_ (.A1(net1534),
    .A2(net2157),
    .B1(net1763),
    .B2(net1533),
    .C1(net1522),
    .C2(net1755),
    .ZN(_07482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22272_ (.I(_07482_),
    .ZN(_07483_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22273_ (.I0(net1792),
    .I1(_07483_),
    .S(net1520),
    .Z(net218));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22274_ (.A1(net1534),
    .A2(net2192),
    .B1(net1762),
    .B2(net1533),
    .C1(net1522),
    .C2(net1753),
    .ZN(_07484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22275_ (.I(_07484_),
    .ZN(_07485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22276_ (.I0(net1790),
    .I1(_07485_),
    .S(net1520),
    .Z(net219));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22277_ (.A1(net1534),
    .A2(net2187),
    .B1(net1761),
    .B2(net1533),
    .C1(net1522),
    .C2(net1719),
    .ZN(_07486_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22278_ (.I(_07486_),
    .ZN(_07487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22279_ (.I0(net1788),
    .I1(_07487_),
    .S(net1520),
    .Z(net220));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22280_ (.A1(net1522),
    .A2(net1798),
    .B1(net2190),
    .B2(net1534),
    .C1(net1760),
    .C2(net1533),
    .ZN(_07488_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22281_ (.I(_07488_),
    .ZN(_07489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22282_ (.I0(net1713),
    .I1(_07489_),
    .S(net1520),
    .Z(net221));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _22283_ (.A1(net1522),
    .A2(net2185),
    .B1(net1769),
    .B2(net1534),
    .C1(net1759),
    .C2(net1533),
    .ZN(_07490_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22284_ (.I(_07490_),
    .ZN(_07491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22285_ (.I0(net1709),
    .I1(_07491_),
    .S(net1520),
    .Z(net222));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22286_ (.A1(_10128_),
    .A2(_05798_),
    .Z(\id_stage_i.branch_set_d ));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _22287_ (.A1(net133),
    .A2(_10012_),
    .Z(_07492_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22288_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(_07492_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .ZN(_07493_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22289_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_10012_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .ZN(_07494_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22290_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net133),
    .A3(_07494_),
    .Z(_07495_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22291_ (.A1(net100),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .ZN(_07496_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22292_ (.A1(_07493_),
    .A2(_07495_),
    .B(_07496_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22293_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net100),
    .Z(_07497_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22294_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .A2(_07497_),
    .ZN(_07498_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22295_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net133),
    .B1(_07494_),
    .B2(_07498_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22296_ (.I0(_06450_),
    .I1(net1819),
    .S(_06469_),
    .Z(_07499_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _22297_ (.A1(net1819),
    .A2(_06670_),
    .B1(_07499_),
    .B2(_10023_),
    .C(_10012_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22298_ (.A1(net1393),
    .A2(net1819),
    .A3(_06457_),
    .Z(_07500_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22299_ (.A1(net2023),
    .A2(net1393),
    .A3(_06457_),
    .ZN(_07501_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _22300_ (.A1(_06448_),
    .A2(_06458_),
    .B1(_07500_),
    .B2(_06450_),
    .C(_07501_),
    .ZN(_07502_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22301_ (.A1(net1589),
    .A2(_07502_),
    .Z(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _22302_ (.A1(net1589),
    .A2(_06469_),
    .A3(_06488_),
    .Z(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22303_ (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .ZN(_07503_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22304_ (.A1(_07503_),
    .A2(net133),
    .ZN(_07504_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22305_ (.A1(net100),
    .A2(net254),
    .B1(_07504_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .ZN(_07505_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _22306_ (.I(_07505_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _22307_ (.A1(net254),
    .A2(_07497_),
    .ZN(_07506_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _22308_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net133),
    .B1(_07506_),
    .B2(_07503_),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _22309_ (.A1(net1834),
    .A2(_10080_),
    .B(net100),
    .ZN(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _22310_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_05745_),
    .A3(_05794_),
    .ZN(_07507_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _22311_ (.A1(_06478_),
    .A2(_05777_),
    .B(net1809),
    .ZN(_07508_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _22312_ (.A1(_03436_),
    .A2(_07508_),
    .Z(_07509_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _22313_ (.A1(_09911_),
    .A2(_07507_),
    .A3(_07509_),
    .B1(_10012_),
    .B2(net1386),
    .ZN(\if_stage_i.instr_valid_id_d ));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22314_ (.A(_00007_),
    .B(_00008_),
    .CI(_00009_),
    .CO(_00010_),
    .S(_00011_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22315_ (.A(_00012_),
    .B(_00013_),
    .CI(_00014_),
    .CO(_00015_),
    .S(_00016_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22316_ (.A(_00017_),
    .B(_00018_),
    .CI(_00019_),
    .CO(_11106_),
    .S(_00020_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22317_ (.A(_00021_),
    .B(_00022_),
    .CI(_00023_),
    .CO(_11107_),
    .S(_11108_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22318_ (.A(_00024_),
    .B(_00025_),
    .CI(_00026_),
    .CO(_11109_),
    .S(_11110_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22319_ (.A(_00027_),
    .B(_11106_),
    .CI(_11110_),
    .CO(_00028_),
    .S(_00029_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22320_ (.A(_00030_),
    .B(_00031_),
    .CI(_00032_),
    .CO(_11111_),
    .S(_11112_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22321_ (.A(_00033_),
    .B(_00034_),
    .CI(_00035_),
    .CO(_11113_),
    .S(_00036_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22322_ (.A(_00037_),
    .B(_11112_),
    .CI(_11109_),
    .CO(_11114_),
    .S(_00038_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22323_ (.A(_00039_),
    .B(_00040_),
    .CI(_11115_),
    .CO(_11116_),
    .S(_11117_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22324_ (.A(_00041_),
    .B(_00042_),
    .CI(_00043_),
    .CO(_11118_),
    .S(_11119_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22325_ (.A(_00044_),
    .B(_00045_),
    .CI(_00046_),
    .CO(_00047_),
    .S(_11120_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22326_ (.A(_11119_),
    .B(_11111_),
    .CI(_11120_),
    .CO(_11121_),
    .S(_11122_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22327_ (.A(_11122_),
    .B(_11114_),
    .CI(_00048_),
    .CO(_00049_),
    .S(_00050_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22328_ (.A(_00051_),
    .B(_00052_),
    .CI(_00053_),
    .CO(_11123_),
    .S(_11124_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22329_ (.A(_00054_),
    .B(_00055_),
    .CI(_00056_),
    .CO(_11125_),
    .S(_00057_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22330_ (.A(_11124_),
    .B(_11118_),
    .CI(_00058_),
    .CO(_11126_),
    .S(_11127_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22331_ (.A(_11127_),
    .B(_11121_),
    .CI(_00059_),
    .CO(_00060_),
    .S(_00061_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22332_ (.A(_00062_),
    .B(_00063_),
    .CI(_11128_),
    .CO(_11129_),
    .S(_11130_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22333_ (.A(_00064_),
    .B(_00065_),
    .CI(_00066_),
    .CO(_11131_),
    .S(_11132_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22334_ (.A(_00067_),
    .B(_00068_),
    .CI(_00069_),
    .CO(_11133_),
    .S(_00070_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22335_ (.A(_00071_),
    .B(_11123_),
    .CI(_11132_),
    .CO(_11134_),
    .S(_11135_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22336_ (.A(_00072_),
    .B(_00073_),
    .CI(_00074_),
    .CO(_00075_),
    .S(_00076_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22337_ (.A(_11125_),
    .B(_00077_),
    .CI(_11136_),
    .CO(_11137_),
    .S(_00078_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22338_ (.A(_11135_),
    .B(_11126_),
    .CI(_00079_),
    .CO(_11138_),
    .S(_00080_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22339_ (.A(_00081_),
    .B(_00082_),
    .CI(_11139_),
    .CO(_11140_),
    .S(_11141_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22340_ (.A(_00083_),
    .B(_00084_),
    .CI(_00085_),
    .CO(_00086_),
    .S(_00087_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22341_ (.A(_00088_),
    .B(_00089_),
    .CI(_00090_),
    .CO(_11142_),
    .S(_11143_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22342_ (.A(_00091_),
    .B(_00092_),
    .CI(_00093_),
    .CO(_11144_),
    .S(_00094_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22343_ (.A(_11143_),
    .B(_11131_),
    .CI(_00095_),
    .CO(_11145_),
    .S(_11146_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22344_ (.A(_00096_),
    .B(_00097_),
    .CI(_00098_),
    .CO(_00099_),
    .S(_00100_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22345_ (.A(_11133_),
    .B(_00101_),
    .CI(_00102_),
    .CO(_11147_),
    .S(_00103_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22346_ (.A(_11146_),
    .B(_11134_),
    .CI(_00104_),
    .CO(_11148_),
    .S(_11149_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22347_ (.A(_11138_),
    .B(_11149_),
    .CI(_00105_),
    .CO(_00106_),
    .S(_00107_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22348_ (.A(_00108_),
    .B(_00109_),
    .CI(_00110_),
    .CO(_11150_),
    .S(_11151_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22349_ (.A(_00111_),
    .B(_00112_),
    .CI(_00113_),
    .CO(_00114_),
    .S(_00115_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22350_ (.A(_11151_),
    .B(_00116_),
    .CI(_11142_),
    .CO(_11152_),
    .S(_11153_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22351_ (.A(_00117_),
    .B(_00118_),
    .CI(_00119_),
    .CO(_11154_),
    .S(_00120_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22352_ (.A(_00121_),
    .B(_00122_),
    .CI(_11144_),
    .CO(_11155_),
    .S(_00123_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22353_ (.A(_00124_),
    .B(_11145_),
    .CI(_11153_),
    .CO(_11156_),
    .S(_11157_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22354_ (.A(_11157_),
    .B(_11148_),
    .CI(_00125_),
    .CO(_00126_),
    .S(_00127_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22355_ (.A(_00128_),
    .B(_00129_),
    .CI(_11158_),
    .CO(_11159_),
    .S(_11160_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22356_ (.A(_00130_),
    .B(_00131_),
    .CI(_00132_),
    .CO(_11161_),
    .S(_11162_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22357_ (.A(_00133_),
    .B(_00134_),
    .CI(_00135_),
    .CO(_00136_),
    .S(_00137_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22358_ (.A(_11162_),
    .B(_11150_),
    .CI(_00138_),
    .CO(_11163_),
    .S(_11164_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22359_ (.A(_00139_),
    .B(_00140_),
    .CI(_00141_),
    .CO(_11165_),
    .S(_11166_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22360_ (.A(_11154_),
    .B(_11166_),
    .CI(_00142_),
    .CO(_00143_),
    .S(_11167_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22361_ (.A(_11152_),
    .B(_11164_),
    .CI(_11167_),
    .CO(_11168_),
    .S(_11169_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22362_ (.A(_00144_),
    .B(_00145_),
    .CI(_00146_),
    .CO(_00147_),
    .S(_00148_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22363_ (.A(_00149_),
    .B(_11156_),
    .CI(_11169_),
    .CO(_00150_),
    .S(_00151_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22364_ (.A(_11170_),
    .B(_00152_),
    .CI(_00153_),
    .CO(_11171_),
    .S(_11172_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22365_ (.A(_00154_),
    .B(_00155_),
    .CI(_00156_),
    .CO(_11173_),
    .S(_11174_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22366_ (.A(_00157_),
    .B(_00158_),
    .CI(_00159_),
    .CO(_00160_),
    .S(_00161_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22367_ (.A(_00162_),
    .B(_11161_),
    .CI(_11174_),
    .CO(_11175_),
    .S(_11176_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22368_ (.A(_00163_),
    .B(_00164_),
    .CI(_00165_),
    .CO(_11177_),
    .S(_11178_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22369_ (.A(_11165_),
    .B(_11178_),
    .CI(_00166_),
    .CO(_11179_),
    .S(_11180_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22370_ (.A(_11180_),
    .B(_11163_),
    .CI(_11176_),
    .CO(_11181_),
    .S(_11182_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22371_ (.A(_00167_),
    .B(_00168_),
    .CI(_00169_),
    .CO(_11183_),
    .S(_00170_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22372_ (.A(_00171_),
    .B(_00172_),
    .CI(_00173_),
    .CO(_00174_),
    .S(_11184_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22373_ (.A(_00175_),
    .B(_11185_),
    .CI(_11184_),
    .CO(_00176_),
    .S(_00177_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22374_ (.A(_11168_),
    .B(_11182_),
    .CI(_00178_),
    .CO(_11186_),
    .S(_00179_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22375_ (.A(_11187_),
    .B(_00180_),
    .CI(_00181_),
    .CO(_11188_),
    .S(_11189_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22376_ (.A(_00182_),
    .B(_00183_),
    .CI(_00184_),
    .CO(_11190_),
    .S(_11191_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22377_ (.A(_00185_),
    .B(_00186_),
    .CI(_00187_),
    .CO(_00188_),
    .S(_00189_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22378_ (.A(_00190_),
    .B(_11173_),
    .CI(_11191_),
    .CO(_11192_),
    .S(_11193_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22379_ (.A(_00191_),
    .B(_00192_),
    .CI(_00193_),
    .CO(_11194_),
    .S(_11195_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22380_ (.A(_11177_),
    .B(_11195_),
    .CI(_00194_),
    .CO(_00195_),
    .S(_11196_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22381_ (.A(_11196_),
    .B(_11175_),
    .CI(_11193_),
    .CO(_11197_),
    .S(_11198_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22382_ (.A(_00196_),
    .B(_00197_),
    .CI(_00198_),
    .CO(_11199_),
    .S(_11200_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22383_ (.A(_00199_),
    .B(_11183_),
    .CI(_11200_),
    .CO(_00200_),
    .S(_11201_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22384_ (.A(_00201_),
    .B(_11201_),
    .CI(_11179_),
    .CO(_00202_),
    .S(_11202_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22385_ (.A(_11181_),
    .B(_11198_),
    .CI(_11202_),
    .CO(_11203_),
    .S(_11204_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22386_ (.A(_00203_),
    .B(_11186_),
    .CI(_11204_),
    .CO(_00204_),
    .S(_00205_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22387_ (.A(_00206_),
    .B(_00207_),
    .CI(_00208_),
    .CO(_11205_),
    .S(_11206_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22388_ (.A(_00209_),
    .B(_00210_),
    .CI(_00211_),
    .CO(_00212_),
    .S(_00213_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22389_ (.A(_00214_),
    .B(_11190_),
    .CI(_11206_),
    .CO(_11207_),
    .S(_11208_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22390_ (.A(_00215_),
    .B(_00216_),
    .CI(_00217_),
    .CO(_11209_),
    .S(_11210_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22391_ (.A(_11194_),
    .B(_11210_),
    .CI(_00218_),
    .CO(_00219_),
    .S(_11211_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22392_ (.A(_11211_),
    .B(_11192_),
    .CI(_11208_),
    .CO(_11212_),
    .S(_11213_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22393_ (.A(_00220_),
    .B(_00221_),
    .CI(_00222_),
    .CO(_11214_),
    .S(_11215_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22394_ (.A(_00223_),
    .B(_00224_),
    .CI(_00225_),
    .CO(_11216_),
    .S(_00226_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22395_ (.A(_11199_),
    .B(_11215_),
    .CI(_00227_),
    .CO(_00228_),
    .S(_00229_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22396_ (.A(_00230_),
    .B(_00231_),
    .CI(_00232_),
    .CO(_11217_),
    .S(_00233_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22397_ (.A(_11197_),
    .B(_11213_),
    .CI(_00234_),
    .CO(_11218_),
    .S(_11219_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22398_ (.A(_00235_),
    .B(_11203_),
    .CI(_11219_),
    .CO(_00236_),
    .S(_00237_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22399_ (.A(_00238_),
    .B(_00239_),
    .CI(_00240_),
    .CO(_11220_),
    .S(_11221_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22400_ (.A(_00241_),
    .B(_00242_),
    .CI(_00243_),
    .CO(_11222_),
    .S(_11223_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22401_ (.A(_11223_),
    .B(_11205_),
    .CI(_11221_),
    .CO(_11224_),
    .S(_11225_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22402_ (.A(_00244_),
    .B(_00245_),
    .CI(_00246_),
    .CO(_11226_),
    .S(_11227_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22403_ (.A(_11209_),
    .B(_11227_),
    .CI(_00247_),
    .CO(_11228_),
    .S(_11229_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22404_ (.A(_11229_),
    .B(_11207_),
    .CI(_11225_),
    .CO(_11230_),
    .S(_11231_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22405_ (.A(_00248_),
    .B(_00249_),
    .CI(_00250_),
    .CO(_11232_),
    .S(_11233_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22406_ (.A(_00253_),
    .B(_00252_),
    .CI(_00251_),
    .CO(_11234_),
    .S(_00254_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22407_ (.A(_00255_),
    .B(_11214_),
    .CI(_11233_),
    .CO(_11235_),
    .S(_00256_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22408_ (.A(_00257_),
    .B(_00258_),
    .CI(_00259_),
    .CO(_11236_),
    .S(_00260_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22409_ (.A(_11231_),
    .B(_00261_),
    .CI(_11212_),
    .CO(_11237_),
    .S(_11238_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22410_ (.A(_00262_),
    .B(_11218_),
    .CI(_11238_),
    .CO(_00263_),
    .S(_00264_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22411_ (.A(_11239_),
    .B(_00265_),
    .CI(_00266_),
    .CO(_11240_),
    .S(_11241_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22412_ (.A(_00267_),
    .B(_00268_),
    .CI(_00269_),
    .CO(_11242_),
    .S(_11243_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22413_ (.A(_00270_),
    .B(_00271_),
    .CI(_00272_),
    .CO(_00273_),
    .S(_00274_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22414_ (.A(_11220_),
    .B(_11243_),
    .CI(_00275_),
    .CO(_11244_),
    .S(_11245_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22415_ (.A(_00276_),
    .B(_00277_),
    .CI(_00278_),
    .CO(_11246_),
    .S(_11247_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22416_ (.A(_11226_),
    .B(_11247_),
    .CI(_11222_),
    .CO(_11248_),
    .S(_11249_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22417_ (.A(_11249_),
    .B(_11224_),
    .CI(_11245_),
    .CO(_11250_),
    .S(_11251_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22418_ (.A(_00279_),
    .B(_00280_),
    .CI(_00281_),
    .CO(_11252_),
    .S(_11253_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22419_ (.A(_00282_),
    .B(_00283_),
    .CI(_00284_),
    .CO(_11254_),
    .S(_00285_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22420_ (.A(_11253_),
    .B(_11232_),
    .CI(_00286_),
    .CO(_11255_),
    .S(_11256_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22421_ (.A(_11256_),
    .B(_11235_),
    .CI(_11228_),
    .CO(_00287_),
    .S(_11257_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22422_ (.A(_11251_),
    .B(_11230_),
    .CI(_11257_),
    .CO(_11258_),
    .S(_11259_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22423_ (.A(_11259_),
    .B(_11237_),
    .CI(_00288_),
    .CO(_00289_),
    .S(_00290_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22424_ (.A(_00292_),
    .B(_00291_),
    .CI(_11260_),
    .CO(_11261_),
    .S(_11262_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22425_ (.A(net1575),
    .B(_09894_),
    .CI(_00295_),
    .CO(_00296_),
    .S(_00297_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22426_ (.A(_00298_),
    .B(_00299_),
    .CI(_00300_),
    .CO(_00301_),
    .S(_00302_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22427_ (.A(_00303_),
    .B(_11242_),
    .CI(_00304_),
    .CO(_11263_),
    .S(_11264_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22428_ (.A(_00305_),
    .B(_00306_),
    .CI(_00307_),
    .CO(_11265_),
    .S(_11266_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22429_ (.A(_11246_),
    .B(_11266_),
    .CI(_00308_),
    .CO(_11267_),
    .S(_11268_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22430_ (.A(_11268_),
    .B(_11244_),
    .CI(_11264_),
    .CO(_11269_),
    .S(_11270_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22431_ (.A(_00309_),
    .B(_00310_),
    .CI(_00311_),
    .CO(_11271_),
    .S(_11272_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22432_ (.A(_00312_),
    .B(_00313_),
    .CI(_00314_),
    .CO(_00315_),
    .S(_00316_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22433_ (.A(_00317_),
    .B(_11252_),
    .CI(_11272_),
    .CO(_11273_),
    .S(_11274_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22434_ (.A(_11255_),
    .B(_11274_),
    .CI(_11248_),
    .CO(_11275_),
    .S(_11276_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22435_ (.A(_11276_),
    .B(_11250_),
    .CI(_11270_),
    .CO(_11277_),
    .S(_11278_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22436_ (.A(_00318_),
    .B(_00319_),
    .CI(_00320_),
    .CO(_11279_),
    .S(_00321_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22437_ (.A(_11280_),
    .B(_00322_),
    .CI(_11254_),
    .CO(_11281_),
    .S(_00323_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22438_ (.A(_00324_),
    .B(_00325_),
    .CI(_00326_),
    .CO(_11282_),
    .S(_00327_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22439_ (.A(_11283_),
    .B(_00328_),
    .CI(_00329_),
    .CO(_00330_),
    .S(_00331_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22440_ (.A(_00332_),
    .B(_11258_),
    .CI(_11278_),
    .CO(_11284_),
    .S(_00333_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22441_ (.A(_11285_),
    .B(_00334_),
    .CI(_00335_),
    .CO(_11286_),
    .S(_11287_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22442_ (.A(net1570),
    .B(_00337_),
    .CI(net1575),
    .CO(_00338_),
    .S(_00339_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22443_ (.A(_00340_),
    .B(_00341_),
    .CI(_00342_),
    .CO(_00343_),
    .S(_00344_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22444_ (.A(_00347_),
    .B(_00346_),
    .CI(_00345_),
    .CO(_11288_),
    .S(_11289_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22445_ (.A(_00348_),
    .B(_00349_),
    .CI(_00350_),
    .CO(_11290_),
    .S(_11291_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22446_ (.A(_11265_),
    .B(_11291_),
    .CI(_00351_),
    .CO(_11292_),
    .S(_11293_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22447_ (.A(_11289_),
    .B(_11263_),
    .CI(_11293_),
    .CO(_11294_),
    .S(_11295_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22448_ (.A(_00352_),
    .B(_00353_),
    .CI(_00354_),
    .CO(_11296_),
    .S(_11297_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22449_ (.A(_00355_),
    .B(_00356_),
    .CI(_00357_),
    .CO(_00358_),
    .S(_00359_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22450_ (.A(_00360_),
    .B(_11271_),
    .CI(_11297_),
    .CO(_11298_),
    .S(_11299_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22451_ (.A(_11273_),
    .B(_11299_),
    .CI(_11267_),
    .CO(_00361_),
    .S(_11300_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22452_ (.A(_11295_),
    .B(_11269_),
    .CI(_11300_),
    .CO(_11301_),
    .S(_11302_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22453_ (.A(_00362_),
    .B(_00363_),
    .CI(_00364_),
    .CO(_11303_),
    .S(_11304_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22454_ (.A(_11279_),
    .B(_11304_),
    .CI(_00365_),
    .CO(_00366_),
    .S(_00367_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22455_ (.A(_11282_),
    .B(_00368_),
    .CI(_11275_),
    .CO(_11305_),
    .S(_11306_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22456_ (.A(_11306_),
    .B(_11277_),
    .CI(_11302_),
    .CO(_11307_),
    .S(_11308_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22457_ (.A(_00369_),
    .B(_11284_),
    .CI(_11308_),
    .CO(_00370_),
    .S(_00371_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22458_ (.A(net1570),
    .B(_00372_),
    .CI(net1575),
    .CO(_00373_),
    .S(_00374_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22459_ (.A(_00375_),
    .B(_00376_),
    .CI(_00377_),
    .CO(_00378_),
    .S(_00379_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22460_ (.A(_00380_),
    .B(_00381_),
    .CI(_00382_),
    .CO(_11309_),
    .S(_11310_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22461_ (.A(_00383_),
    .B(_00384_),
    .CI(_00385_),
    .CO(_11311_),
    .S(_11312_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22462_ (.A(_11290_),
    .B(_11312_),
    .CI(_00386_),
    .CO(_11313_),
    .S(_11314_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22463_ (.A(_11314_),
    .B(_11288_),
    .CI(_11310_),
    .CO(_11315_),
    .S(_11316_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22464_ (.A(_00387_),
    .B(_00388_),
    .CI(_00389_),
    .CO(_11317_),
    .S(_11318_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22465_ (.A(_00390_),
    .B(_00391_),
    .CI(_00392_),
    .CO(_00393_),
    .S(_00394_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22466_ (.A(_00395_),
    .B(_11296_),
    .CI(_11318_),
    .CO(_11319_),
    .S(_11320_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22467_ (.A(_11298_),
    .B(_11320_),
    .CI(_11292_),
    .CO(_00396_),
    .S(_11321_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22468_ (.A(_11321_),
    .B(_11294_),
    .CI(_11316_),
    .CO(_11322_),
    .S(_11323_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22469_ (.A(_00397_),
    .B(_00398_),
    .CI(_00399_),
    .CO(_11324_),
    .S(_11325_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22470_ (.A(_11303_),
    .B(_11325_),
    .CI(_00400_),
    .CO(_00401_),
    .S(_00402_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22471_ (.A(_11326_),
    .B(_11327_),
    .CI(_00403_),
    .CO(_00404_),
    .S(_00405_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22472_ (.A(_00406_),
    .B(_11301_),
    .CI(_11323_),
    .CO(_11328_),
    .S(_11329_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22473_ (.A(_11329_),
    .B(_11305_),
    .CI(_11307_),
    .CO(_00407_),
    .S(_00408_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22474_ (.A(net1570),
    .B(_00409_),
    .CI(net1575),
    .CO(_11330_),
    .S(_00410_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22475_ (.A(_00411_),
    .B(net1569),
    .CI(_00377_),
    .CO(_00413_),
    .S(_00414_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22476_ (.A(_00417_),
    .B(_00416_),
    .CI(_00415_),
    .CO(_11331_),
    .S(_11332_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22477_ (.A(_00418_),
    .B(_00419_),
    .CI(_00420_),
    .CO(_11333_),
    .S(_11334_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22478_ (.A(_11311_),
    .B(_11334_),
    .CI(_00421_),
    .CO(_11335_),
    .S(_11336_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22479_ (.A(_11332_),
    .B(_11309_),
    .CI(_11336_),
    .CO(_11337_),
    .S(_11338_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22480_ (.A(_00422_),
    .B(_00423_),
    .CI(_00424_),
    .CO(_11339_),
    .S(_11340_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22481_ (.A(_00425_),
    .B(_00426_),
    .CI(_00427_),
    .CO(_00428_),
    .S(_00429_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22482_ (.A(_00430_),
    .B(_11317_),
    .CI(_11340_),
    .CO(_11341_),
    .S(_11342_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22483_ (.A(_11342_),
    .B(_11313_),
    .CI(_11319_),
    .CO(_00431_),
    .S(_11343_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22484_ (.A(_11338_),
    .B(_11315_),
    .CI(_11343_),
    .CO(_11344_),
    .S(_11345_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22485_ (.A(_00432_),
    .B(_00433_),
    .CI(_00434_),
    .CO(_11346_),
    .S(_11347_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22486_ (.A(_11324_),
    .B(_11347_),
    .CI(_00435_),
    .CO(_00436_),
    .S(_00437_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22487_ (.A(_11348_),
    .B(_11349_),
    .CI(_00438_),
    .CO(_00439_),
    .S(_00440_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22488_ (.A(_11345_),
    .B(_11322_),
    .CI(_00441_),
    .CO(_11350_),
    .S(_11351_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22489_ (.A(_11351_),
    .B(_11328_),
    .CI(_00442_),
    .CO(_00443_),
    .S(_00444_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22490_ (.A(net1570),
    .B(_00445_),
    .CI(net1575),
    .CO(_00446_),
    .S(_11352_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22491_ (.A(_00377_),
    .B(_00447_),
    .CI(_00412_),
    .CO(_00448_),
    .S(_00449_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22492_ (.A(_11352_),
    .B(_11330_),
    .CI(_00449_),
    .CO(_00450_),
    .S(_00451_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22493_ (.A(_00453_),
    .B(_00454_),
    .CI(_00455_),
    .CO(_11353_),
    .S(_11354_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22494_ (.A(_00456_),
    .B(_11333_),
    .CI(_11354_),
    .CO(_11355_),
    .S(_11356_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22495_ (.A(_11331_),
    .B(_00457_),
    .CI(_11356_),
    .CO(_11357_),
    .S(_11358_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22496_ (.A(_00458_),
    .B(_00459_),
    .CI(_00460_),
    .CO(_11359_),
    .S(_11360_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22497_ (.A(_00461_),
    .B(_00462_),
    .CI(_00463_),
    .CO(_00464_),
    .S(_00465_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22498_ (.A(_00466_),
    .B(_11339_),
    .CI(_11360_),
    .CO(_11361_),
    .S(_11362_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22499_ (.A(_11341_),
    .B(_11362_),
    .CI(_11335_),
    .CO(_00467_),
    .S(_11363_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22500_ (.A(_11363_),
    .B(_11337_),
    .CI(_11358_),
    .CO(_11364_),
    .S(_11365_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22501_ (.A(_00468_),
    .B(_00469_),
    .CI(_00470_),
    .CO(_11366_),
    .S(_11367_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22502_ (.A(_11346_),
    .B(_11367_),
    .CI(_00471_),
    .CO(_00472_),
    .S(_00473_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22503_ (.A(_11368_),
    .B(_11369_),
    .CI(_00474_),
    .CO(_00475_),
    .S(_00476_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22504_ (.A(_00477_),
    .B(_11344_),
    .CI(_11365_),
    .CO(_11370_),
    .S(_11371_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22505_ (.A(_00478_),
    .B(_11350_),
    .CI(_11371_),
    .CO(_00479_),
    .S(_00480_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22506_ (.A(net1571),
    .B(_00481_),
    .CI(net1575),
    .CO(_11372_),
    .S(_00482_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22507_ (.A(_00483_),
    .B(_00452_),
    .CI(_00484_),
    .CO(_11373_),
    .S(_11374_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22508_ (.A(_00485_),
    .B(net1568),
    .CI(_00487_),
    .CO(_00488_),
    .S(_00489_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22509_ (.A(net1545),
    .B(_11353_),
    .CI(_00491_),
    .CO(_11375_),
    .S(_11376_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22510_ (.A(_00492_),
    .B(_11374_),
    .CI(_11376_),
    .CO(_11377_),
    .S(_11378_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22511_ (.A(_00493_),
    .B(_00494_),
    .CI(_00495_),
    .CO(_11379_),
    .S(_11380_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22512_ (.A(_00496_),
    .B(_00497_),
    .CI(_00498_),
    .CO(_00499_),
    .S(_00500_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22513_ (.A(_00501_),
    .B(_11359_),
    .CI(_11380_),
    .CO(_11381_),
    .S(_11382_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22514_ (.A(_11361_),
    .B(_11382_),
    .CI(_11355_),
    .CO(_00502_),
    .S(_11383_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22515_ (.A(_11383_),
    .B(_11357_),
    .CI(_11378_),
    .CO(_11384_),
    .S(_11385_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22516_ (.A(_00503_),
    .B(_00504_),
    .CI(_00505_),
    .CO(_11386_),
    .S(_11387_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22517_ (.A(_11366_),
    .B(_11387_),
    .CI(_00506_),
    .CO(_00507_),
    .S(_00508_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22518_ (.A(_11388_),
    .B(_11389_),
    .CI(_00509_),
    .CO(_00510_),
    .S(_00511_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22519_ (.A(_00512_),
    .B(_11364_),
    .CI(_11385_),
    .CO(_11390_),
    .S(_11391_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22520_ (.A(_00513_),
    .B(_11370_),
    .CI(_11391_),
    .CO(_00514_),
    .S(_00515_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22521_ (.A(net1571),
    .B(_00516_),
    .CI(net1575),
    .CO(_11392_),
    .S(_11393_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22522_ (.A(net2492),
    .B(_11372_),
    .CI(_11393_),
    .CO(_00517_),
    .S(_00518_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22523_ (.A(net1568),
    .B(_00519_),
    .CI(_00520_),
    .CO(_00521_),
    .S(_00522_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22524_ (.A(net1545),
    .B(_00523_),
    .CI(_00524_),
    .CO(_11394_),
    .S(_11395_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22525_ (.A(_11395_),
    .B(_11373_),
    .CI(_00525_),
    .CO(_11396_),
    .S(_11397_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22526_ (.A(_00526_),
    .B(_00527_),
    .CI(_00528_),
    .CO(_11398_),
    .S(_11399_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22527_ (.A(_00529_),
    .B(_00530_),
    .CI(_00531_),
    .CO(_00532_),
    .S(_00533_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22528_ (.A(_00534_),
    .B(_11379_),
    .CI(_11399_),
    .CO(_11400_),
    .S(_11401_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22529_ (.A(_11375_),
    .B(_11381_),
    .CI(_11401_),
    .CO(_00535_),
    .S(_11402_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22530_ (.A(_11377_),
    .B(_11397_),
    .CI(_11402_),
    .CO(_11403_),
    .S(_11404_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22531_ (.A(_00536_),
    .B(_00537_),
    .CI(_00538_),
    .CO(_11405_),
    .S(_11406_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22532_ (.A(_11386_),
    .B(_11406_),
    .CI(_00539_),
    .CO(_00540_),
    .S(_00541_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22533_ (.A(_11407_),
    .B(_11408_),
    .CI(_00542_),
    .CO(_00543_),
    .S(_00544_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22534_ (.A(_00545_),
    .B(_11384_),
    .CI(_11404_),
    .CO(_11409_),
    .S(_11410_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22535_ (.A(_00546_),
    .B(_11390_),
    .CI(_11410_),
    .CO(_00547_),
    .S(_00548_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22536_ (.A(net1570),
    .B(_00549_),
    .CI(net1575),
    .CO(_11411_),
    .S(_11412_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22537_ (.A(net2492),
    .B(_11392_),
    .CI(_11412_),
    .CO(_11413_),
    .S(_00550_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22538_ (.A(_00486_),
    .B(_00520_),
    .CI(_00551_),
    .CO(_00552_),
    .S(_00553_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22539_ (.A(net1545),
    .B(_00554_),
    .CI(_00555_),
    .CO(_11414_),
    .S(_11415_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22540_ (.A(_00556_),
    .B(_00557_),
    .CI(_11415_),
    .CO(_11416_),
    .S(_11417_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22541_ (.A(_00558_),
    .B(_00559_),
    .CI(_00560_),
    .CO(_11418_),
    .S(_11419_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22542_ (.A(_00561_),
    .B(_00562_),
    .CI(_00563_),
    .CO(_00564_),
    .S(_00565_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22543_ (.A(_00566_),
    .B(_11398_),
    .CI(_11419_),
    .CO(_11420_),
    .S(_11421_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22544_ (.A(_11400_),
    .B(_11421_),
    .CI(_11394_),
    .CO(_00567_),
    .S(_11422_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22545_ (.A(_11422_),
    .B(_11396_),
    .CI(_11417_),
    .CO(_11423_),
    .S(_11424_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22546_ (.A(_00568_),
    .B(_00569_),
    .CI(_00570_),
    .CO(_11425_),
    .S(_11426_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22547_ (.A(_11405_),
    .B(_11426_),
    .CI(_00571_),
    .CO(_00572_),
    .S(_00573_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22548_ (.A(_11427_),
    .B(_11428_),
    .CI(_00574_),
    .CO(_00575_),
    .S(_00576_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22549_ (.A(_00577_),
    .B(_11403_),
    .CI(_11424_),
    .CO(_11429_),
    .S(_11430_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22550_ (.A(_00578_),
    .B(_11409_),
    .CI(_11430_),
    .CO(_00579_),
    .S(_00580_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22551_ (.A(net1570),
    .B(_00581_),
    .CI(net1575),
    .CO(_11431_),
    .S(_11432_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22552_ (.A(net2492),
    .B(_11411_),
    .CI(_11432_),
    .CO(_00582_),
    .S(_11433_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _22553_ (.A(_00490_),
    .B(_00583_),
    .CI(_00555_),
    .CO(_11434_),
    .S(_00584_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22554_ (.A(_00585_),
    .B(_11413_),
    .CI(_11433_),
    .CO(_00586_),
    .S(_00587_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22555_ (.A(_00588_),
    .B(_00589_),
    .CI(_00590_),
    .CO(_00591_),
    .S(_00592_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22556_ (.A(_00593_),
    .B(_00594_),
    .CI(_00595_),
    .CO(_00596_),
    .S(_00597_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22557_ (.A(_00598_),
    .B(_11418_),
    .CI(_00599_),
    .CO(_11435_),
    .S(_11436_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22558_ (.A(_11414_),
    .B(_11420_),
    .CI(_11436_),
    .CO(_00600_),
    .S(_11437_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22559_ (.A(_11416_),
    .B(_00601_),
    .CI(_11437_),
    .CO(_11438_),
    .S(_11439_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22560_ (.A(_00602_),
    .B(_00603_),
    .CI(_00604_),
    .CO(_11440_),
    .S(_11441_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22561_ (.A(_11425_),
    .B(_11441_),
    .CI(_00605_),
    .CO(_00606_),
    .S(_00607_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22562_ (.A(_11442_),
    .B(_11443_),
    .CI(_00608_),
    .CO(_00609_),
    .S(_00610_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22563_ (.A(_00611_),
    .B(_11423_),
    .CI(_11439_),
    .CO(_11444_),
    .S(_11445_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22564_ (.A(_00612_),
    .B(_11429_),
    .CI(_11445_),
    .CO(_00613_),
    .S(_00614_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22565_ (.A(net1572),
    .B(_00615_),
    .CI(net1576),
    .CO(_11446_),
    .S(_11447_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22566_ (.A(net2492),
    .B(_11431_),
    .CI(_11447_),
    .CO(_11448_),
    .S(_00616_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22567_ (.A(_00617_),
    .B(_00618_),
    .CI(net1537),
    .CO(_11449_),
    .S(_11450_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22568_ (.A(net1567),
    .B(_00619_),
    .CI(_00620_),
    .CO(_00621_),
    .S(_00622_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22569_ (.A(_00623_),
    .B(_00624_),
    .CI(_00625_),
    .CO(_00626_),
    .S(_00627_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22570_ (.A(_00628_),
    .B(_00629_),
    .CI(_00630_),
    .CO(_11451_),
    .S(_11452_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22571_ (.A(_11435_),
    .B(_11452_),
    .CI(_11434_),
    .CO(_00631_),
    .S(_11453_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22572_ (.A(_11453_),
    .B(_00632_),
    .CI(_11450_),
    .CO(_11454_),
    .S(_11455_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22573_ (.A(_00633_),
    .B(_00634_),
    .CI(_00635_),
    .CO(_11456_),
    .S(_11457_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22574_ (.A(_11440_),
    .B(_11457_),
    .CI(_00636_),
    .CO(_00637_),
    .S(_00638_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22575_ (.A(_11458_),
    .B(_11459_),
    .CI(_00639_),
    .CO(_00640_),
    .S(_00641_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22576_ (.A(_00642_),
    .B(_11438_),
    .CI(_11455_),
    .CO(_11460_),
    .S(_11461_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22577_ (.A(_00643_),
    .B(_11444_),
    .CI(_11461_),
    .CO(_00644_),
    .S(_00645_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22578_ (.A(net1573),
    .B(_00646_),
    .CI(net1576),
    .CO(_11462_),
    .S(_11463_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22579_ (.A(net1550),
    .B(_11463_),
    .CI(_11446_),
    .CO(_11464_),
    .S(_11465_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22580_ (.A(net1536),
    .B(_11448_),
    .CI(_11465_),
    .CO(_00647_),
    .S(_00648_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22581_ (.A(net1567),
    .B(_00620_),
    .CI(_00649_),
    .CO(_00650_),
    .S(_00651_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22582_ (.A(_00652_),
    .B(_00653_),
    .CI(_00654_),
    .CO(_00655_),
    .S(_00656_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22583_ (.A(_00657_),
    .B(_00658_),
    .CI(_00659_),
    .CO(_11466_),
    .S(_11467_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22584_ (.A(_11434_),
    .B(_11451_),
    .CI(_11467_),
    .CO(_00660_),
    .S(_11468_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22585_ (.A(_11468_),
    .B(_11449_),
    .CI(_00661_),
    .CO(_11469_),
    .S(_11470_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22586_ (.A(_00662_),
    .B(_00663_),
    .CI(_00664_),
    .CO(_11471_),
    .S(_11472_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22587_ (.A(_11456_),
    .B(_11472_),
    .CI(_00665_),
    .CO(_00666_),
    .S(_00667_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22588_ (.A(_11473_),
    .B(_11474_),
    .CI(_00668_),
    .CO(_00669_),
    .S(_00670_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22589_ (.A(_00671_),
    .B(_11454_),
    .CI(_11470_),
    .CO(_11475_),
    .S(_11476_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22590_ (.A(_00672_),
    .B(_11460_),
    .CI(_11476_),
    .CO(_00673_),
    .S(_00674_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22591_ (.A(net1573),
    .B(_00675_),
    .CI(net1576),
    .CO(_11477_),
    .S(_11478_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22592_ (.A(net1550),
    .B(_11462_),
    .CI(_11478_),
    .CO(_11479_),
    .S(_11480_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22593_ (.A(net1536),
    .B(_11464_),
    .CI(_11480_),
    .CO(_00676_),
    .S(_00677_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22594_ (.A(_00678_),
    .B(_00679_),
    .CI(_00680_),
    .CO(_00681_),
    .S(_00682_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22595_ (.A(_00683_),
    .B(_00684_),
    .CI(_00659_),
    .CO(_11481_),
    .S(_11482_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22596_ (.A(_11466_),
    .B(_11482_),
    .CI(net1538),
    .CO(_00685_),
    .S(_11483_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22597_ (.A(_11483_),
    .B(_00686_),
    .CI(_00687_),
    .CO(_11484_),
    .S(_11485_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22598_ (.A(_00688_),
    .B(_00689_),
    .CI(_00690_),
    .CO(_11486_),
    .S(_11487_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22599_ (.A(_11471_),
    .B(_11487_),
    .CI(_00691_),
    .CO(_00692_),
    .S(_00693_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22600_ (.A(_11488_),
    .B(_11489_),
    .CI(_00694_),
    .CO(_00695_),
    .S(_00696_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22601_ (.A(_00697_),
    .B(_11469_),
    .CI(_11485_),
    .CO(_11490_),
    .S(_11491_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22602_ (.A(_00698_),
    .B(_11475_),
    .CI(_11491_),
    .CO(_00699_),
    .S(_00700_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22603_ (.A(net1574),
    .B(net1577),
    .CI(_00701_),
    .CO(_11492_),
    .S(_11493_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22604_ (.A(net1550),
    .B(_11477_),
    .CI(_11493_),
    .CO(_11494_),
    .S(_11495_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22605_ (.A(net1536),
    .B(_11479_),
    .CI(_11495_),
    .CO(_00702_),
    .S(_00703_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22606_ (.A(net1566),
    .B(_00704_),
    .CI(_00705_),
    .CO(_00706_),
    .S(_00707_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22607_ (.A(net1544),
    .B(net1546),
    .CI(_00708_),
    .CO(_11496_),
    .S(_11497_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22608_ (.A(net1538),
    .B(_11481_),
    .CI(_11497_),
    .CO(_00709_),
    .S(_11498_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22609_ (.A(_11498_),
    .B(_00710_),
    .CI(_00711_),
    .CO(_11499_),
    .S(_11500_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22610_ (.A(_00712_),
    .B(_00713_),
    .CI(_00714_),
    .CO(_11501_),
    .S(_11502_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22611_ (.A(_11486_),
    .B(_11502_),
    .CI(_00715_),
    .CO(_00716_),
    .S(_00717_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22612_ (.A(_11503_),
    .B(_11504_),
    .CI(_00718_),
    .CO(_00719_),
    .S(_00720_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22613_ (.A(_00721_),
    .B(_11484_),
    .CI(_11500_),
    .CO(_11505_),
    .S(_11506_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22614_ (.A(_00722_),
    .B(_11490_),
    .CI(_11506_),
    .CO(_00723_),
    .S(_00724_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22615_ (.A(net1574),
    .B(net1577),
    .CI(_00725_),
    .CO(_11507_),
    .S(_11508_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22616_ (.A(net1550),
    .B(_11492_),
    .CI(_11508_),
    .CO(_11509_),
    .S(_11510_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22617_ (.A(net1536),
    .B(_11494_),
    .CI(_11510_),
    .CO(_11511_),
    .S(_00726_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22618_ (.A(net1566),
    .B(_00705_),
    .CI(_00727_),
    .CO(_00728_),
    .S(_00729_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22619_ (.A(net1544),
    .B(net1546),
    .CI(_00730_),
    .CO(_11512_),
    .S(_11513_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22620_ (.A(net1538),
    .B(_11496_),
    .CI(_11513_),
    .CO(_00731_),
    .S(_11514_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22621_ (.A(_11514_),
    .B(_00732_),
    .CI(_00733_),
    .CO(_11515_),
    .S(_11516_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22622_ (.A(_00734_),
    .B(_00735_),
    .CI(_00736_),
    .CO(_11517_),
    .S(_11518_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22623_ (.A(_11501_),
    .B(_11518_),
    .CI(_00737_),
    .CO(_00738_),
    .S(_00739_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22624_ (.A(_11519_),
    .B(_11520_),
    .CI(_00740_),
    .CO(_00741_),
    .S(_00742_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22625_ (.A(_00743_),
    .B(_11499_),
    .CI(_11516_),
    .CO(_11521_),
    .S(_11522_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22626_ (.A(_00744_),
    .B(_11505_),
    .CI(_11522_),
    .CO(_00745_),
    .S(_00746_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22627_ (.A(net1574),
    .B(net1577),
    .CI(_00747_),
    .CO(_11523_),
    .S(_11524_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22628_ (.A(net1550),
    .B(_11507_),
    .CI(_11524_),
    .CO(_11525_),
    .S(_11526_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22629_ (.A(net1536),
    .B(_11509_),
    .CI(_11526_),
    .CO(_00748_),
    .S(_11527_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22630_ (.A(net1538),
    .B(_11513_),
    .CI(_11512_),
    .CO(_00749_),
    .S(_00750_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22631_ (.A(_00751_),
    .B(_11511_),
    .CI(_11527_),
    .CO(_00752_),
    .S(_00753_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22632_ (.A(_00754_),
    .B(_00755_),
    .CI(_00756_),
    .CO(_00757_),
    .S(_00758_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22633_ (.A(_11517_),
    .B(_00759_),
    .CI(_00760_),
    .CO(_00761_),
    .S(_00762_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22634_ (.A(_11528_),
    .B(_11529_),
    .CI(_00763_),
    .CO(_00764_),
    .S(_00765_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22635_ (.A(_00766_),
    .B(_11515_),
    .CI(_00767_),
    .CO(_11530_),
    .S(_11531_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22636_ (.A(_00768_),
    .B(_11521_),
    .CI(_11531_),
    .CO(_00769_),
    .S(_00770_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22637_ (.A(net1574),
    .B(net1577),
    .CI(_00771_),
    .CO(_11532_),
    .S(_11533_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22638_ (.A(net1550),
    .B(_11523_),
    .CI(_11533_),
    .CO(_11534_),
    .S(_11535_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22639_ (.A(net1536),
    .B(_11525_),
    .CI(_11535_),
    .CO(_00772_),
    .S(_00773_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22640_ (.A(_00774_),
    .B(_00775_),
    .CI(_00750_),
    .CO(_11536_),
    .S(_11537_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22641_ (.A(_00776_),
    .B(_00756_),
    .CI(_00777_),
    .CO(_11538_),
    .S(_00778_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22642_ (.A(_00760_),
    .B(_00779_),
    .CI(_00780_),
    .CO(_00781_),
    .S(_00782_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22643_ (.A(_00783_),
    .B(_11539_),
    .CI(_11540_),
    .CO(_00784_),
    .S(_00785_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22644_ (.A(_00786_),
    .B(_11537_),
    .CI(_00787_),
    .CO(_11541_),
    .S(_11542_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22645_ (.A(_00788_),
    .B(_11530_),
    .CI(_11542_),
    .CO(_00789_),
    .S(_00790_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22646_ (.A(net1574),
    .B(net1577),
    .CI(_00791_),
    .CO(_00792_),
    .S(_11543_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22647_ (.A(net1550),
    .B(_11532_),
    .CI(_11543_),
    .CO(_00793_),
    .S(_11544_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22648_ (.A(net1536),
    .B(_11534_),
    .CI(_11544_),
    .CO(_00794_),
    .S(_00795_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22649_ (.A(_00796_),
    .B(_00797_),
    .CI(_00750_),
    .CO(_00798_),
    .S(_11545_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22650_ (.A(_00776_),
    .B(_00799_),
    .CI(_00756_),
    .CO(_00800_),
    .S(_11546_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22651_ (.A(_11538_),
    .B(_11546_),
    .CI(_00728_),
    .CO(_00801_),
    .S(_11547_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22652_ (.A(_00783_),
    .B(_11548_),
    .CI(_11549_),
    .CO(_00802_),
    .S(_00803_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22653_ (.A(_00804_),
    .B(_11536_),
    .CI(_11545_),
    .CO(_00805_),
    .S(_11550_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22654_ (.A(_00806_),
    .B(_11541_),
    .CI(_11550_),
    .CO(_00807_),
    .S(_00808_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _22655_ (.A(_00809_),
    .B(_00810_),
    .CI(_00811_),
    .CO(_00812_),
    .S(_00813_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22656_ (.A(_00814_),
    .B(_00815_),
    .CO(_00816_),
    .S(_00817_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22657_ (.A(_00819_),
    .B(_00818_),
    .CO(_00820_),
    .S(_00821_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22658_ (.A(_00822_),
    .B(_00823_),
    .CO(_00824_),
    .S(_00825_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22659_ (.A(_00826_),
    .B(_00827_),
    .CO(_00828_),
    .S(_00829_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22660_ (.A(_00831_),
    .B(_00830_),
    .CO(_00832_),
    .S(_00833_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22661_ (.A(_00834_),
    .B(_00835_),
    .CO(_00836_),
    .S(_00837_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22662_ (.A(_00838_),
    .B(_00839_),
    .CO(_00840_),
    .S(_00841_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22663_ (.A(_00843_),
    .B(_00842_),
    .CO(_00844_),
    .S(_00845_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22664_ (.A(_00847_),
    .B(_00846_),
    .CO(_00848_),
    .S(_00849_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22665_ (.A(_00850_),
    .B(_00851_),
    .CO(_00852_),
    .S(_00853_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22666_ (.A(_00855_),
    .B(_00854_),
    .CO(_00856_),
    .S(_00857_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22667_ (.A(_00859_),
    .B(_00858_),
    .CO(_00860_),
    .S(_00861_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22668_ (.A(_00862_),
    .B(_00863_),
    .CO(_00864_),
    .S(_00865_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _22669_ (.A(_00866_),
    .B(_00867_),
    .CO(_00868_),
    .S(_00869_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22670_ (.A(_00871_),
    .B(_00870_),
    .CO(_00872_),
    .S(_00873_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22671_ (.A(_00875_),
    .B(_00874_),
    .CO(_00876_),
    .S(_00877_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22672_ (.A(_00879_),
    .B(_00878_),
    .CO(_00880_),
    .S(_00881_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22673_ (.A(_00882_),
    .B(_00883_),
    .CO(_00884_),
    .S(_00885_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22674_ (.A(_00886_),
    .B(_00887_),
    .CO(_00888_),
    .S(_00889_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22675_ (.A(_00890_),
    .B(_00891_),
    .CO(_00892_),
    .S(_00893_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22676_ (.A(_00895_),
    .B(_00894_),
    .CO(_00896_),
    .S(_00897_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22677_ (.A(_00898_),
    .B(_00899_),
    .CO(_00900_),
    .S(_00901_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22678_ (.A(_00903_),
    .B(_00902_),
    .CO(_00904_),
    .S(_00905_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22679_ (.A(_00906_),
    .B(_00907_),
    .CO(_00908_),
    .S(_00909_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22680_ (.A(_00911_),
    .B(_00910_),
    .CO(_00912_),
    .S(_00913_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22681_ (.A(_00914_),
    .B(_00915_),
    .CO(_00916_),
    .S(_00917_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22682_ (.A(_00918_),
    .B(_00919_),
    .CO(_00920_),
    .S(_00921_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22683_ (.A(_00922_),
    .B(_00923_),
    .CO(_00924_),
    .S(_00925_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22684_ (.A(_00926_),
    .B(_00927_),
    .CO(_00928_),
    .S(_00929_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22685_ (.A(_00930_),
    .B(_00931_),
    .CO(_00932_),
    .S(_00933_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22686_ (.A(_00934_),
    .B(_00935_),
    .CO(_00936_),
    .S(_00937_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22687_ (.A(_00938_),
    .B(_00939_),
    .CO(_00940_),
    .S(_00941_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22688_ (.A(_09470_),
    .B(_00943_),
    .CO(_00944_),
    .S(_11551_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22689_ (.A(_08008_),
    .B(_00946_),
    .CO(_00947_),
    .S(_00948_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22690_ (.A(_08008_),
    .B(_00949_),
    .CO(_00950_),
    .S(_11552_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22691_ (.A(_08009_),
    .B(_00946_),
    .CO(_00952_),
    .S(_11553_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22692_ (.A(_00953_),
    .B(_00954_),
    .CO(_00955_),
    .S(_00956_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22693_ (.A(\cs_registers_i.priv_mode_id_o[0] ),
    .B(_00957_),
    .CO(_00958_),
    .S(_00959_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22694_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CO(_00960_),
    .S(_00961_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22695_ (.A(_00962_),
    .B(_00963_),
    .CO(_00964_),
    .S(_00965_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22696_ (.A(_00962_),
    .B(_00963_),
    .CO(_00966_),
    .S(_11554_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22697_ (.A(_00962_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_00967_),
    .S(_11555_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22698_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_00963_),
    .CO(_00968_),
    .S(_11556_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22699_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CO(_00969_),
    .S(_11557_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22700_ (.A(_00970_),
    .B(_00971_),
    .CO(_11558_),
    .S(_00972_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22701_ (.A(_11558_),
    .B(_00973_),
    .CO(_11559_),
    .S(_00974_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22702_ (.A(_11559_),
    .B(_11108_),
    .CO(_11560_),
    .S(_00975_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22703_ (.A(_00976_),
    .B(_00977_),
    .CO(_11115_),
    .S(_00978_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22704_ (.A(_11107_),
    .B(_00979_),
    .CO(_11561_),
    .S(_11562_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22705_ (.A(_11560_),
    .B(_11562_),
    .CO(_11563_),
    .S(_00980_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22706_ (.A(_11117_),
    .B(_11561_),
    .CO(_11564_),
    .S(_11565_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22707_ (.A(_11565_),
    .B(_11563_),
    .CO(_11566_),
    .S(_00981_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22708_ (.A(_11113_),
    .B(_00982_),
    .CO(_11128_),
    .S(_00983_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22709_ (.A(_11116_),
    .B(_00984_),
    .CO(_11567_),
    .S(_11568_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22710_ (.A(_11568_),
    .B(_11564_),
    .CO(_11569_),
    .S(_11570_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22711_ (.A(_11570_),
    .B(_11566_),
    .CO(_11571_),
    .S(_00985_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22712_ (.A(_00986_),
    .B(_00987_),
    .CO(_11136_),
    .S(_11572_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22713_ (.A(_00988_),
    .B(_11572_),
    .CO(_11139_),
    .S(_00989_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22714_ (.A(_11130_),
    .B(_11567_),
    .CO(_11573_),
    .S(_11574_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22715_ (.A(_11569_),
    .B(_11574_),
    .CO(_00990_),
    .S(_11575_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22716_ (.A(_11571_),
    .B(_11575_),
    .CO(_00991_),
    .S(_00992_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22717_ (.A(_11141_),
    .B(_11129_),
    .CO(_11576_),
    .S(_11577_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22718_ (.A(_11577_),
    .B(_11573_),
    .CO(_11578_),
    .S(_00993_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22719_ (.A(_00990_),
    .B(_00993_),
    .CO(_00994_),
    .S(_00995_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22720_ (.A(_00996_),
    .B(_11137_),
    .CO(_11158_),
    .S(_00997_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22721_ (.A(_11140_),
    .B(_00998_),
    .CO(_11579_),
    .S(_11580_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22722_ (.A(_11576_),
    .B(_11580_),
    .CO(_11581_),
    .S(_11582_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22723_ (.A(_11578_),
    .B(_11582_),
    .CO(_00999_),
    .S(_01000_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22724_ (.A(_01001_),
    .B(_01002_),
    .CO(_11583_),
    .S(_11584_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22725_ (.A(_11584_),
    .B(_11147_),
    .CO(_11170_),
    .S(_01003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22726_ (.A(_11160_),
    .B(_11579_),
    .CO(_11585_),
    .S(_11586_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22727_ (.A(_11581_),
    .B(_11586_),
    .CO(_01004_),
    .S(_01005_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22728_ (.A(_11583_),
    .B(_01006_),
    .CO(_11185_),
    .S(_11587_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22729_ (.A(_11587_),
    .B(_11155_),
    .CO(_11187_),
    .S(_01007_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22730_ (.A(_11159_),
    .B(_11172_),
    .CO(_11588_),
    .S(_11589_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22731_ (.A(_11585_),
    .B(_11589_),
    .CO(_01008_),
    .S(_01009_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22732_ (.A(_11171_),
    .B(_11189_),
    .CO(_11590_),
    .S(_11591_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22733_ (.A(_11588_),
    .B(_11591_),
    .CO(_01010_),
    .S(_01011_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22734_ (.A(_01012_),
    .B(_01013_),
    .CO(_11592_),
    .S(_01014_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22735_ (.A(_11188_),
    .B(_01015_),
    .CO(_11593_),
    .S(_11594_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22736_ (.A(_11590_),
    .B(_11594_),
    .CO(_01016_),
    .S(_01017_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22737_ (.A(_11592_),
    .B(_01018_),
    .CO(_11239_),
    .S(_01019_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22738_ (.A(_01020_),
    .B(_01021_),
    .CO(_11595_),
    .S(_11596_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22739_ (.A(_11593_),
    .B(_11596_),
    .CO(_01022_),
    .S(_01023_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22740_ (.A(_01024_),
    .B(_11216_),
    .CO(_11597_),
    .S(_11598_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22741_ (.A(_11598_),
    .B(_11217_),
    .CO(_11260_),
    .S(_01025_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22742_ (.A(_11595_),
    .B(_11241_),
    .CO(_01026_),
    .S(_01027_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22743_ (.A(_01028_),
    .B(_01029_),
    .CO(_11280_),
    .S(_11599_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22744_ (.A(_11599_),
    .B(_11234_),
    .CO(_01030_),
    .S(_11600_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22745_ (.A(_11597_),
    .B(_11600_),
    .CO(_11283_),
    .S(_11601_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22746_ (.A(_11601_),
    .B(_11236_),
    .CO(_11285_),
    .S(_01031_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22747_ (.A(_11262_),
    .B(_11240_),
    .CO(_01032_),
    .S(_01033_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22748_ (.A(_11261_),
    .B(_11287_),
    .CO(_01034_),
    .S(_01035_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22749_ (.A(_11281_),
    .B(_01036_),
    .CO(_11326_),
    .S(_01037_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22750_ (.A(_01038_),
    .B(_11286_),
    .CO(_01039_),
    .S(_01040_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22751_ (.A(_01041_),
    .B(_01042_),
    .CO(_11348_),
    .S(_11327_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22752_ (.A(_01043_),
    .B(_01044_),
    .CO(_01045_),
    .S(_01046_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22753_ (.A(_01047_),
    .B(_01048_),
    .CO(_11368_),
    .S(_11349_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22754_ (.A(_01049_),
    .B(_01050_),
    .CO(_01051_),
    .S(_01052_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22755_ (.A(_01053_),
    .B(_01054_),
    .CO(_11388_),
    .S(_11369_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22756_ (.A(_01055_),
    .B(_01056_),
    .CO(_01057_),
    .S(_01058_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22757_ (.A(_01059_),
    .B(_01060_),
    .CO(_11407_),
    .S(_11389_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22758_ (.A(_01061_),
    .B(_01062_),
    .CO(_01063_),
    .S(_01064_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22759_ (.A(_01065_),
    .B(_01066_),
    .CO(_11427_),
    .S(_11408_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22760_ (.A(_01067_),
    .B(_01068_),
    .CO(_01069_),
    .S(_01070_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22761_ (.A(_01071_),
    .B(_01072_),
    .CO(_11442_),
    .S(_11428_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22762_ (.A(_01073_),
    .B(_01074_),
    .CO(_01075_),
    .S(_01076_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22763_ (.A(_01077_),
    .B(_01078_),
    .CO(_11458_),
    .S(_11443_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22764_ (.A(_01079_),
    .B(_01080_),
    .CO(_01081_),
    .S(_01082_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22765_ (.A(_01083_),
    .B(_01084_),
    .CO(_11473_),
    .S(_11459_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22766_ (.A(_01085_),
    .B(_01086_),
    .CO(_01087_),
    .S(_01088_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22767_ (.A(_01089_),
    .B(_01090_),
    .CO(_11488_),
    .S(_11474_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22768_ (.A(_01091_),
    .B(_01092_),
    .CO(_01093_),
    .S(_01094_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22769_ (.A(_01095_),
    .B(_01096_),
    .CO(_11503_),
    .S(_11489_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22770_ (.A(_01097_),
    .B(_01098_),
    .CO(_01099_),
    .S(_01100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22771_ (.A(_01101_),
    .B(_01102_),
    .CO(_11519_),
    .S(_11504_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22772_ (.A(_01103_),
    .B(_01104_),
    .CO(_01105_),
    .S(_01106_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22773_ (.A(_01107_),
    .B(_01108_),
    .CO(_11528_),
    .S(_11520_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22774_ (.A(_01109_),
    .B(_01110_),
    .CO(_01111_),
    .S(_01112_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22775_ (.A(_01113_),
    .B(_01114_),
    .CO(_11539_),
    .S(_11529_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22776_ (.A(_01115_),
    .B(_01116_),
    .CO(_01117_),
    .S(_01118_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22777_ (.A(_01119_),
    .B(_01120_),
    .CO(_11548_),
    .S(_11540_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22778_ (.A(_01121_),
    .B(_01122_),
    .CO(_01123_),
    .S(_01124_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22779_ (.A(_11546_),
    .B(_00728_),
    .CO(_11602_),
    .S(_01125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22780_ (.A(_01126_),
    .B(_11547_),
    .CO(_01127_),
    .S(_11549_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22781_ (.A(_01128_),
    .B(_01129_),
    .CO(_01130_),
    .S(_01131_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22782_ (.A(\cs_registers_i.pc_if_i[2] ),
    .B(_01132_),
    .CO(_01133_),
    .S(_01134_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22783_ (.A(net2289),
    .B(net1703),
    .CO(_01137_),
    .S(_01138_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22784_ (.A(_01139_),
    .B(net1612),
    .CO(_01141_),
    .S(_01142_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22785_ (.A(_01143_),
    .B(net1703),
    .CO(_01144_),
    .S(_11603_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22786_ (.A(_01145_),
    .B(net1586),
    .CO(_01147_),
    .S(_01148_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22787_ (.A(_01149_),
    .B(net2289),
    .CO(_01150_),
    .S(_11604_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22788_ (.A(_01151_),
    .B(net1611),
    .CO(_01153_),
    .S(_01154_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22789_ (.A(_01155_),
    .B(_07773_),
    .CO(_01157_),
    .S(_11605_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22790_ (.A(net2103),
    .B(_01159_),
    .CO(_01160_),
    .S(_01161_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22791_ (.A(_01162_),
    .B(net1702),
    .CO(_01164_),
    .S(_11606_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22792_ (.A(_01165_),
    .B(_01166_),
    .CO(_01167_),
    .S(_01168_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22793_ (.A(_01169_),
    .B(net1701),
    .CO(_01171_),
    .S(_11607_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22794_ (.A(net1692),
    .B(net1700),
    .CO(_01174_),
    .S(_01175_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22795_ (.A(_01176_),
    .B(_07859_),
    .CO(_01178_),
    .S(_11608_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22796_ (.A(net1691),
    .B(_01180_),
    .CO(_01181_),
    .S(_01182_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22797_ (.A(_01183_),
    .B(_01184_),
    .CO(_01185_),
    .S(_11609_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22798_ (.A(net2116),
    .B(_01187_),
    .CO(_01188_),
    .S(_01189_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22799_ (.A(_01190_),
    .B(net2068),
    .CO(_01192_),
    .S(_11610_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22800_ (.A(net2072),
    .B(net1699),
    .CO(_01195_),
    .S(_01196_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22801_ (.A(_01197_),
    .B(_01198_),
    .CO(_01199_),
    .S(_11611_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22802_ (.A(net2097),
    .B(net1698),
    .CO(_01202_),
    .S(_01203_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22803_ (.A(_01204_),
    .B(_01205_),
    .CO(_01206_),
    .S(_11612_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22804_ (.A(net2102),
    .B(net1697),
    .CO(_01209_),
    .S(_01210_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22805_ (.A(_01211_),
    .B(_01212_),
    .CO(_01213_),
    .S(_11613_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22806_ (.A(net2159),
    .B(net1610),
    .CO(_01216_),
    .S(_01217_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22807_ (.A(_01218_),
    .B(net1696),
    .CO(_01220_),
    .S(_11614_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22808_ (.A(_01221_),
    .B(_01222_),
    .CO(_01223_),
    .S(_01224_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22809_ (.A(net2150),
    .B(net1704),
    .CO(_01227_),
    .S(_11615_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22810_ (.A(net2070),
    .B(net2096),
    .CO(_01230_),
    .S(_01231_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22811_ (.A(_01232_),
    .B(_01233_),
    .CO(_01234_),
    .S(_11616_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22812_ (.A(net1685),
    .B(net2176),
    .CO(_01237_),
    .S(_01238_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22813_ (.A(_01239_),
    .B(_01240_),
    .CO(_01241_),
    .S(_11617_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22814_ (.A(net1684),
    .B(_01243_),
    .CO(_01244_),
    .S(_01245_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22815_ (.A(_01246_),
    .B(_01247_),
    .CO(_01248_),
    .S(_11618_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22816_ (.A(net1683),
    .B(_01250_),
    .CO(_01251_),
    .S(_01252_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22817_ (.A(_01253_),
    .B(_01254_),
    .CO(_01255_),
    .S(_11619_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22818_ (.A(_01256_),
    .B(_01257_),
    .CO(_01258_),
    .S(_01259_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22819_ (.A(_01260_),
    .B(_01261_),
    .CO(_01262_),
    .S(_11620_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22820_ (.A(net1682),
    .B(net2482),
    .CO(_01265_),
    .S(_01266_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22821_ (.A(_01267_),
    .B(_01268_),
    .CO(_01269_),
    .S(_11621_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22822_ (.A(net1681),
    .B(_01271_),
    .CO(_01272_),
    .S(_01273_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22823_ (.A(_01274_),
    .B(_01275_),
    .CO(_01276_),
    .S(_11622_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22824_ (.A(net2135),
    .B(_01278_),
    .CO(_01279_),
    .S(_01280_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22825_ (.A(_01281_),
    .B(_01282_),
    .CO(_01283_),
    .S(_11623_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22826_ (.A(net1680),
    .B(_01285_),
    .CO(_01286_),
    .S(_01287_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22827_ (.A(_01288_),
    .B(_01289_),
    .CO(_01290_),
    .S(_11624_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22828_ (.A(net1679),
    .B(_01292_),
    .CO(_01293_),
    .S(_01294_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22829_ (.A(_01295_),
    .B(_01296_),
    .CO(_01297_),
    .S(_11625_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22830_ (.A(net1678),
    .B(_01299_),
    .CO(_01300_),
    .S(_01301_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22831_ (.A(_01302_),
    .B(_01303_),
    .CO(_01304_),
    .S(_11626_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22832_ (.A(net1677),
    .B(_01306_),
    .CO(_01307_),
    .S(_01308_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22833_ (.A(_01309_),
    .B(_01310_),
    .CO(_01311_),
    .S(_11627_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22834_ (.A(_01312_),
    .B(_01313_),
    .CO(_01314_),
    .S(_01315_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22835_ (.A(_01316_),
    .B(_01317_),
    .CO(_01318_),
    .S(_11628_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22836_ (.A(_01319_),
    .B(_01320_),
    .CO(_01321_),
    .S(_01322_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22837_ (.A(_01323_),
    .B(_01324_),
    .CO(_01325_),
    .S(_11629_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22838_ (.A(_01326_),
    .B(_01327_),
    .CO(_01328_),
    .S(_01329_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22839_ (.A(_01330_),
    .B(_01331_),
    .CO(_01332_),
    .S(_11630_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22840_ (.A(net1676),
    .B(_01334_),
    .CO(_01335_),
    .S(_01336_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22841_ (.A(_01337_),
    .B(_01338_),
    .CO(_01339_),
    .S(_11631_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22842_ (.A(net1675),
    .B(_01341_),
    .CO(_01342_),
    .S(_01343_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22843_ (.A(_01344_),
    .B(_01345_),
    .CO(_01346_),
    .S(_11632_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22844_ (.A(_01347_),
    .B(_01348_),
    .CO(_01349_),
    .S(_01350_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22845_ (.A(_01351_),
    .B(_01352_),
    .CO(_01353_),
    .S(_11633_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22846_ (.A(net1885),
    .B(net1520),
    .CO(_01356_),
    .S(_01357_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22847_ (.A(net1539),
    .B(\alu_adder_result_ex[0] ),
    .CO(_01358_),
    .S(_01359_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22848_ (.A(net1539),
    .B(\alu_adder_result_ex[0] ),
    .CO(_01360_),
    .S(_11634_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22849_ (.A(net1539),
    .B(net1540),
    .CO(_01361_),
    .S(_11635_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22850_ (.A(net1539),
    .B(net1540),
    .CO(_01362_),
    .S(_11636_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22851_ (.A(_01363_),
    .B(\alu_adder_result_ex[0] ),
    .CO(_01364_),
    .S(_11637_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _22852_ (.A(_01363_),
    .B(\alu_adder_result_ex[0] ),
    .CO(_01365_),
    .S(_11638_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22853_ (.A(_01363_),
    .B(net1540),
    .CO(_01366_),
    .S(_11639_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22854_ (.A(\cs_registers_i.mhpmcounter[1856] ),
    .B(\cs_registers_i.mhpmcounter[1857] ),
    .CO(_01367_),
    .S(_01368_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22855_ (.A(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ),
    .CO(_01369_),
    .S(_01370_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22856_ (.A(_01371_),
    .B(_01372_),
    .CO(_01373_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _22857_ (.A(_01373_),
    .B(_01374_),
    .CO(_01375_),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22858_ (.D(_01376_),
    .RN(net2037),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.data_type_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22859_ (.D(_01377_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.data_type_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22860_ (.D(_01378_),
    .RN(net2037),
    .CLK(clknet_leaf_29_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22861_ (.D(_01379_),
    .RN(net2037),
    .CLK(clknet_leaf_29_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22862_ (.D(_01380_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 _22863_ (.D(_01381_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 _22864_ (.D(_01382_),
    .SETN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(data_rdata_i[18]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(data_rdata_i[17]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(data_rdata_i[16]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input39 (.I(data_rdata_i[15]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(data_rdata_i[14]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(data_rdata_i[13]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(data_rdata_i[12]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(data_rdata_i[11]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(data_rdata_i[10]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(data_rdata_i[0]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(data_gnt_i),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(data_err_i),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(boot_addr_i[9]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(boot_addr_i[8]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(boot_addr_i[31]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(boot_addr_i[30]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(boot_addr_i[29]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(boot_addr_i[28]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(boot_addr_i[27]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(boot_addr_i[26]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(boot_addr_i[25]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(boot_addr_i[24]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(boot_addr_i[23]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(boot_addr_i[22]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(boot_addr_i[21]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(boot_addr_i[20]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(boot_addr_i[19]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(boot_addr_i[18]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(boot_addr_i[17]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(boot_addr_i[16]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(boot_addr_i[15]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(boot_addr_i[14]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(boot_addr_i[13]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(boot_addr_i[12]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(boot_addr_i[11]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(boot_addr_i[10]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(core_busy_q));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00006_),
    .E(clknet_leaf_2_clk_i_regs),
    .Q(\core_clock_gate_i.en_latch ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_01383_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.mcountinhibit_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_01384_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.mcountinhibit_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_01385_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_01386_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_01387_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_01388_),
    .RN(net2034),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_01389_),
    .RN(net2034),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_01390_),
    .RN(net2034),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_01391_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_01392_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_01393_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_01394_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_01395_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_01396_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_01397_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_01398_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_01399_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_01400_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_01401_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_01402_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_01403_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_01404_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_01405_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_01406_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_01407_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_01408_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_01409_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_01410_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_01411_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_01412_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_01413_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_01414_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_01415_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_01416_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_01417_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_01418_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_01419_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_01420_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_01421_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_01422_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_01423_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_01424_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_01425_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_01426_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_01427_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_01428_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_01429_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_01430_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_01431_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_01432_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_01433_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_01434_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_01435_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_01436_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_01437_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_01438_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_01439_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_01440_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_01441_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_01442_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_01443_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_01444_),
    .RN(net2037),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_01445_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_01446_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_01447_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.mcycle_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_01448_),
    .RN(net2037),
    .CLK(clknet_leaf_23_clk),
    .Q(\cs_registers_i.mcycle_counter_i.counter_val_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[0]$_DFFE_PN0P_  (.D(_01449_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1856] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[10]$_DFFE_PN0P_  (.D(_01450_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1866] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[11]$_DFFE_PN0P_  (.D(_01451_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1867] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[12]$_DFFE_PN0P_  (.D(_01452_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1868] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[13]$_DFFE_PN0P_  (.D(_01453_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1869] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[14]$_DFFE_PN0P_  (.D(_01454_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1870] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[15]$_DFFE_PN0P_  (.D(_01455_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1871] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[16]$_DFFE_PN0P_  (.D(_01456_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1872] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[17]$_DFFE_PN0P_  (.D(_01457_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1873] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[18]$_DFFE_PN0P_  (.D(_01458_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1874] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[19]$_DFFE_PN0P_  (.D(_01459_),
    .RN(net2035),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1875] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[1]$_DFFE_PN0P_  (.D(_01460_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1857] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[20]$_DFFE_PN0P_  (.D(_01461_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mhpmcounter[1876] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[21]$_DFFE_PN0P_  (.D(_01462_),
    .RN(net2035),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1877] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[22]$_DFFE_PN0P_  (.D(_01463_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mhpmcounter[1878] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[23]$_DFFE_PN0P_  (.D(_01464_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mhpmcounter[1879] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[24]$_DFFE_PN0P_  (.D(_01465_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mhpmcounter[1880] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[25]$_DFFE_PN0P_  (.D(_01466_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1881] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[26]$_DFFE_PN0P_  (.D(_01467_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1882] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[27]$_DFFE_PN0P_  (.D(_01468_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1883] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[28]$_DFFE_PN0P_  (.D(_01469_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1884] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[29]$_DFFE_PN0P_  (.D(_01470_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1885] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[2]$_DFFE_PN0P_  (.D(_01471_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1858] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[30]$_DFFE_PN0P_  (.D(_01472_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1886] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[31]$_DFFE_PN0P_  (.D(_01473_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1887] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[32]$_DFFE_PN0P_  (.D(_01474_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1888] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[33]$_DFFE_PN0P_  (.D(_01475_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1889] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[34]$_DFFE_PN0P_  (.D(_01476_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1890] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[35]$_DFFE_PN0P_  (.D(_01477_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1891] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[36]$_DFFE_PN0P_  (.D(_01478_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1892] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[37]$_DFFE_PN0P_  (.D(_01479_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1893] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[38]$_DFFE_PN0P_  (.D(_01480_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1894] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[39]$_DFFE_PN0P_  (.D(_01481_),
    .RN(net2037),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1895] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[3]$_DFFE_PN0P_  (.D(_01482_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1859] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[40]$_DFFE_PN0P_  (.D(_01483_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1896] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[41]$_DFFE_PN0P_  (.D(_01484_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1897] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[42]$_DFFE_PN0P_  (.D(_01485_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1898] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[43]$_DFFE_PN0P_  (.D(_01486_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1899] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[44]$_DFFE_PN0P_  (.D(_01487_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1900] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[45]$_DFFE_PN0P_  (.D(_01488_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1901] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[46]$_DFFE_PN0P_  (.D(_01489_),
    .RN(net2037),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1902] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[47]$_DFFE_PN0P_  (.D(_01490_),
    .RN(net2037),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1903] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[48]$_DFFE_PN0P_  (.D(_01491_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1904] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[49]$_DFFE_PN0P_  (.D(_01492_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1905] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[4]$_DFFE_PN0P_  (.D(_01493_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1860] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[50]$_DFFE_PN0P_  (.D(_01494_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1906] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[51]$_DFFE_PN0P_  (.D(_01495_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1907] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[52]$_DFFE_PN0P_  (.D(_01496_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1908] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[53]$_DFFE_PN0P_  (.D(_01497_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mhpmcounter[1909] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[54]$_DFFE_PN0P_  (.D(_01498_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mhpmcounter[1910] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[55]$_DFFE_PN0P_  (.D(_01499_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mhpmcounter[1911] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[56]$_DFFE_PN0P_  (.D(_01500_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mhpmcounter[1912] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[57]$_DFFE_PN0P_  (.D(_01501_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.mhpmcounter[1913] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[58]$_DFFE_PN0P_  (.D(_01502_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1914] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[59]$_DFFE_PN0P_  (.D(_01503_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1915] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[5]$_DFFE_PN0P_  (.D(_01504_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mhpmcounter[1861] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[60]$_DFFE_PN0P_  (.D(_01505_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1916] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[61]$_DFFE_PN0P_  (.D(_01506_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1917] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[62]$_DFFE_PN0P_  (.D(_01507_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1918] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[63]$_DFFE_PN0P_  (.D(_01508_),
    .RN(net2035),
    .CLK(clknet_leaf_19_clk),
    .Q(\cs_registers_i.mhpmcounter[1919] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[6]$_DFFE_PN0P_  (.D(_01509_),
    .RN(net2034),
    .CLK(clknet_leaf_22_clk),
    .Q(\cs_registers_i.mhpmcounter[1862] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[7]$_DFFE_PN0P_  (.D(_01510_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1863] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[8]$_DFFE_PN0P_  (.D(_01511_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1864] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.minstret_counter_i.counter_val_o[9]$_DFFE_PN0P_  (.D(_01512_),
    .RN(net2034),
    .CLK(clknet_leaf_20_clk),
    .Q(\cs_registers_i.mhpmcounter[1865] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.priv_mode_id_o[0]$_DFFE_PN1P_  (.D(_01513_),
    .SETN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.priv_mode_id_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.priv_mode_id_o[1]$_DFFE_PN1P_  (.D(_01514_),
    .SETN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.priv_mode_id_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[0]$_DFFE_PN1P_  (.D(_01515_),
    .SETN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dcsr_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01516_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dcsr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01517_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dcsr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01518_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dcsr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01519_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dcsr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[1]$_DFFE_PN1P_  (.D(_01520_),
    .SETN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dcsr_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01521_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dcsr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01522_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dcsr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01523_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.dcsr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dcsr_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01524_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dcsr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01525_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_depc_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01526_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.csr_depc_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01527_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_depc_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01528_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01529_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_depc_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01530_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_depc_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01531_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01532_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_depc_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01533_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_depc_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01534_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_depc_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01535_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_depc_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01536_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01537_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01538_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_depc_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01539_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01540_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_depc_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01541_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_depc_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01542_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_depc_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01543_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_depc_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01544_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_depc_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01545_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_depc_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01546_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_depc_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01547_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_depc_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01548_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_depc_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01549_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_depc_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01550_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\cs_registers_i.csr_depc_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01551_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_depc_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01552_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_depc_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01553_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_depc_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01554_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_depc_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_depc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01555_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_depc_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01556_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.dscratch0_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01557_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01558_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.dscratch0_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01559_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.dscratch0_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01560_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch0_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01561_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01562_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch0_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01563_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01564_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dscratch0_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01565_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01566_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01567_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch0_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01568_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01569_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01570_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01571_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01572_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dscratch0_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01573_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01574_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01575_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01576_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01577_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch0_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01578_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01579_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01580_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.dscratch0_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01581_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01582_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.dscratch0_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01583_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.dscratch0_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01584_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01585_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch0_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01586_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch0_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01587_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch0_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01588_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01589_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch1_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01590_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch1_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01591_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch1_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01592_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01593_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01594_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01595_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01596_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01597_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01598_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dscratch1_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01599_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch1_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01600_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01601_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01602_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01603_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01604_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dscratch1_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01605_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01606_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.dscratch1_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01607_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01608_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01609_),
    .RN(net2035),
    .CLK(clknet_leaf_18_clk),
    .Q(\cs_registers_i.dscratch1_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01610_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch1_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01611_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch1_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01612_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch1_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01613_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.dscratch1_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01614_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.dscratch1_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01615_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.dscratch1_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01616_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.dscratch1_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01617_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01618_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_dscratch1_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01619_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.dscratch1_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01620_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mcause_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01621_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mcause_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01622_),
    .RN(net2035),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mcause_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01623_),
    .RN(net2035),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mcause_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01624_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mcause_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mcause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01625_),
    .RN(net2035),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mcause_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01626_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_mepc_o[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01627_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mepc_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01628_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.csr_mepc_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01629_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_mepc_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01630_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_mepc_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01631_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mepc_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01632_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mepc_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01633_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mepc_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01634_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mepc_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01635_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_mepc_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01636_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_mepc_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01637_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_mepc_o[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01638_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_mepc_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01639_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mepc_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01640_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mepc_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01641_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.csr_mepc_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01642_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.csr_mepc_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01643_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mepc_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01644_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mepc_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01645_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mepc_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01646_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mepc_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01647_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mepc_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01648_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mepc_o[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01649_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.csr_mepc_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01650_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mepc_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01651_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mepc_o[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01652_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_mepc_o[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01653_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_mepc_o[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01654_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_mepc_o[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01655_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_mepc_o[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01656_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_mepc_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mepc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01657_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mepc_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01658_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01659_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mie_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01660_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mie_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01661_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mie_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01662_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mie_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01663_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mie_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01664_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mie_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01665_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mie_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01666_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mie_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01667_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01668_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01669_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01670_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01671_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mie_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01672_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01673_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mie_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01674_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mie_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mie_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01675_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mie_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01676_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mscratch_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01677_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mscratch_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01678_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mscratch_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01679_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mscratch_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01680_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mscratch_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01681_),
    .RN(net2035),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mscratch_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01682_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mscratch_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01683_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mscratch_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01684_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mscratch_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01685_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mscratch_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01686_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mscratch_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01687_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mscratch_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01688_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mscratch_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01689_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mscratch_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01690_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mscratch_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01691_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mscratch_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01692_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mscratch_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01693_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mscratch_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01694_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mscratch_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01695_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mscratch_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01696_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mscratch_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01697_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mscratch_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01698_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk),
    .Q(\cs_registers_i.mscratch_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01699_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mscratch_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01700_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mscratch_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01701_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mscratch_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01702_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mscratch_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01703_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\cs_registers_i.mscratch_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01704_),
    .RN(net2034),
    .CLK(clknet_leaf_21_clk),
    .Q(\cs_registers_i.mscratch_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01705_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mscratch_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01706_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mscratch_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mscratch_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01707_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mscratch_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01708_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_cause_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01709_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mstack_cause_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01710_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mstack_cause_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01711_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mstack_cause_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01712_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_cause_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_cause_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01713_),
    .RN(net2035),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_cause_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01714_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstack_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01715_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.u_mstack_csr.rd_data_o[2]$_DFFE_PN1P_  (.D(_01716_),
    .SETN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstack_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01717_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstack_epc_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01718_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mstack_epc_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01719_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mstack_epc_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01720_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_epc_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01721_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mstack_epc_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01722_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mstack_epc_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01723_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mstack_epc_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01724_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mstack_epc_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01725_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mstack_epc_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01726_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mstack_epc_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01727_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mstack_epc_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01728_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_epc_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01729_),
    .RN(net2035),
    .CLK(clknet_leaf_16_clk),
    .Q(\cs_registers_i.mstack_epc_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01730_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mstack_epc_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01731_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mstack_epc_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01732_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mstack_epc_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01733_),
    .RN(net2035),
    .CLK(clknet_leaf_15_clk),
    .Q(\cs_registers_i.mstack_epc_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01734_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mstack_epc_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01735_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.mstack_epc_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01736_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.mstack_epc_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01737_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.mstack_epc_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01738_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mstack_epc_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01739_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mstack_epc_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01740_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstack_epc_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01741_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mstack_epc_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01742_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_epc_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01743_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_epc_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01744_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstack_epc_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01745_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_epc_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01746_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_epc_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01747_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mstack_epc_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstack_epc_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01748_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mstack_epc_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01749_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.csr_mstatus_tw_o ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01750_),
    .RN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstatus_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[2]$_DFFE_PN0N_  (.D(_01751_),
    .RN(net2034),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstatus_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[3]$_DFFE_PN0N_  (.D(_01752_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mstatus_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[4]$_DFFE_PN1N_  (.D(_01753_),
    .SETN(net2035),
    .CLK(clknet_leaf_11_clk),
    .Q(\cs_registers_i.mstatus_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mstatus_csr.rd_data_o[5]$_DFFE_PN0N_  (.D(_01754_),
    .RN(net2035),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.csr_mstatus_mie_o ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[0]$_DFFE_PN0P_  (.D(_01755_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01756_),
    .RN(net2035),
    .CLK(clknet_leaf_9_clk),
    .Q(\cs_registers_i.mtval_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01757_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01758_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01759_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mtval_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01760_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mtval_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01761_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mtval_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01762_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01763_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mtval_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01764_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01765_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[1]$_DFFE_PN0P_  (.D(_01766_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mtval_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01767_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01768_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mtval_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01769_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.mtval_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01770_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.mtval_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01771_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mtval_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01772_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01773_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01774_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01775_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01776_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[2]$_DFFE_PN0P_  (.D(_01777_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01778_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.mtval_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01779_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[3]$_DFFE_PN0P_  (.D(_01780_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[4]$_DFFE_PN0P_  (.D(_01781_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\cs_registers_i.mtval_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[5]$_DFFE_PN0P_  (.D(_01782_),
    .RN(net2034),
    .CLK(clknet_leaf_10_clk),
    .Q(\cs_registers_i.mtval_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[6]$_DFFE_PN0P_  (.D(_01783_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mtval_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[7]$_DFFE_PN0P_  (.D(_01784_),
    .RN(net2035),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.mtval_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01785_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.mtval_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtval_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01786_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.mtval_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[10]$_DFFE_PN0P_  (.D(_01787_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mtvec_o[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[11]$_DFFE_PN0P_  (.D(_01788_),
    .RN(net2035),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.csr_mtvec_o[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[12]$_DFFE_PN0P_  (.D(_01789_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mtvec_o[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[13]$_DFFE_PN0P_  (.D(_01790_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[14]$_DFFE_PN0P_  (.D(_01791_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mtvec_o[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[15]$_DFFE_PN0P_  (.D(_01792_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mtvec_o[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[16]$_DFFE_PN0P_  (.D(_01793_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[17]$_DFFE_PN0P_  (.D(_01794_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mtvec_o[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[18]$_DFFE_PN0P_  (.D(_01795_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[19]$_DFFE_PN0P_  (.D(_01796_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mtvec_o[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[20]$_DFFE_PN0P_  (.D(_01797_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[21]$_DFFE_PN0P_  (.D(_01798_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[22]$_DFFE_PN0P_  (.D(_01799_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mtvec_o[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[23]$_DFFE_PN0P_  (.D(_01800_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[24]$_DFFE_PN0P_  (.D(_01801_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mtvec_o[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[25]$_DFFE_PN0P_  (.D(_01802_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mtvec_o[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[26]$_DFFE_PN0P_  (.D(_01803_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mtvec_o[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[27]$_DFFE_PN0P_  (.D(_01804_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mtvec_o[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[28]$_DFFE_PN0P_  (.D(_01805_),
    .RN(net2035),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.csr_mtvec_o[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[29]$_DFFE_PN0P_  (.D(_01806_),
    .RN(net2035),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.csr_mtvec_o[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[30]$_DFFE_PN0P_  (.D(_01807_),
    .RN(net2035),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.csr_mtvec_o[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[31]$_DFFE_PN0P_  (.D(_01808_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.csr_mtvec_o[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[8]$_DFFE_PN0P_  (.D(_01809_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mtvec_o[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \cs_registers_i.u_mtvec_csr.rd_data_o[9]$_DFFE_PN0P_  (.D(_01810_),
    .RN(net2035),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.csr_mtvec_o[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_01811_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_01812_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_01813_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_01814_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_01815_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_01816_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .SETN(net2037),
    .CLK(clknet_leaf_29_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .RN(net2037),
    .CLK(clknet_leaf_29_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_01817_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_01818_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_01819_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_01820_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_01821_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_01822_),
    .RN(net2037),
    .CLK(clknet_leaf_29_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_01823_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_01824_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_01825_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_01826_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_01827_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_01828_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_01829_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_01830_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_01831_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_01832_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_01833_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_01834_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_01835_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_01836_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_01837_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_01838_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_01839_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_01840_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_01841_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_01842_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_01843_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_01844_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_01845_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_01846_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_01847_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_01848_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_01849_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_01850_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_01851_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_01852_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_01853_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_01854_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_01855_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_01856_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_01857_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_01858_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_01859_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_01860_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_01861_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_01862_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_01863_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_01864_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_01865_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_01866_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_01867_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_01868_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_01869_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_01870_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_01871_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_01872_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_01873_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_01874_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_01875_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_01876_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_01877_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_01878_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_01879_),
    .RN(net2037),
    .CLK(clknet_leaf_27_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_01880_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \fetch_enable_q$_DFFE_PN0P_  (.D(_01881_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(fetch_enable_q));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1000]$_DFFE_PN0P_  (.D(_01882_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1001]$_DFFE_PN0P_  (.D(_01883_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1002]$_DFFE_PN0P_  (.D(_01884_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1003]$_DFFE_PN0P_  (.D(_01885_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1004]$_DFFE_PN0P_  (.D(_01886_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1005]$_DFFE_PN0P_  (.D(_01887_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1006]$_DFFE_PN0P_  (.D(_01888_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1007]$_DFFE_PN0P_  (.D(_01889_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1008]$_DFFE_PN0P_  (.D(_01890_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1009]$_DFFE_PN0P_  (.D(_01891_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[100]$_DFFE_PN0P_  (.D(_01892_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1010]$_DFFE_PN0P_  (.D(_01893_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1011]$_DFFE_PN0P_  (.D(_01894_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1012]$_DFFE_PN0P_  (.D(_01895_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1013]$_DFFE_PN0P_  (.D(_01896_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1014]$_DFFE_PN0P_  (.D(_01897_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1015]$_DFFE_PN0P_  (.D(_01898_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1016]$_DFFE_PN0P_  (.D(_01899_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1017]$_DFFE_PN0P_  (.D(_01900_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1018]$_DFFE_PN0P_  (.D(_01901_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1019]$_DFFE_PN0P_  (.D(_01902_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[101]$_DFFE_PN0P_  (.D(_01903_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1020]$_DFFE_PN0P_  (.D(_01904_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1021]$_DFFE_PN0P_  (.D(_01905_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1022]$_DFFE_PN0P_  (.D(_01906_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[1023]$_DFFE_PN0P_  (.D(_01907_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[102]$_DFFE_PN0P_  (.D(_01908_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[103]$_DFFE_PN0P_  (.D(_01909_),
    .RN(net153),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[104]$_DFFE_PN0P_  (.D(_01910_),
    .RN(net153),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[105]$_DFFE_PN0P_  (.D(_01911_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[106]$_DFFE_PN0P_  (.D(_01912_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[107]$_DFFE_PN0P_  (.D(_01913_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[108]$_DFFE_PN0P_  (.D(_01914_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[109]$_DFFE_PN0P_  (.D(_01915_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[110]$_DFFE_PN0P_  (.D(_01916_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[111]$_DFFE_PN0P_  (.D(_01917_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[112]$_DFFE_PN0P_  (.D(_01918_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[113]$_DFFE_PN0P_  (.D(_01919_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[114]$_DFFE_PN0P_  (.D(_01920_),
    .RN(net2036),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[115]$_DFFE_PN0P_  (.D(_01921_),
    .RN(net2037),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[116]$_DFFE_PN0P_  (.D(_01922_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[117]$_DFFE_PN0P_  (.D(_01923_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[118]$_DFFE_PN0P_  (.D(_01924_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[119]$_DFFE_PN0P_  (.D(_01925_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[120]$_DFFE_PN0P_  (.D(_01926_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[121]$_DFFE_PN0P_  (.D(_01927_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[122]$_DFFE_PN0P_  (.D(_01928_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[123]$_DFFE_PN0P_  (.D(_01929_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[124]$_DFFE_PN0P_  (.D(_01930_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[125]$_DFFE_PN0P_  (.D(_01931_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[126]$_DFFE_PN0P_  (.D(_01932_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[127]$_DFFE_PN0P_  (.D(_01933_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[128]$_DFFE_PN0P_  (.D(_01934_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[129]$_DFFE_PN0P_  (.D(_01935_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[130]$_DFFE_PN0P_  (.D(_01936_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[131]$_DFFE_PN0P_  (.D(_01937_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[132]$_DFFE_PN0P_  (.D(_01938_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[133]$_DFFE_PN0P_  (.D(_01939_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[134]$_DFFE_PN0P_  (.D(_01940_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[135]$_DFFE_PN0P_  (.D(_01941_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[136]$_DFFE_PN0P_  (.D(_01942_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[137]$_DFFE_PN0P_  (.D(_01943_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[138]$_DFFE_PN0P_  (.D(_01944_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[139]$_DFFE_PN0P_  (.D(_01945_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[140]$_DFFE_PN0P_  (.D(_01946_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[141]$_DFFE_PN0P_  (.D(_01947_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[142]$_DFFE_PN0P_  (.D(_01948_),
    .RN(net2033),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[143]$_DFFE_PN0P_  (.D(_01949_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[144]$_DFFE_PN0P_  (.D(_01950_),
    .RN(net153),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[145]$_DFFE_PN0P_  (.D(_01951_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[146]$_DFFE_PN0P_  (.D(_01952_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[147]$_DFFE_PN0P_  (.D(_01953_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[148]$_DFFE_PN0P_  (.D(_01954_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[149]$_DFFE_PN0P_  (.D(_01955_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[150]$_DFFE_PN0P_  (.D(_01956_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[151]$_DFFE_PN0P_  (.D(_01957_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[152]$_DFFE_PN0P_  (.D(_01958_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[153]$_DFFE_PN0P_  (.D(_01959_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[154]$_DFFE_PN0P_  (.D(_01960_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[155]$_DFFE_PN0P_  (.D(_01961_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[156]$_DFFE_PN0P_  (.D(_01962_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[157]$_DFFE_PN0P_  (.D(_01963_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[158]$_DFFE_PN0P_  (.D(_01964_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[159]$_DFFE_PN0P_  (.D(_01965_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[160]$_DFFE_PN0P_  (.D(_01966_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[161]$_DFFE_PN0P_  (.D(_01967_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[162]$_DFFE_PN0P_  (.D(_01968_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[163]$_DFFE_PN0P_  (.D(_01969_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[164]$_DFFE_PN0P_  (.D(_01970_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[165]$_DFFE_PN0P_  (.D(_01971_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[166]$_DFFE_PN0P_  (.D(_01972_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[167]$_DFFE_PN0P_  (.D(_01973_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[168]$_DFFE_PN0P_  (.D(_01974_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[169]$_DFFE_PN0P_  (.D(_01975_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[170]$_DFFE_PN0P_  (.D(_01976_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[171]$_DFFE_PN0P_  (.D(_01977_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[172]$_DFFE_PN0P_  (.D(_01978_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[173]$_DFFE_PN0P_  (.D(_01979_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[174]$_DFFE_PN0P_  (.D(_01980_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[175]$_DFFE_PN0P_  (.D(_01981_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[176]$_DFFE_PN0P_  (.D(_01982_),
    .RN(net153),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[177]$_DFFE_PN0P_  (.D(_01983_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[178]$_DFFE_PN0P_  (.D(_01984_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[179]$_DFFE_PN0P_  (.D(_01985_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[180]$_DFFE_PN0P_  (.D(_01986_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[181]$_DFFE_PN0P_  (.D(_01987_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[182]$_DFFE_PN0P_  (.D(_01988_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[183]$_DFFE_PN0P_  (.D(_01989_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[184]$_DFFE_PN0P_  (.D(_01990_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[185]$_DFFE_PN0P_  (.D(_01991_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[186]$_DFFE_PN0P_  (.D(_01992_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[187]$_DFFE_PN0P_  (.D(_01993_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[188]$_DFFE_PN0P_  (.D(_01994_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[189]$_DFFE_PN0P_  (.D(_01995_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[190]$_DFFE_PN0P_  (.D(_01996_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[191]$_DFFE_PN0P_  (.D(_01997_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[192]$_DFFE_PN0P_  (.D(_01998_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[193]$_DFFE_PN0P_  (.D(_01999_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[194]$_DFFE_PN0P_  (.D(_02000_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[195]$_DFFE_PN0P_  (.D(_02001_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[196]$_DFFE_PN0P_  (.D(_02002_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[197]$_DFFE_PN0P_  (.D(_02003_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[198]$_DFFE_PN0P_  (.D(_02004_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[199]$_DFFE_PN0P_  (.D(_02005_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[200]$_DFFE_PN0P_  (.D(_02006_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[201]$_DFFE_PN0P_  (.D(_02007_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[202]$_DFFE_PN0P_  (.D(_02008_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[203]$_DFFE_PN0P_  (.D(_02009_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[204]$_DFFE_PN0P_  (.D(_02010_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[205]$_DFFE_PN0P_  (.D(_02011_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[206]$_DFFE_PN0P_  (.D(_02012_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[207]$_DFFE_PN0P_  (.D(_02013_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[208]$_DFFE_PN0P_  (.D(_02014_),
    .RN(net153),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[209]$_DFFE_PN0P_  (.D(_02015_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[210]$_DFFE_PN0P_  (.D(_02016_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[211]$_DFFE_PN0P_  (.D(_02017_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[212]$_DFFE_PN0P_  (.D(_02018_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[213]$_DFFE_PN0P_  (.D(_02019_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[214]$_DFFE_PN0P_  (.D(_02020_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[215]$_DFFE_PN0P_  (.D(_02021_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[216]$_DFFE_PN0P_  (.D(_02022_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[217]$_DFFE_PN0P_  (.D(_02023_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[218]$_DFFE_PN0P_  (.D(_02024_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[219]$_DFFE_PN0P_  (.D(_02025_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[220]$_DFFE_PN0P_  (.D(_02026_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[221]$_DFFE_PN0P_  (.D(_02027_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[222]$_DFFE_PN0P_  (.D(_02028_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[223]$_DFFE_PN0P_  (.D(_02029_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[224]$_DFFE_PN0P_  (.D(_02030_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[225]$_DFFE_PN0P_  (.D(_02031_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[226]$_DFFE_PN0P_  (.D(_02032_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[227]$_DFFE_PN0P_  (.D(_02033_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[228]$_DFFE_PN0P_  (.D(_02034_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[229]$_DFFE_PN0P_  (.D(_02035_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[230]$_DFFE_PN0P_  (.D(_02036_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[231]$_DFFE_PN0P_  (.D(_02037_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[232]$_DFFE_PN0P_  (.D(_02038_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[233]$_DFFE_PN0P_  (.D(_02039_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[234]$_DFFE_PN0P_  (.D(_02040_),
    .RN(net2034),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[235]$_DFFE_PN0P_  (.D(_02041_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[236]$_DFFE_PN0P_  (.D(_02042_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[237]$_DFFE_PN0P_  (.D(_02043_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[238]$_DFFE_PN0P_  (.D(_02044_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[239]$_DFFE_PN0P_  (.D(_02045_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[240]$_DFFE_PN0P_  (.D(_02046_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[241]$_DFFE_PN0P_  (.D(_02047_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[242]$_DFFE_PN0P_  (.D(_02048_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[243]$_DFFE_PN0P_  (.D(_02049_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[244]$_DFFE_PN0P_  (.D(_02050_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[245]$_DFFE_PN0P_  (.D(_02051_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[246]$_DFFE_PN0P_  (.D(_02052_),
    .RN(net2034),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[247]$_DFFE_PN0P_  (.D(_02053_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[248]$_DFFE_PN0P_  (.D(_02054_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[249]$_DFFE_PN0P_  (.D(_02055_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[250]$_DFFE_PN0P_  (.D(_02056_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[251]$_DFFE_PN0P_  (.D(_02057_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[252]$_DFFE_PN0P_  (.D(_02058_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[253]$_DFFE_PN0P_  (.D(_02059_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[254]$_DFFE_PN0P_  (.D(_02060_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[255]$_DFFE_PN0P_  (.D(_02061_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[256]$_DFFE_PN0P_  (.D(_02062_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[257]$_DFFE_PN0P_  (.D(_02063_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[258]$_DFFE_PN0P_  (.D(_02064_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[259]$_DFFE_PN0P_  (.D(_02065_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[260]$_DFFE_PN0P_  (.D(_02066_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[261]$_DFFE_PN0P_  (.D(_02067_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[262]$_DFFE_PN0P_  (.D(_02068_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[263]$_DFFE_PN0P_  (.D(_02069_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[264]$_DFFE_PN0P_  (.D(_02070_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[265]$_DFFE_PN0P_  (.D(_02071_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[266]$_DFFE_PN0P_  (.D(_02072_),
    .RN(net2033),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[267]$_DFFE_PN0P_  (.D(_02073_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[268]$_DFFE_PN0P_  (.D(_02074_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[269]$_DFFE_PN0P_  (.D(_02075_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[270]$_DFFE_PN0P_  (.D(_02076_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[271]$_DFFE_PN0P_  (.D(_02077_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[272]$_DFFE_PN0P_  (.D(_02078_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[273]$_DFFE_PN0P_  (.D(_02079_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[274]$_DFFE_PN0P_  (.D(_02080_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[275]$_DFFE_PN0P_  (.D(_02081_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[276]$_DFFE_PN0P_  (.D(_02082_),
    .RN(net2037),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[277]$_DFFE_PN0P_  (.D(_02083_),
    .RN(net153),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[278]$_DFFE_PN0P_  (.D(_02084_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[279]$_DFFE_PN0P_  (.D(_02085_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[280]$_DFFE_PN0P_  (.D(_02086_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[281]$_DFFE_PN0P_  (.D(_02087_),
    .RN(net153),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[282]$_DFFE_PN0P_  (.D(_02088_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[283]$_DFFE_PN0P_  (.D(_02089_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[284]$_DFFE_PN0P_  (.D(_02090_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[285]$_DFFE_PN0P_  (.D(_02091_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[286]$_DFFE_PN0P_  (.D(_02092_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[287]$_DFFE_PN0P_  (.D(_02093_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[288]$_DFFE_PN0P_  (.D(_02094_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[289]$_DFFE_PN0P_  (.D(_02095_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[290]$_DFFE_PN0P_  (.D(_02096_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[291]$_DFFE_PN0P_  (.D(_02097_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[292]$_DFFE_PN0P_  (.D(_02098_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[293]$_DFFE_PN0P_  (.D(_02099_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[294]$_DFFE_PN0P_  (.D(_02100_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[295]$_DFFE_PN0P_  (.D(_02101_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[296]$_DFFE_PN0P_  (.D(_02102_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[297]$_DFFE_PN0P_  (.D(_02103_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[298]$_DFFE_PN0P_  (.D(_02104_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[299]$_DFFE_PN0P_  (.D(_02105_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[300]$_DFFE_PN0P_  (.D(_02106_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[301]$_DFFE_PN0P_  (.D(_02107_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[302]$_DFFE_PN0P_  (.D(_02108_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[303]$_DFFE_PN0P_  (.D(_02109_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[304]$_DFFE_PN0P_  (.D(_02110_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[305]$_DFFE_PN0P_  (.D(_02111_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[306]$_DFFE_PN0P_  (.D(_02112_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[307]$_DFFE_PN0P_  (.D(_02113_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[308]$_DFFE_PN0P_  (.D(_02114_),
    .RN(net2037),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[309]$_DFFE_PN0P_  (.D(_02115_),
    .RN(net153),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[310]$_DFFE_PN0P_  (.D(_02116_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[311]$_DFFE_PN0P_  (.D(_02117_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[312]$_DFFE_PN0P_  (.D(_02118_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[313]$_DFFE_PN0P_  (.D(_02119_),
    .RN(net153),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[314]$_DFFE_PN0P_  (.D(_02120_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[315]$_DFFE_PN0P_  (.D(_02121_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[316]$_DFFE_PN0P_  (.D(_02122_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[317]$_DFFE_PN0P_  (.D(_02123_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[318]$_DFFE_PN0P_  (.D(_02124_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[319]$_DFFE_PN0P_  (.D(_02125_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[320]$_DFFE_PN0P_  (.D(_02126_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[321]$_DFFE_PN0P_  (.D(_02127_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[322]$_DFFE_PN0P_  (.D(_02128_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[323]$_DFFE_PN0P_  (.D(_02129_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[324]$_DFFE_PN0P_  (.D(_02130_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[325]$_DFFE_PN0P_  (.D(_02131_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[326]$_DFFE_PN0P_  (.D(_02132_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[327]$_DFFE_PN0P_  (.D(_02133_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[328]$_DFFE_PN0P_  (.D(_02134_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[329]$_DFFE_PN0P_  (.D(_02135_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[32]$_DFFE_PN0P_  (.D(_02136_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[330]$_DFFE_PN0P_  (.D(_02137_),
    .RN(net2033),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[331]$_DFFE_PN0P_  (.D(_02138_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[332]$_DFFE_PN0P_  (.D(_02139_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[333]$_DFFE_PN0P_  (.D(_02140_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[334]$_DFFE_PN0P_  (.D(_02141_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[335]$_DFFE_PN0P_  (.D(_02142_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[336]$_DFFE_PN0P_  (.D(_02143_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[337]$_DFFE_PN0P_  (.D(_02144_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[338]$_DFFE_PN0P_  (.D(_02145_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[339]$_DFFE_PN0P_  (.D(_02146_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[33]$_DFFE_PN0P_  (.D(_02147_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[340]$_DFFE_PN0P_  (.D(_02148_),
    .RN(net2037),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[341]$_DFFE_PN0P_  (.D(_02149_),
    .RN(net153),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[342]$_DFFE_PN0P_  (.D(_02150_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[343]$_DFFE_PN0P_  (.D(_02151_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[344]$_DFFE_PN0P_  (.D(_02152_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[345]$_DFFE_PN0P_  (.D(_02153_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[346]$_DFFE_PN0P_  (.D(_02154_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[347]$_DFFE_PN0P_  (.D(_02155_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[348]$_DFFE_PN0P_  (.D(_02156_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[349]$_DFFE_PN0P_  (.D(_02157_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[34]$_DFFE_PN0P_  (.D(_02158_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[350]$_DFFE_PN0P_  (.D(_02159_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[351]$_DFFE_PN0P_  (.D(_02160_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[352]$_DFFE_PN0P_  (.D(_02161_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[353]$_DFFE_PN0P_  (.D(_02162_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[354]$_DFFE_PN0P_  (.D(_02163_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[355]$_DFFE_PN0P_  (.D(_02164_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[356]$_DFFE_PN0P_  (.D(_02165_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[357]$_DFFE_PN0P_  (.D(_02166_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[358]$_DFFE_PN0P_  (.D(_02167_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[359]$_DFFE_PN0P_  (.D(_02168_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[35]$_DFFE_PN0P_  (.D(_02169_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[360]$_DFFE_PN0P_  (.D(_02170_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[361]$_DFFE_PN0P_  (.D(_02171_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[362]$_DFFE_PN0P_  (.D(_02172_),
    .RN(net2033),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[363]$_DFFE_PN0P_  (.D(_02173_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[364]$_DFFE_PN0P_  (.D(_02174_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[365]$_DFFE_PN0P_  (.D(_02175_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[366]$_DFFE_PN0P_  (.D(_02176_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[367]$_DFFE_PN0P_  (.D(_02177_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[368]$_DFFE_PN0P_  (.D(_02178_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[369]$_DFFE_PN0P_  (.D(_02179_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[36]$_DFFE_PN0P_  (.D(_02180_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[370]$_DFFE_PN0P_  (.D(_02181_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[371]$_DFFE_PN0P_  (.D(_02182_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[372]$_DFFE_PN0P_  (.D(_02183_),
    .RN(net2037),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[373]$_DFFE_PN0P_  (.D(_02184_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[374]$_DFFE_PN0P_  (.D(_02185_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[375]$_DFFE_PN0P_  (.D(_02186_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[376]$_DFFE_PN0P_  (.D(_02187_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[377]$_DFFE_PN0P_  (.D(_02188_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[378]$_DFFE_PN0P_  (.D(_02189_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[379]$_DFFE_PN0P_  (.D(_02190_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[37]$_DFFE_PN0P_  (.D(_02191_),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[380]$_DFFE_PN0P_  (.D(_02192_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[381]$_DFFE_PN0P_  (.D(_02193_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[382]$_DFFE_PN0P_  (.D(_02194_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[383]$_DFFE_PN0P_  (.D(_02195_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[384]$_DFFE_PN0P_  (.D(_02196_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[385]$_DFFE_PN0P_  (.D(_02197_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[386]$_DFFE_PN0P_  (.D(_02198_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[387]$_DFFE_PN0P_  (.D(_02199_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[388]$_DFFE_PN0P_  (.D(_02200_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[389]$_DFFE_PN0P_  (.D(_02201_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[38]$_DFFE_PN0P_  (.D(_02202_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[390]$_DFFE_PN0P_  (.D(_02203_),
    .RN(net2033),
    .CLK(clknet_leaf_2_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[391]$_DFFE_PN0P_  (.D(_02204_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[392]$_DFFE_PN0P_  (.D(_02205_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[393]$_DFFE_PN0P_  (.D(_02206_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[394]$_DFFE_PN0P_  (.D(_02207_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[395]$_DFFE_PN0P_  (.D(_02208_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[396]$_DFFE_PN0P_  (.D(_02209_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[397]$_DFFE_PN0P_  (.D(_02210_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[398]$_DFFE_PN0P_  (.D(_02211_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[399]$_DFFE_PN0P_  (.D(_02212_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[39]$_DFFE_PN0P_  (.D(_02213_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[400]$_DFFE_PN0P_  (.D(_02214_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[401]$_DFFE_PN0P_  (.D(_02215_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[402]$_DFFE_PN0P_  (.D(_02216_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[403]$_DFFE_PN0P_  (.D(_02217_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[404]$_DFFE_PN0P_  (.D(_02218_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[405]$_DFFE_PN0P_  (.D(_02219_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[406]$_DFFE_PN0P_  (.D(_02220_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[407]$_DFFE_PN0P_  (.D(_02221_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[408]$_DFFE_PN0P_  (.D(_02222_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[409]$_DFFE_PN0P_  (.D(_02223_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[40]$_DFFE_PN0P_  (.D(_02224_),
    .RN(net153),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[410]$_DFFE_PN0P_  (.D(_02225_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[411]$_DFFE_PN0P_  (.D(_02226_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[412]$_DFFE_PN0P_  (.D(_02227_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[413]$_DFFE_PN0P_  (.D(_02228_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[414]$_DFFE_PN0P_  (.D(_02229_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[415]$_DFFE_PN0P_  (.D(_02230_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[416]$_DFFE_PN0P_  (.D(_02231_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[417]$_DFFE_PN0P_  (.D(_02232_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[418]$_DFFE_PN0P_  (.D(_02233_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[419]$_DFFE_PN0P_  (.D(_02234_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[41]$_DFFE_PN0P_  (.D(_02235_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[420]$_DFFE_PN0P_  (.D(_02236_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[421]$_DFFE_PN0P_  (.D(_02237_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[422]$_DFFE_PN0P_  (.D(_02238_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[423]$_DFFE_PN0P_  (.D(_02239_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[424]$_DFFE_PN0P_  (.D(_02240_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[425]$_DFFE_PN0P_  (.D(_02241_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[426]$_DFFE_PN0P_  (.D(_02242_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[427]$_DFFE_PN0P_  (.D(_02243_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[428]$_DFFE_PN0P_  (.D(_02244_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[429]$_DFFE_PN0P_  (.D(_02245_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[42]$_DFFE_PN0P_  (.D(_02246_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[430]$_DFFE_PN0P_  (.D(_02247_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[431]$_DFFE_PN0P_  (.D(_02248_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[432]$_DFFE_PN0P_  (.D(_02249_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[433]$_DFFE_PN0P_  (.D(_02250_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[434]$_DFFE_PN0P_  (.D(_02251_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[435]$_DFFE_PN0P_  (.D(_02252_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[436]$_DFFE_PN0P_  (.D(_02253_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[437]$_DFFE_PN0P_  (.D(_02254_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[438]$_DFFE_PN0P_  (.D(_02255_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[439]$_DFFE_PN0P_  (.D(_02256_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[43]$_DFFE_PN0P_  (.D(_02257_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[440]$_DFFE_PN0P_  (.D(_02258_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[441]$_DFFE_PN0P_  (.D(_02259_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[442]$_DFFE_PN0P_  (.D(_02260_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[443]$_DFFE_PN0P_  (.D(_02261_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[444]$_DFFE_PN0P_  (.D(_02262_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[445]$_DFFE_PN0P_  (.D(_02263_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[446]$_DFFE_PN0P_  (.D(_02264_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[447]$_DFFE_PN0P_  (.D(_02265_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[448]$_DFFE_PN0P_  (.D(_02266_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[449]$_DFFE_PN0P_  (.D(_02267_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[44]$_DFFE_PN0P_  (.D(_02268_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[450]$_DFFE_PN0P_  (.D(_02269_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[451]$_DFFE_PN0P_  (.D(_02270_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[452]$_DFFE_PN0P_  (.D(_02271_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[453]$_DFFE_PN0P_  (.D(_02272_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[454]$_DFFE_PN0P_  (.D(_02273_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[455]$_DFFE_PN0P_  (.D(_02274_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[456]$_DFFE_PN0P_  (.D(_02275_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[457]$_DFFE_PN0P_  (.D(_02276_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[458]$_DFFE_PN0P_  (.D(_02277_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[459]$_DFFE_PN0P_  (.D(_02278_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[45]$_DFFE_PN0P_  (.D(_02279_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[460]$_DFFE_PN0P_  (.D(_02280_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[461]$_DFFE_PN0P_  (.D(_02281_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[462]$_DFFE_PN0P_  (.D(_02282_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[463]$_DFFE_PN0P_  (.D(_02283_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[464]$_DFFE_PN0P_  (.D(_02284_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[465]$_DFFE_PN0P_  (.D(_02285_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[466]$_DFFE_PN0P_  (.D(_02286_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[467]$_DFFE_PN0P_  (.D(_02287_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[468]$_DFFE_PN0P_  (.D(_02288_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[469]$_DFFE_PN0P_  (.D(_02289_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[46]$_DFFE_PN0P_  (.D(_02290_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[470]$_DFFE_PN0P_  (.D(_02291_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[471]$_DFFE_PN0P_  (.D(_02292_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[472]$_DFFE_PN0P_  (.D(_02293_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[473]$_DFFE_PN0P_  (.D(_02294_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[474]$_DFFE_PN0P_  (.D(_02295_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[475]$_DFFE_PN0P_  (.D(_02296_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[476]$_DFFE_PN0P_  (.D(_02297_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[477]$_DFFE_PN0P_  (.D(_02298_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[478]$_DFFE_PN0P_  (.D(_02299_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[479]$_DFFE_PN0P_  (.D(_02300_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[47]$_DFFE_PN0P_  (.D(_02301_),
    .RN(net2033),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[480]$_DFFE_PN0P_  (.D(_02302_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[481]$_DFFE_PN0P_  (.D(_02303_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[482]$_DFFE_PN0P_  (.D(_02304_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[483]$_DFFE_PN0P_  (.D(_02305_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[484]$_DFFE_PN0P_  (.D(_02306_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[485]$_DFFE_PN0P_  (.D(_02307_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[486]$_DFFE_PN0P_  (.D(_02308_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[487]$_DFFE_PN0P_  (.D(_02309_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[488]$_DFFE_PN0P_  (.D(_02310_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[489]$_DFFE_PN0P_  (.D(_02311_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[48]$_DFFE_PN0P_  (.D(_02312_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[490]$_DFFE_PN0P_  (.D(_02313_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[491]$_DFFE_PN0P_  (.D(_02314_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[492]$_DFFE_PN0P_  (.D(_02315_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[493]$_DFFE_PN0P_  (.D(_02316_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[494]$_DFFE_PN0P_  (.D(_02317_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[495]$_DFFE_PN0P_  (.D(_02318_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[496]$_DFFE_PN0P_  (.D(_02319_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[497]$_DFFE_PN0P_  (.D(_02320_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[498]$_DFFE_PN0P_  (.D(_02321_),
    .RN(net2037),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[499]$_DFFE_PN0P_  (.D(_02322_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[49]$_DFFE_PN0P_  (.D(_02323_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[500]$_DFFE_PN0P_  (.D(_02324_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[501]$_DFFE_PN0P_  (.D(_02325_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[502]$_DFFE_PN0P_  (.D(_02326_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[503]$_DFFE_PN0P_  (.D(_02327_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[504]$_DFFE_PN0P_  (.D(_02328_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[505]$_DFFE_PN0P_  (.D(_02329_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[506]$_DFFE_PN0P_  (.D(_02330_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[507]$_DFFE_PN0P_  (.D(_02331_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[508]$_DFFE_PN0P_  (.D(_02332_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[509]$_DFFE_PN0P_  (.D(_02333_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[50]$_DFFE_PN0P_  (.D(_02334_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[510]$_DFFE_PN0P_  (.D(_02335_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[511]$_DFFE_PN0P_  (.D(_02336_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[512]$_DFFE_PN0P_  (.D(_02337_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[513]$_DFFE_PN0P_  (.D(_02338_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[514]$_DFFE_PN0P_  (.D(_02339_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[515]$_DFFE_PN0P_  (.D(_02340_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[516]$_DFFE_PN0P_  (.D(_02341_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[517]$_DFFE_PN0P_  (.D(_02342_),
    .RN(net2034),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[518]$_DFFE_PN0P_  (.D(_02343_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[519]$_DFFE_PN0P_  (.D(_02344_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[51]$_DFFE_PN0P_  (.D(_02345_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[520]$_DFFE_PN0P_  (.D(_02346_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[521]$_DFFE_PN0P_  (.D(_02347_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[522]$_DFFE_PN0P_  (.D(_02348_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[523]$_DFFE_PN0P_  (.D(_02349_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[524]$_DFFE_PN0P_  (.D(_02350_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[525]$_DFFE_PN0P_  (.D(_02351_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[526]$_DFFE_PN0P_  (.D(_02352_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[527]$_DFFE_PN0P_  (.D(_02353_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[528]$_DFFE_PN0P_  (.D(_02354_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[529]$_DFFE_PN0P_  (.D(_02355_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[52]$_DFFE_PN0P_  (.D(_02356_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[530]$_DFFE_PN0P_  (.D(_02357_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[531]$_DFFE_PN0P_  (.D(_02358_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[532]$_DFFE_PN0P_  (.D(_02359_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[533]$_DFFE_PN0P_  (.D(_02360_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[534]$_DFFE_PN0P_  (.D(_02361_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[535]$_DFFE_PN0P_  (.D(_02362_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[536]$_DFFE_PN0P_  (.D(_02363_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[537]$_DFFE_PN0P_  (.D(_02364_),
    .RN(net153),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[538]$_DFFE_PN0P_  (.D(_02365_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[539]$_DFFE_PN0P_  (.D(_02366_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[53]$_DFFE_PN0P_  (.D(_02367_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[540]$_DFFE_PN0P_  (.D(_02368_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[541]$_DFFE_PN0P_  (.D(_02369_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[542]$_DFFE_PN0P_  (.D(_02370_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[543]$_DFFE_PN0P_  (.D(_02371_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[544]$_DFFE_PN0P_  (.D(_02372_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[545]$_DFFE_PN0P_  (.D(_02373_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[546]$_DFFE_PN0P_  (.D(_02374_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[547]$_DFFE_PN0P_  (.D(_02375_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[548]$_DFFE_PN0P_  (.D(_02376_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[549]$_DFFE_PN0P_  (.D(_02377_),
    .RN(net2034),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[54]$_DFFE_PN0P_  (.D(_02378_),
    .RN(net2034),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[550]$_DFFE_PN0P_  (.D(_02379_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[551]$_DFFE_PN0P_  (.D(_02380_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[552]$_DFFE_PN0P_  (.D(_02381_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[553]$_DFFE_PN0P_  (.D(_02382_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[554]$_DFFE_PN0P_  (.D(_02383_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[555]$_DFFE_PN0P_  (.D(_02384_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[556]$_DFFE_PN0P_  (.D(_02385_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[557]$_DFFE_PN0P_  (.D(_02386_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[558]$_DFFE_PN0P_  (.D(_02387_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[559]$_DFFE_PN0P_  (.D(_02388_),
    .RN(net2036),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[55]$_DFFE_PN0P_  (.D(_02389_),
    .RN(net2036),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[560]$_DFFE_PN0P_  (.D(_02390_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[561]$_DFFE_PN0P_  (.D(_02391_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[562]$_DFFE_PN0P_  (.D(_02392_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[563]$_DFFE_PN0P_  (.D(_02393_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[564]$_DFFE_PN0P_  (.D(_02394_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[565]$_DFFE_PN0P_  (.D(_02395_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[566]$_DFFE_PN0P_  (.D(_02396_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[567]$_DFFE_PN0P_  (.D(_02397_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[568]$_DFFE_PN0P_  (.D(_02398_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[569]$_DFFE_PN0P_  (.D(_02399_),
    .RN(net153),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[56]$_DFFE_PN0P_  (.D(_02400_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[570]$_DFFE_PN0P_  (.D(_02401_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[571]$_DFFE_PN0P_  (.D(_02402_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[572]$_DFFE_PN0P_  (.D(_02403_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[573]$_DFFE_PN0P_  (.D(_02404_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[574]$_DFFE_PN0P_  (.D(_02405_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[575]$_DFFE_PN0P_  (.D(_02406_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[576]$_DFFE_PN0P_  (.D(_02407_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[577]$_DFFE_PN0P_  (.D(_02408_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[578]$_DFFE_PN0P_  (.D(_02409_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[579]$_DFFE_PN0P_  (.D(_02410_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[57]$_DFFE_PN0P_  (.D(_02411_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[580]$_DFFE_PN0P_  (.D(_02412_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[581]$_DFFE_PN0P_  (.D(_02413_),
    .RN(net2034),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[582]$_DFFE_PN0P_  (.D(_02414_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[583]$_DFFE_PN0P_  (.D(_02415_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[584]$_DFFE_PN0P_  (.D(_02416_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[585]$_DFFE_PN0P_  (.D(_02417_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[586]$_DFFE_PN0P_  (.D(_02418_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[587]$_DFFE_PN0P_  (.D(_02419_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[588]$_DFFE_PN0P_  (.D(_02420_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[589]$_DFFE_PN0P_  (.D(_02421_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[58]$_DFFE_PN0P_  (.D(_02422_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[590]$_DFFE_PN0P_  (.D(_02423_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[591]$_DFFE_PN0P_  (.D(_02424_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[592]$_DFFE_PN0P_  (.D(_02425_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[593]$_DFFE_PN0P_  (.D(_02426_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[594]$_DFFE_PN0P_  (.D(_02427_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[595]$_DFFE_PN0P_  (.D(_02428_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[596]$_DFFE_PN0P_  (.D(_02429_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[597]$_DFFE_PN0P_  (.D(_02430_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[598]$_DFFE_PN0P_  (.D(_02431_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[599]$_DFFE_PN0P_  (.D(_02432_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[59]$_DFFE_PN0P_  (.D(_02433_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[600]$_DFFE_PN0P_  (.D(_02434_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[601]$_DFFE_PN0P_  (.D(_02435_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[602]$_DFFE_PN0P_  (.D(_02436_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[603]$_DFFE_PN0P_  (.D(_02437_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[604]$_DFFE_PN0P_  (.D(_02438_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[605]$_DFFE_PN0P_  (.D(_02439_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[606]$_DFFE_PN0P_  (.D(_02440_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[607]$_DFFE_PN0P_  (.D(_02441_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[608]$_DFFE_PN0P_  (.D(_02442_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[609]$_DFFE_PN0P_  (.D(_02443_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[60]$_DFFE_PN0P_  (.D(_02444_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[610]$_DFFE_PN0P_  (.D(_02445_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[611]$_DFFE_PN0P_  (.D(_02446_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[612]$_DFFE_PN0P_  (.D(_02447_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[613]$_DFFE_PN0P_  (.D(_02448_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[614]$_DFFE_PN0P_  (.D(_02449_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[615]$_DFFE_PN0P_  (.D(_02450_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[616]$_DFFE_PN0P_  (.D(_02451_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[617]$_DFFE_PN0P_  (.D(_02452_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[618]$_DFFE_PN0P_  (.D(_02453_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[619]$_DFFE_PN0P_  (.D(_02454_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[61]$_DFFE_PN0P_  (.D(_02455_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[620]$_DFFE_PN0P_  (.D(_02456_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[621]$_DFFE_PN0P_  (.D(_02457_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[622]$_DFFE_PN0P_  (.D(_02458_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[623]$_DFFE_PN0P_  (.D(_02459_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[624]$_DFFE_PN0P_  (.D(_02460_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[625]$_DFFE_PN0P_  (.D(_02461_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[626]$_DFFE_PN0P_  (.D(_02462_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[627]$_DFFE_PN0P_  (.D(_02463_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[628]$_DFFE_PN0P_  (.D(_02464_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[629]$_DFFE_PN0P_  (.D(_02465_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[62]$_DFFE_PN0P_  (.D(_02466_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[630]$_DFFE_PN0P_  (.D(_02467_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[631]$_DFFE_PN0P_  (.D(_02468_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[632]$_DFFE_PN0P_  (.D(_02469_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[633]$_DFFE_PN0P_  (.D(_02470_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[634]$_DFFE_PN0P_  (.D(_02471_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[635]$_DFFE_PN0P_  (.D(_02472_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[636]$_DFFE_PN0P_  (.D(_02473_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[637]$_DFFE_PN0P_  (.D(_02474_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[638]$_DFFE_PN0P_  (.D(_02475_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[639]$_DFFE_PN0P_  (.D(_02476_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[63]$_DFFE_PN0P_  (.D(_02477_),
    .RN(net2034),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[640]$_DFFE_PN0P_  (.D(_02478_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[641]$_DFFE_PN0P_  (.D(_02479_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[642]$_DFFE_PN0P_  (.D(_02480_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[643]$_DFFE_PN0P_  (.D(_02481_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[644]$_DFFE_PN0P_  (.D(_02482_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[645]$_DFFE_PN0P_  (.D(_02483_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[646]$_DFFE_PN0P_  (.D(_02484_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[647]$_DFFE_PN0P_  (.D(_02485_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[648]$_DFFE_PN0P_  (.D(_02486_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[649]$_DFFE_PN0P_  (.D(_02487_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[64]$_DFFE_PN0P_  (.D(_02488_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[650]$_DFFE_PN0P_  (.D(_02489_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[651]$_DFFE_PN0P_  (.D(_02490_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[652]$_DFFE_PN0P_  (.D(_02491_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[653]$_DFFE_PN0P_  (.D(_02492_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[654]$_DFFE_PN0P_  (.D(_02493_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[655]$_DFFE_PN0P_  (.D(_02494_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[656]$_DFFE_PN0P_  (.D(_02495_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[657]$_DFFE_PN0P_  (.D(_02496_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[658]$_DFFE_PN0P_  (.D(_02497_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[659]$_DFFE_PN0P_  (.D(_02498_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[65]$_DFFE_PN0P_  (.D(_02499_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[660]$_DFFE_PN0P_  (.D(_02500_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[661]$_DFFE_PN0P_  (.D(_02501_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[662]$_DFFE_PN0P_  (.D(_02502_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[663]$_DFFE_PN0P_  (.D(_02503_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[664]$_DFFE_PN0P_  (.D(_02504_),
    .RN(net2033),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[665]$_DFFE_PN0P_  (.D(_02505_),
    .RN(net153),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[666]$_DFFE_PN0P_  (.D(_02506_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[667]$_DFFE_PN0P_  (.D(_02507_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[668]$_DFFE_PN0P_  (.D(_02508_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[669]$_DFFE_PN0P_  (.D(_02509_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[66]$_DFFE_PN0P_  (.D(_02510_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[670]$_DFFE_PN0P_  (.D(_02511_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[671]$_DFFE_PN0P_  (.D(_02512_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[672]$_DFFE_PN0P_  (.D(_02513_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[673]$_DFFE_PN0P_  (.D(_02514_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[674]$_DFFE_PN0P_  (.D(_02515_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[675]$_DFFE_PN0P_  (.D(_02516_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[676]$_DFFE_PN0P_  (.D(_02517_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[677]$_DFFE_PN0P_  (.D(_02518_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[678]$_DFFE_PN0P_  (.D(_02519_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[679]$_DFFE_PN0P_  (.D(_02520_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[67]$_DFFE_PN0P_  (.D(_02521_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[680]$_DFFE_PN0P_  (.D(_02522_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[681]$_DFFE_PN0P_  (.D(_02523_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[682]$_DFFE_PN0P_  (.D(_02524_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[683]$_DFFE_PN0P_  (.D(_02525_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[684]$_DFFE_PN0P_  (.D(_02526_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[685]$_DFFE_PN0P_  (.D(_02527_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[686]$_DFFE_PN0P_  (.D(_02528_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[687]$_DFFE_PN0P_  (.D(_02529_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[688]$_DFFE_PN0P_  (.D(_02530_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[689]$_DFFE_PN0P_  (.D(_02531_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[68]$_DFFE_PN0P_  (.D(_02532_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[690]$_DFFE_PN0P_  (.D(_02533_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[691]$_DFFE_PN0P_  (.D(_02534_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[692]$_DFFE_PN0P_  (.D(_02535_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[693]$_DFFE_PN0P_  (.D(_02536_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[694]$_DFFE_PN0P_  (.D(_02537_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[695]$_DFFE_PN0P_  (.D(_02538_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[696]$_DFFE_PN0P_  (.D(_02539_),
    .RN(net2033),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[697]$_DFFE_PN0P_  (.D(_02540_),
    .RN(net153),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[698]$_DFFE_PN0P_  (.D(_02541_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[699]$_DFFE_PN0P_  (.D(_02542_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[69]$_DFFE_PN0P_  (.D(_02543_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[700]$_DFFE_PN0P_  (.D(_02544_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[701]$_DFFE_PN0P_  (.D(_02545_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[702]$_DFFE_PN0P_  (.D(_02546_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[703]$_DFFE_PN0P_  (.D(_02547_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[704]$_DFFE_PN0P_  (.D(_02548_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[705]$_DFFE_PN0P_  (.D(_02549_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[706]$_DFFE_PN0P_  (.D(_02550_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[707]$_DFFE_PN0P_  (.D(_02551_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[708]$_DFFE_PN0P_  (.D(_02552_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[709]$_DFFE_PN0P_  (.D(_02553_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[70]$_DFFE_PN0P_  (.D(_02554_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[710]$_DFFE_PN0P_  (.D(_02555_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[711]$_DFFE_PN0P_  (.D(_02556_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[712]$_DFFE_PN0P_  (.D(_02557_),
    .RN(net153),
    .CLK(clknet_leaf_5_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[713]$_DFFE_PN0P_  (.D(_02558_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[714]$_DFFE_PN0P_  (.D(_02559_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[715]$_DFFE_PN0P_  (.D(_02560_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[716]$_DFFE_PN0P_  (.D(_02561_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[717]$_DFFE_PN0P_  (.D(_02562_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[718]$_DFFE_PN0P_  (.D(_02563_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[719]$_DFFE_PN0P_  (.D(_02564_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[71]$_DFFE_PN0P_  (.D(_02565_),
    .RN(net153),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[720]$_DFFE_PN0P_  (.D(_02566_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[721]$_DFFE_PN0P_  (.D(_02567_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[722]$_DFFE_PN0P_  (.D(_02568_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[723]$_DFFE_PN0P_  (.D(_02569_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[724]$_DFFE_PN0P_  (.D(_02570_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[725]$_DFFE_PN0P_  (.D(_02571_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[726]$_DFFE_PN0P_  (.D(_02572_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[727]$_DFFE_PN0P_  (.D(_02573_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[728]$_DFFE_PN0P_  (.D(_02574_),
    .RN(net2033),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[729]$_DFFE_PN0P_  (.D(_02575_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[72]$_DFFE_PN0P_  (.D(_02576_),
    .RN(net153),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[730]$_DFFE_PN0P_  (.D(_02577_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[731]$_DFFE_PN0P_  (.D(_02578_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[732]$_DFFE_PN0P_  (.D(_02579_),
    .RN(net2037),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[733]$_DFFE_PN0P_  (.D(_02580_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[734]$_DFFE_PN0P_  (.D(_02581_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[735]$_DFFE_PN0P_  (.D(_02582_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[736]$_DFFE_PN0P_  (.D(_02583_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[737]$_DFFE_PN0P_  (.D(_02584_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[738]$_DFFE_PN0P_  (.D(_02585_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[739]$_DFFE_PN0P_  (.D(_02586_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[73]$_DFFE_PN0P_  (.D(_02587_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[740]$_DFFE_PN0P_  (.D(_02588_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[741]$_DFFE_PN0P_  (.D(_02589_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[742]$_DFFE_PN0P_  (.D(_02590_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[743]$_DFFE_PN0P_  (.D(_02591_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[744]$_DFFE_PN0P_  (.D(_02592_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[745]$_DFFE_PN0P_  (.D(_02593_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[746]$_DFFE_PN0P_  (.D(_02594_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[747]$_DFFE_PN0P_  (.D(_02595_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[748]$_DFFE_PN0P_  (.D(_02596_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[749]$_DFFE_PN0P_  (.D(_02597_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[74]$_DFFE_PN0P_  (.D(_02598_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[750]$_DFFE_PN0P_  (.D(_02599_),
    .RN(net153),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[751]$_DFFE_PN0P_  (.D(_02600_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[752]$_DFFE_PN0P_  (.D(_02601_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[753]$_DFFE_PN0P_  (.D(_02602_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[754]$_DFFE_PN0P_  (.D(_02603_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[755]$_DFFE_PN0P_  (.D(_02604_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[756]$_DFFE_PN0P_  (.D(_02605_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[757]$_DFFE_PN0P_  (.D(_02606_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[758]$_DFFE_PN0P_  (.D(_02607_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[759]$_DFFE_PN0P_  (.D(_02608_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[75]$_DFFE_PN0P_  (.D(_02609_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[760]$_DFFE_PN0P_  (.D(_02610_),
    .RN(net2033),
    .CLK(clknet_leaf_23_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[761]$_DFFE_PN0P_  (.D(_02611_),
    .RN(net153),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[762]$_DFFE_PN0P_  (.D(_02612_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[763]$_DFFE_PN0P_  (.D(_02613_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[764]$_DFFE_PN0P_  (.D(_02614_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[765]$_DFFE_PN0P_  (.D(_02615_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[766]$_DFFE_PN0P_  (.D(_02616_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[767]$_DFFE_PN0P_  (.D(_02617_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[768]$_DFFE_PN0P_  (.D(_02618_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[769]$_DFFE_PN0P_  (.D(_02619_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[76]$_DFFE_PN0P_  (.D(_02620_),
    .RN(net2033),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[770]$_DFFE_PN0P_  (.D(_02621_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[771]$_DFFE_PN0P_  (.D(_02622_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[772]$_DFFE_PN0P_  (.D(_02623_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[773]$_DFFE_PN0P_  (.D(_02624_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[774]$_DFFE_PN0P_  (.D(_02625_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[775]$_DFFE_PN0P_  (.D(_02626_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[776]$_DFFE_PN0P_  (.D(_02627_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[777]$_DFFE_PN0P_  (.D(_02628_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[778]$_DFFE_PN0P_  (.D(_02629_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[779]$_DFFE_PN0P_  (.D(_02630_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[77]$_DFFE_PN0P_  (.D(_02631_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[780]$_DFFE_PN0P_  (.D(_02632_),
    .RN(net153),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[781]$_DFFE_PN0P_  (.D(_02633_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[782]$_DFFE_PN0P_  (.D(_02634_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[783]$_DFFE_PN0P_  (.D(_02635_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[784]$_DFFE_PN0P_  (.D(_02636_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[785]$_DFFE_PN0P_  (.D(_02637_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[786]$_DFFE_PN0P_  (.D(_02638_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[787]$_DFFE_PN0P_  (.D(_02639_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[788]$_DFFE_PN0P_  (.D(_02640_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[789]$_DFFE_PN0P_  (.D(_02641_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[78]$_DFFE_PN0P_  (.D(_02642_),
    .RN(net2033),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[790]$_DFFE_PN0P_  (.D(_02643_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[791]$_DFFE_PN0P_  (.D(_02644_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[792]$_DFFE_PN0P_  (.D(_02645_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[793]$_DFFE_PN0P_  (.D(_02646_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[794]$_DFFE_PN0P_  (.D(_02647_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[795]$_DFFE_PN0P_  (.D(_02648_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[796]$_DFFE_PN0P_  (.D(_02649_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[797]$_DFFE_PN0P_  (.D(_02650_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[798]$_DFFE_PN0P_  (.D(_02651_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[799]$_DFFE_PN0P_  (.D(_02652_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[79]$_DFFE_PN0P_  (.D(_02653_),
    .RN(net153),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[800]$_DFFE_PN0P_  (.D(_02654_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[801]$_DFFE_PN0P_  (.D(_02655_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[802]$_DFFE_PN0P_  (.D(_02656_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[803]$_DFFE_PN0P_  (.D(_02657_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[804]$_DFFE_PN0P_  (.D(_02658_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[805]$_DFFE_PN0P_  (.D(_02659_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[806]$_DFFE_PN0P_  (.D(_02660_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[807]$_DFFE_PN0P_  (.D(_02661_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[808]$_DFFE_PN0P_  (.D(_02662_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[809]$_DFFE_PN0P_  (.D(_02663_),
    .RN(net2033),
    .CLK(clknet_leaf_25_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[80]$_DFFE_PN0P_  (.D(_02664_),
    .RN(net153),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[810]$_DFFE_PN0P_  (.D(_02665_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[811]$_DFFE_PN0P_  (.D(_02666_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[812]$_DFFE_PN0P_  (.D(_02667_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[813]$_DFFE_PN0P_  (.D(_02668_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[814]$_DFFE_PN0P_  (.D(_02669_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[815]$_DFFE_PN0P_  (.D(_02670_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[816]$_DFFE_PN0P_  (.D(_02671_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[817]$_DFFE_PN0P_  (.D(_02672_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[818]$_DFFE_PN0P_  (.D(_02673_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[819]$_DFFE_PN0P_  (.D(_02674_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[81]$_DFFE_PN0P_  (.D(_02675_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[820]$_DFFE_PN0P_  (.D(_02676_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[821]$_DFFE_PN0P_  (.D(_02677_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[822]$_DFFE_PN0P_  (.D(_02678_),
    .RN(net153),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[823]$_DFFE_PN0P_  (.D(_02679_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[824]$_DFFE_PN0P_  (.D(_02680_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[825]$_DFFE_PN0P_  (.D(_02681_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[826]$_DFFE_PN0P_  (.D(_02682_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[827]$_DFFE_PN0P_  (.D(_02683_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[828]$_DFFE_PN0P_  (.D(_02684_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[829]$_DFFE_PN0P_  (.D(_02685_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[82]$_DFFE_PN0P_  (.D(_02686_),
    .RN(net2037),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[830]$_DFFE_PN0P_  (.D(_02687_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[831]$_DFFE_PN0P_  (.D(_02688_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[832]$_DFFE_PN0P_  (.D(_02689_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[833]$_DFFE_PN0P_  (.D(_02690_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[834]$_DFFE_PN0P_  (.D(_02691_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[835]$_DFFE_PN0P_  (.D(_02692_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[836]$_DFFE_PN0P_  (.D(_02693_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[837]$_DFFE_PN0P_  (.D(_02694_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[838]$_DFFE_PN0P_  (.D(_02695_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[839]$_DFFE_PN0P_  (.D(_02696_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[83]$_DFFE_PN0P_  (.D(_02697_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[840]$_DFFE_PN0P_  (.D(_02698_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[841]$_DFFE_PN0P_  (.D(_02699_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[842]$_DFFE_PN0P_  (.D(_02700_),
    .RN(net2034),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[843]$_DFFE_PN0P_  (.D(_02701_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[844]$_DFFE_PN0P_  (.D(_02702_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[845]$_DFFE_PN0P_  (.D(_02703_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[846]$_DFFE_PN0P_  (.D(_02704_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[847]$_DFFE_PN0P_  (.D(_02705_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[848]$_DFFE_PN0P_  (.D(_02706_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[849]$_DFFE_PN0P_  (.D(_02707_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[84]$_DFFE_PN0P_  (.D(_02708_),
    .RN(net2037),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[850]$_DFFE_PN0P_  (.D(_02709_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[851]$_DFFE_PN0P_  (.D(_02710_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[852]$_DFFE_PN0P_  (.D(_02711_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[853]$_DFFE_PN0P_  (.D(_02712_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[854]$_DFFE_PN0P_  (.D(_02713_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[855]$_DFFE_PN0P_  (.D(_02714_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[856]$_DFFE_PN0P_  (.D(_02715_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[857]$_DFFE_PN0P_  (.D(_02716_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[858]$_DFFE_PN0P_  (.D(_02717_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[859]$_DFFE_PN0P_  (.D(_02718_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[85]$_DFFE_PN0P_  (.D(_02719_),
    .RN(net2033),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[860]$_DFFE_PN0P_  (.D(_02720_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[861]$_DFFE_PN0P_  (.D(_02721_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[862]$_DFFE_PN0P_  (.D(_02722_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[863]$_DFFE_PN0P_  (.D(_02723_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[864]$_DFFE_PN0P_  (.D(_02724_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[865]$_DFFE_PN0P_  (.D(_02725_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[866]$_DFFE_PN0P_  (.D(_02726_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[867]$_DFFE_PN0P_  (.D(_02727_),
    .RN(net2034),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[868]$_DFFE_PN0P_  (.D(_02728_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[869]$_DFFE_PN0P_  (.D(_02729_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[86]$_DFFE_PN0P_  (.D(_02730_),
    .RN(net2034),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[870]$_DFFE_PN0P_  (.D(_02731_),
    .RN(net2033),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[871]$_DFFE_PN0P_  (.D(_02732_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[872]$_DFFE_PN0P_  (.D(_02733_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[873]$_DFFE_PN0P_  (.D(_02734_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[874]$_DFFE_PN0P_  (.D(_02735_),
    .RN(net2034),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[875]$_DFFE_PN0P_  (.D(_02736_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[876]$_DFFE_PN0P_  (.D(_02737_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[877]$_DFFE_PN0P_  (.D(_02738_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[878]$_DFFE_PN0P_  (.D(_02739_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[879]$_DFFE_PN0P_  (.D(_02740_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[87]$_DFFE_PN0P_  (.D(_02741_),
    .RN(net2036),
    .CLK(clknet_leaf_18_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[880]$_DFFE_PN0P_  (.D(_02742_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[881]$_DFFE_PN0P_  (.D(_02743_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[882]$_DFFE_PN0P_  (.D(_02744_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[883]$_DFFE_PN0P_  (.D(_02745_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[884]$_DFFE_PN0P_  (.D(_02746_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[885]$_DFFE_PN0P_  (.D(_02747_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[886]$_DFFE_PN0P_  (.D(_02748_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[887]$_DFFE_PN0P_  (.D(_02749_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[888]$_DFFE_PN0P_  (.D(_02750_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[889]$_DFFE_PN0P_  (.D(_02751_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[88]$_DFFE_PN0P_  (.D(_02752_),
    .RN(net2034),
    .CLK(clknet_leaf_26_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[890]$_DFFE_PN0P_  (.D(_02753_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[891]$_DFFE_PN0P_  (.D(_02754_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[892]$_DFFE_PN0P_  (.D(_02755_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[893]$_DFFE_PN0P_  (.D(_02756_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[894]$_DFFE_PN0P_  (.D(_02757_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[895]$_DFFE_PN0P_  (.D(_02758_),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[896]$_DFFE_PN0P_  (.D(_02759_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[897]$_DFFE_PN0P_  (.D(_02760_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[898]$_DFFE_PN0P_  (.D(_02761_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[899]$_DFFE_PN0P_  (.D(_02762_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[89]$_DFFE_PN0P_  (.D(_02763_),
    .RN(net2037),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[900]$_DFFE_PN0P_  (.D(_02764_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[901]$_DFFE_PN0P_  (.D(_02765_),
    .RN(net2034),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[902]$_DFFE_PN0P_  (.D(_02766_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[903]$_DFFE_PN0P_  (.D(_02767_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[904]$_DFFE_PN0P_  (.D(_02768_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[905]$_DFFE_PN0P_  (.D(_02769_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[906]$_DFFE_PN0P_  (.D(_02770_),
    .RN(net2034),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[907]$_DFFE_PN0P_  (.D(_02771_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[908]$_DFFE_PN0P_  (.D(_02772_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[909]$_DFFE_PN0P_  (.D(_02773_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[90]$_DFFE_PN0P_  (.D(_02774_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[910]$_DFFE_PN0P_  (.D(_02775_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[911]$_DFFE_PN0P_  (.D(_02776_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[912]$_DFFE_PN0P_  (.D(_02777_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[913]$_DFFE_PN0P_  (.D(_02778_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[914]$_DFFE_PN0P_  (.D(_02779_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[915]$_DFFE_PN0P_  (.D(_02780_),
    .RN(net2037),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[916]$_DFFE_PN0P_  (.D(_02781_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[917]$_DFFE_PN0P_  (.D(_02782_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[918]$_DFFE_PN0P_  (.D(_02783_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[919]$_DFFE_PN0P_  (.D(_02784_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[91]$_DFFE_PN0P_  (.D(_02785_),
    .RN(net2036),
    .CLK(clknet_leaf_14_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[920]$_DFFE_PN0P_  (.D(_02786_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[921]$_DFFE_PN0P_  (.D(_02787_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[922]$_DFFE_PN0P_  (.D(_02788_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[923]$_DFFE_PN0P_  (.D(_02789_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[924]$_DFFE_PN0P_  (.D(_02790_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[925]$_DFFE_PN0P_  (.D(_02791_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[926]$_DFFE_PN0P_  (.D(_02792_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[927]$_DFFE_PN0P_  (.D(_02793_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[928]$_DFFE_PN0P_  (.D(_02794_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[929]$_DFFE_PN0P_  (.D(_02795_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[92]$_DFFE_PN0P_  (.D(_02796_),
    .RN(net153),
    .CLK(clknet_leaf_6_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[930]$_DFFE_PN0P_  (.D(_02797_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[931]$_DFFE_PN0P_  (.D(_02798_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[932]$_DFFE_PN0P_  (.D(_02799_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[933]$_DFFE_PN0P_  (.D(_02800_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[934]$_DFFE_PN0P_  (.D(_02801_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[935]$_DFFE_PN0P_  (.D(_02802_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[936]$_DFFE_PN0P_  (.D(_02803_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[937]$_DFFE_PN0P_  (.D(_02804_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[938]$_DFFE_PN0P_  (.D(_02805_),
    .RN(net2034),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[939]$_DFFE_PN0P_  (.D(_02806_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[93]$_DFFE_PN0P_  (.D(_02807_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[940]$_DFFE_PN0P_  (.D(_02808_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[941]$_DFFE_PN0P_  (.D(_02809_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[942]$_DFFE_PN0P_  (.D(_02810_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[943]$_DFFE_PN0P_  (.D(_02811_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[944]$_DFFE_PN0P_  (.D(_02812_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[945]$_DFFE_PN0P_  (.D(_02813_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[946]$_DFFE_PN0P_  (.D(_02814_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[947]$_DFFE_PN0P_  (.D(_02815_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[948]$_DFFE_PN0P_  (.D(_02816_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[949]$_DFFE_PN0P_  (.D(_02817_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[94]$_DFFE_PN0P_  (.D(_02818_),
    .RN(net2036),
    .CLK(clknet_leaf_11_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[950]$_DFFE_PN0P_  (.D(_02819_),
    .RN(net153),
    .CLK(clknet_leaf_17_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[951]$_DFFE_PN0P_  (.D(_02820_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[952]$_DFFE_PN0P_  (.D(_02821_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[953]$_DFFE_PN0P_  (.D(_02822_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[954]$_DFFE_PN0P_  (.D(_02823_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[955]$_DFFE_PN0P_  (.D(_02824_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[956]$_DFFE_PN0P_  (.D(_02825_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[957]$_DFFE_PN0P_  (.D(_02826_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[958]$_DFFE_PN0P_  (.D(_02827_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[959]$_DFFE_PN0P_  (.D(_02828_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[95]$_DFFE_PN0P_  (.D(_02829_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[960]$_DFFE_PN0P_  (.D(_02830_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[961]$_DFFE_PN0P_  (.D(_02831_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[962]$_DFFE_PN0P_  (.D(_02832_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[963]$_DFFE_PN0P_  (.D(_02833_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[964]$_DFFE_PN0P_  (.D(_02834_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[965]$_DFFE_PN0P_  (.D(_02835_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[966]$_DFFE_PN0P_  (.D(_02836_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[967]$_DFFE_PN0P_  (.D(_02837_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[968]$_DFFE_PN0P_  (.D(_02838_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[969]$_DFFE_PN0P_  (.D(_02839_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[96]$_DFFE_PN0P_  (.D(_02840_),
    .RN(net2033),
    .CLK(clknet_leaf_33_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[970]$_DFFE_PN0P_  (.D(_02841_),
    .RN(net2034),
    .CLK(clknet_leaf_27_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[971]$_DFFE_PN0P_  (.D(_02842_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[972]$_DFFE_PN0P_  (.D(_02843_),
    .RN(net153),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[973]$_DFFE_PN0P_  (.D(_02844_),
    .RN(net2036),
    .CLK(clknet_leaf_20_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[974]$_DFFE_PN0P_  (.D(_02845_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[975]$_DFFE_PN0P_  (.D(_02846_),
    .RN(net153),
    .CLK(clknet_leaf_21_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[976]$_DFFE_PN0P_  (.D(_02847_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[977]$_DFFE_PN0P_  (.D(_02848_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[978]$_DFFE_PN0P_  (.D(_02849_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[979]$_DFFE_PN0P_  (.D(_02850_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[97]$_DFFE_PN0P_  (.D(_02851_),
    .RN(net2033),
    .CLK(clknet_leaf_30_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[980]$_DFFE_PN0P_  (.D(_02852_),
    .RN(net2037),
    .CLK(clknet_leaf_8_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[981]$_DFFE_PN0P_  (.D(_02853_),
    .RN(net153),
    .CLK(clknet_leaf_22_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[982]$_DFFE_PN0P_  (.D(_02854_),
    .RN(net153),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[983]$_DFFE_PN0P_  (.D(_02855_),
    .RN(net2036),
    .CLK(clknet_leaf_19_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[984]$_DFFE_PN0P_  (.D(_02856_),
    .RN(net153),
    .CLK(clknet_leaf_24_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[985]$_DFFE_PN0P_  (.D(_02857_),
    .RN(net153),
    .CLK(clknet_leaf_15_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[986]$_DFFE_PN0P_  (.D(_02858_),
    .RN(net2036),
    .CLK(clknet_leaf_9_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[987]$_DFFE_PN0P_  (.D(_02859_),
    .RN(net2036),
    .CLK(clknet_leaf_13_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[988]$_DFFE_PN0P_  (.D(_02860_),
    .RN(net153),
    .CLK(clknet_leaf_7_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[989]$_DFFE_PN0P_  (.D(_02861_),
    .RN(net2036),
    .CLK(clknet_leaf_10_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[98]$_DFFE_PN0P_  (.D(_02862_),
    .RN(net2033),
    .CLK(clknet_leaf_28_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[990]$_DFFE_PN0P_  (.D(_02863_),
    .RN(net2036),
    .CLK(clknet_leaf_12_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[991]$_DFFE_PN0P_  (.D(_02864_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[992]$_DFFE_PN0P_  (.D(_02865_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[993]$_DFFE_PN0P_  (.D(_02866_),
    .RN(net2033),
    .CLK(clknet_leaf_32_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[994]$_DFFE_PN0P_  (.D(_02867_),
    .RN(net2033),
    .CLK(clknet_leaf_31_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[995]$_DFFE_PN0P_  (.D(_02868_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[996]$_DFFE_PN0P_  (.D(_02869_),
    .RN(net2033),
    .CLK(clknet_leaf_29_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[997]$_DFFE_PN0P_  (.D(_02870_),
    .RN(net2034),
    .CLK(clknet_leaf_4_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[998]$_DFFE_PN0P_  (.D(_02871_),
    .RN(net2033),
    .CLK(clknet_leaf_0_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[999]$_DFFE_PN0P_  (.D(_02872_),
    .RN(net153),
    .CLK(clknet_leaf_3_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gen_regfile_ff.register_file_i.rf_reg[99]$_DFFE_PN0P_  (.D(_02873_),
    .RN(net2034),
    .CLK(clknet_leaf_16_clk_i_regs),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.branch_set$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .RN(net2034),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.branch_set ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_02874_),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_02875_),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_02876_),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_02877_),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.debug_mode_o$_DFFE_PN0P_  (.D(_02878_),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.debug_mode_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.exc_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.illegal_insn_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_i ),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.load_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.nmi_mode_o$_DFFE_PN0P_  (.D(_02879_),
    .RN(net2035),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.nmi_mode_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_i ),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.store_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_02880_),
    .RN(net2034),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.id_fsm_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[0]$_DFFE_PN0P_  (.D(_02881_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[10]$_DFFE_PN0P_  (.D(_02882_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[11]$_DFFE_PN0P_  (.D(_02883_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[12]$_DFFE_PN0P_  (.D(_02884_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[13]$_DFFE_PN0P_  (.D(_02885_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[14]$_DFFE_PN0P_  (.D(_02886_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[15]$_DFFE_PN0P_  (.D(_02887_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[16]$_DFFE_PN0P_  (.D(_02888_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[17]$_DFFE_PN0P_  (.D(_02889_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[18]$_DFFE_PN0P_  (.D(_02890_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[19]$_DFFE_PN0P_  (.D(_02891_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[1]$_DFFE_PN0P_  (.D(_02892_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[20]$_DFFE_PN0P_  (.D(_02893_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[21]$_DFFE_PN0P_  (.D(_02894_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[22]$_DFFE_PN0P_  (.D(_02895_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[23]$_DFFE_PN0P_  (.D(_02896_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[24]$_DFFE_PN0P_  (.D(_02897_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[25]$_DFFE_PN0P_  (.D(_02898_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[26]$_DFFE_PN0P_  (.D(_02899_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[27]$_DFFE_PN0P_  (.D(_02900_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[28]$_DFFE_PN0P_  (.D(_02901_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[29]$_DFFE_PN0P_  (.D(_02902_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[2]$_DFFE_PN0P_  (.D(_02903_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[30]$_DFFE_PN0P_  (.D(_02904_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[31]$_DFFE_PN0P_  (.D(_02905_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[34]$_DFFE_PN0P_  (.D(_02906_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[35]$_DFFE_PN0P_  (.D(_02907_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[36]$_DFFE_PN0P_  (.D(_02908_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[37]$_DFFE_PN0P_  (.D(_02909_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[38]$_DFFE_PN0P_  (.D(_02910_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[39]$_DFFE_PN0P_  (.D(_02911_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[3]$_DFFE_PN0P_  (.D(_02912_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[40]$_DFFE_PN0P_  (.D(_02913_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[41]$_DFFE_PN0P_  (.D(_02914_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[42]$_DFFE_PN0P_  (.D(_02915_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[43]$_DFFE_PN0P_  (.D(_02916_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[44]$_DFFE_PN0P_  (.D(_02917_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[45]$_DFFE_PN0P_  (.D(_02918_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[46]$_DFFE_PN0P_  (.D(_02919_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[47]$_DFFE_PN0P_  (.D(_02920_),
    .RN(net2037),
    .CLK(clknet_leaf_30_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[48]$_DFFE_PN0P_  (.D(_02921_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[49]$_DFFE_PN0P_  (.D(_02922_),
    .RN(net2037),
    .CLK(clknet_leaf_25_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[4]$_DFFE_PN0P_  (.D(_02923_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[50]$_DFFE_PN0P_  (.D(_02924_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[51]$_DFFE_PN0P_  (.D(_02925_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[52]$_DFFE_PN0P_  (.D(_02926_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[53]$_DFFE_PN0P_  (.D(_02927_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[54]$_DFFE_PN0P_  (.D(_02928_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[55]$_DFFE_PN0P_  (.D(_02929_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[56]$_DFFE_PN0P_  (.D(_02930_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[57]$_DFFE_PN0P_  (.D(_02931_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[58]$_DFFE_PN0P_  (.D(_02932_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[59]$_DFFE_PN0P_  (.D(_02933_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[5]$_DFFE_PN0P_  (.D(_02934_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[60]$_DFFE_PN0P_  (.D(_02935_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[61]$_DFFE_PN0P_  (.D(_02936_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[62]$_DFFE_PN0P_  (.D(_02937_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[63]$_DFFE_PN0P_  (.D(_02938_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[64]$_DFFE_PN0P_  (.D(_02939_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[65]$_DFFE_PN0P_  (.D(_02940_),
    .RN(net2037),
    .CLK(clknet_leaf_26_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[66]$_DFFE_PN0P_  (.D(_02941_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[67]$_DFFE_PN0P_  (.D(_02942_),
    .RN(net2037),
    .CLK(clknet_leaf_28_clk),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[6]$_DFFE_PN0P_  (.D(_02943_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[7]$_DFFE_PN0P_  (.D(_02944_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[8]$_DFFE_PN0P_  (.D(_02945_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \id_stage_i.imd_val_q_ex_o[9]$_DFFE_PN0P_  (.D(_02946_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\ex_block_i.alu_i.imd_val_q_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(_02947_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(_02948_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(_02949_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(_02950_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(_02951_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(_02952_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(_02953_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(_02954_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(_02955_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(_02956_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(_02957_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(_02958_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(_02959_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(_02960_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(_02961_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(_02962_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(_02963_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(_02964_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(_02965_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(_02966_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(_02967_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(_02968_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(_02969_),
    .CLK(clknet_leaf_3_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(_02970_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(_02971_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(_02972_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(_02973_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(_02974_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(_02975_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(_02976_),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(_02977_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(_02978_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(_02979_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(_02980_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(_02981_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_if_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(_02982_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_if_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(_02983_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(_02984_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(_02985_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_if_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(_02986_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(_02987_),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.pc_if_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(_02988_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(_02989_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(_02990_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(_02991_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(_02992_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(_02993_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(_02994_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(_02995_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(_02996_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(_02997_),
    .CLK(clknet_leaf_3_clk),
    .Q(\cs_registers_i.pc_if_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(_02998_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_if_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(_02999_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_if_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(_03000_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_if_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(_03001_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_if_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(_03002_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(_03003_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_if_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(_03004_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(_03005_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(_03006_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(_03007_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_if_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(_03008_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(_03009_),
    .CLK(clknet_leaf_2_clk),
    .Q(\cs_registers_i.pc_if_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(_03010_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_if_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(_03011_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(_03012_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(_03013_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(_03014_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(_03015_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(_03016_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(_03017_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(_03018_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(_03019_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(_03020_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(_03021_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(_03022_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(_03023_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(_03024_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(_03025_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(_03026_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(_03027_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(_03028_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(_03029_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(_03030_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(_03031_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(_03032_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(_03033_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(_03034_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(_03035_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(_03036_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(_03037_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(_03038_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(_03039_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(_03040_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(_03041_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(_03042_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(_03043_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(_03044_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(_03045_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(_03046_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(_03047_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(_03048_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(_03049_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(_03050_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(_03051_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(_03052_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(_03053_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(_03054_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(_03055_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(_03056_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(_03057_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(_03058_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(_03059_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(_03060_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(_03061_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(_03062_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(_03063_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(_03064_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(_03065_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(_03066_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(_03067_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(_03068_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(_03069_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(_03070_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(_03071_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(_03072_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(_03073_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(_03074_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(_03075_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(_03076_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(_03077_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(_03078_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(_03079_),
    .CLK(clknet_leaf_35_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(_03080_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(_03081_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(_03082_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(_03083_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(_03084_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(_03085_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(_03086_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(_03087_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(_03088_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(_03089_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(_03090_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(_03091_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(_03092_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(_03093_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(_03094_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(_03095_),
    .CLK(clknet_leaf_36_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(_03096_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(_03097_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(_03098_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(_03099_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(_03100_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(_03101_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(_03102_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(_03103_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(_03104_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(_03105_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(_03106_),
    .CLK(clknet_leaf_37_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .RN(net2034),
    .CLK(clknet_leaf_2_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(_03107_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(_03108_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(_03109_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(_03110_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(_03111_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(_03112_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(_03113_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(_03114_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(_03115_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(_03116_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(_03117_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(_03118_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(_03119_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(_03120_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(_03121_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(_03122_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(_03123_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(_03124_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(_03125_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(_03126_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(_03127_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(_03128_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(_03129_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(_03130_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(_03131_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(_03132_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(_03133_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(_03134_),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(_03135_),
    .CLK(clknet_leaf_0_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(_03136_),
    .CLK(clknet_leaf_38_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .RN(net2034),
    .CLK(clknet_leaf_1_clk),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(_03137_),
    .CLK(clknet_leaf_34_clk),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(_03138_),
    .CLK(clknet_leaf_2_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_03139_),
    .CLK(clknet_leaf_2_clk),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(_03140_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(_03141_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(_03142_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_03143_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_03144_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_03145_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_03146_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_03147_),
    .CLK(clknet_leaf_34_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_03148_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(_03149_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(_03150_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(_03151_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(_03152_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(_03153_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(_03154_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_03155_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(_03156_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[0]$_DFFE_PN_  (.D(_03157_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[10]$_DFFE_PN_  (.D(_03158_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[11]$_DFFE_PN_  (.D(_03159_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[12]$_DFFE_PN_  (.D(_03160_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[13]$_DFFE_PN_  (.D(_03161_),
    .CLK(clknet_leaf_34_clk),
    .Q(\id_stage_i.controller_i.instr_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[14]$_DFFE_PN_  (.D(_03162_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[15]$_DFFE_PN_  (.D(_03163_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[16]$_DFFE_PN_  (.D(_03164_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[17]$_DFFE_PN_  (.D(_03165_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[18]$_DFFE_PN_  (.D(_03166_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[19]$_DFFE_PN_  (.D(_03167_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[1]$_DFFE_PN_  (.D(_03168_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[20]$_DFFE_PN_  (.D(_03169_),
    .CLK(clknet_leaf_35_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[21]$_DFFE_PN_  (.D(_03170_),
    .CLK(clknet_leaf_35_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[22]$_DFFE_PN_  (.D(_03171_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[23]$_DFFE_PN_  (.D(_03172_),
    .CLK(clknet_leaf_35_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[24]$_DFFE_PN_  (.D(_03173_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[25]$_DFFE_PN_  (.D(_03174_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[26]$_DFFE_PN_  (.D(_03175_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[27]$_DFFE_PN_  (.D(_03176_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[28]$_DFFE_PN_  (.D(_03177_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[29]$_DFFE_PN_  (.D(_03178_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[2]$_DFFE_PN_  (.D(_03179_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[30]$_DFFE_PN_  (.D(_03180_),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.instr_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[31]$_DFFE_PN_  (.D(_03181_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[3]$_DFFE_PN_  (.D(_03182_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[4]$_DFFE_PN_  (.D(_03183_),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_4 \if_stage_i.instr_rdata_id_o[5]$_DFFE_PN_  (.D(_03184_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[6]$_DFFE_PN_  (.D(_03185_),
    .CLK(clknet_leaf_33_clk),
    .Q(\id_stage_i.controller_i.instr_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[7]$_DFFE_PN_  (.D(_03186_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[8]$_DFFE_PN_  (.D(_03187_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.instr_rdata_id_o[9]$_DFFE_PN_  (.D(_03188_),
    .CLK(clknet_leaf_34_clk),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \if_stage_i.instr_valid_id_o$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .RN(net2034),
    .CLK(clknet_leaf_7_clk),
    .Q(\id_stage_i.controller_i.instr_valid_i ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(_03189_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(_03190_),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.pc_id_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(_03191_),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.pc_id_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(_03192_),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.pc_id_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(_03193_),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.pc_id_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(_03194_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_id_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(_03195_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(_03196_),
    .CLK(clknet_leaf_5_clk),
    .Q(\cs_registers_i.pc_id_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(_03197_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(_03198_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(_03199_),
    .CLK(clknet_leaf_7_clk),
    .Q(\cs_registers_i.pc_id_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(_03200_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(_03201_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(_03202_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(_03203_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(_03204_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(_03205_),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.pc_id_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(_03206_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(_03207_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(_03208_),
    .CLK(clknet_leaf_4_clk),
    .Q(\cs_registers_i.pc_id_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(_03209_),
    .CLK(clknet_leaf_14_clk),
    .Q(\cs_registers_i.pc_id_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(_03210_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(_03211_),
    .CLK(clknet_leaf_13_clk),
    .Q(\cs_registers_i.pc_id_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(_03212_),
    .CLK(clknet_leaf_12_clk),
    .Q(\cs_registers_i.pc_id_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(_03213_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(_03214_),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.pc_id_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(_03215_),
    .CLK(clknet_leaf_8_clk),
    .Q(\cs_registers_i.pc_id_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(_03216_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(_03217_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(_03218_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(_03219_),
    .CLK(clknet_leaf_6_clk),
    .Q(\cs_registers_i.pc_id_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[0]$_DFFE_PN0P_  (.D(_03220_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[10]$_DFFE_PN0P_  (.D(_03221_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[11]$_DFFE_PN0P_  (.D(_03222_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[12]$_DFFE_PN0P_  (.D(_03223_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[13]$_DFFE_PN0P_  (.D(_03224_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[14]$_DFFE_PN0P_  (.D(_03225_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[15]$_DFFE_PN0P_  (.D(_03226_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[16]$_DFFE_PN0P_  (.D(_03227_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[17]$_DFFE_PN0P_  (.D(_03228_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[18]$_DFFE_PN0P_  (.D(_03229_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[19]$_DFFE_PN0P_  (.D(_03230_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[1]$_DFFE_PN0P_  (.D(_03231_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[20]$_DFFE_PN0P_  (.D(_03232_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[21]$_DFFE_PN0P_  (.D(_03233_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[22]$_DFFE_PN0P_  (.D(_03234_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[23]$_DFFE_PN0P_  (.D(_03235_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[24]$_DFFE_PN0P_  (.D(_03236_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[25]$_DFFE_PN0P_  (.D(_03237_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[26]$_DFFE_PN0P_  (.D(_03238_),
    .RN(net2034),
    .CLK(clknet_leaf_24_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[27]$_DFFE_PN0P_  (.D(_03239_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[28]$_DFFE_PN0P_  (.D(_03240_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[29]$_DFFE_PN0P_  (.D(_03241_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[2]$_DFFE_PN0P_  (.D(_03242_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[30]$_DFFE_PN0P_  (.D(_03243_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[31]$_DFFE_PN0P_  (.D(_03244_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[3]$_DFFE_PN0P_  (.D(_03245_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[4]$_DFFE_PN0P_  (.D(_03246_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[5]$_DFFE_PN0P_  (.D(_03247_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[6]$_DFFE_PN0P_  (.D(_03248_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[7]$_DFFE_PN0P_  (.D(_03249_),
    .RN(net2034),
    .CLK(clknet_leaf_8_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[8]$_DFFE_PN0P_  (.D(_03250_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.addr_last_o[9]$_DFFE_PN0P_  (.D(_03251_),
    .RN(net2034),
    .CLK(clknet_leaf_9_clk),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_03252_),
    .RN(net2037),
    .CLK(clknet_leaf_31_clk),
    .Q(\load_store_unit_i.data_sign_ext_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_03253_),
    .RN(net2034),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.data_we_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_03254_),
    .RN(net153),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.handle_misaligned_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_03255_),
    .RN(net153),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_03256_),
    .RN(net153),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_03257_),
    .RN(net2034),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_03258_),
    .RN(net2034),
    .CLK(clknet_leaf_33_clk),
    .Q(\load_store_unit_i.lsu_err_q ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_03259_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_offset_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_03260_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_offset_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_03261_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_03262_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_03263_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_03264_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_03265_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_03266_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_03267_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_03268_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_03269_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_03270_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_03271_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_03272_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_03273_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_03274_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_03275_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_03276_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_03277_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_03278_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_03279_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_03280_),
    .RN(net2036),
    .CLK(clknet_leaf_29_clk),
    .Q(\load_store_unit_i.rdata_q[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_03281_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_03282_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_03283_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_03284_),
    .RN(net2036),
    .CLK(clknet_leaf_32_clk),
    .Q(\load_store_unit_i.rdata_q[9] ));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22866__1 (.ZN(alert_major_o));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22867__2 (.ZN(alert_minor_o));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22868__3 (.ZN(data_addr_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22869__4 (.ZN(data_addr_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22900__5 (.ZN(instr_addr_o[0]));
 gf180mcu_fd_sc_mcu9t5v0__tiel _22901__6 (.ZN(instr_addr_o[1]));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1741 (.I(net1739),
    .Z(net1740));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1740 (.I(_07763_),
    .Z(net1739));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1747 (.I(_09965_),
    .Z(net1746));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1742 (.I(net2177),
    .Z(net1741));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1743 (.I(_07603_),
    .Z(net1742));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1744 (.I(_06969_),
    .Z(net1743));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1745 (.I(_06964_),
    .Z(net1744));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1746 (.I(_06936_),
    .Z(net1745));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1748 (.I(_09962_),
    .Z(net1747));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1749 (.I(_09840_),
    .Z(net1748));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1787 (.I(net1785),
    .Z(net1786));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1751 (.I(_09668_),
    .Z(net1750));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1752 (.I(_09660_),
    .Z(net1751));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1781 (.I(net1779),
    .Z(net1780));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1766 (.I(_08954_),
    .Z(net1765));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1753 (.I(_09421_),
    .Z(net1752));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1754 (.I(_09405_),
    .Z(net1753));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1755 (.I(_09374_),
    .Z(net1754));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1756 (.I(_09358_),
    .Z(net1755));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1757 (.I(_09322_),
    .Z(net1756));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1758 (.I(_09258_),
    .Z(net1757));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1759 (.I(_09223_),
    .Z(net1758));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1760 (.I(_09166_),
    .Z(net1759));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1761 (.I(_09131_),
    .Z(net1760));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1762 (.I(_09079_),
    .Z(net1761));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1763 (.I(_09042_),
    .Z(net1762));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1764 (.I(_08981_),
    .Z(net1763));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1765 (.I(_08961_),
    .Z(net1764));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1767 (.I(_08941_),
    .Z(net1766));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1768 (.I(_08889_),
    .Z(net1767));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1769 (.I(_08852_),
    .Z(net1768));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1770 (.I(_08793_),
    .Z(net1769));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1771 (.I(_08775_),
    .Z(net1770));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1772 (.I(_08755_),
    .Z(net1771));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1773 (.I(_08690_),
    .Z(net1772));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1774 (.I(_08649_),
    .Z(net1773));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1775 (.I(_08586_),
    .Z(net1774));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1776 (.I(_08427_),
    .Z(net1775));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1777 (.I(_08378_),
    .Z(net1776));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1778 (.I(_08361_),
    .Z(net1777));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1779 (.I(_08339_),
    .Z(net1778));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1780 (.I(_08291_),
    .Z(net1779));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1782 (.I(_08252_),
    .Z(net1781));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1783 (.I(_08214_),
    .Z(net1782));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1784 (.I(_08187_),
    .Z(net1783));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1785 (.I(_08098_),
    .Z(net1784));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1786 (.I(_08074_),
    .Z(net1785));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1788 (.I(_07993_),
    .Z(net1787));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1795 (.I(net1793),
    .Z(net1794));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1793 (.I(net1791),
    .Z(net1792));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1791 (.I(net1789),
    .Z(net1790));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1789 (.I(_07904_),
    .Z(net1788));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1790 (.I(_07880_),
    .Z(net1789));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1792 (.I(_07857_),
    .Z(net1791));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1794 (.I(_07829_),
    .Z(net1793));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1796 (.I(_07805_),
    .Z(net1795));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2008 (.I(net2005),
    .Z(net2007));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1814 (.I(_08597_),
    .Z(net1813));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1797 (.I(_07740_),
    .Z(net1796));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1798 (.I(_07693_),
    .Z(net1797));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1813 (.I(_08704_),
    .Z(net1812));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1799 (.I(_07691_),
    .Z(net1798));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1800 (.I(_07647_),
    .Z(net1799));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1809 (.I(_09937_),
    .Z(net1808));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 place1801 (.I(_07636_),
    .Z(net1800));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1804 (.I(net1802),
    .Z(net1803));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1802 (.I(_07610_),
    .Z(net1801));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1803 (.I(_07549_),
    .Z(net1802));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1805 (.I(_07030_),
    .Z(net1804));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1807 (.I(_05835_),
    .Z(net1806));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1808 (.I(_04342_),
    .Z(net1807));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1810 (.I(_09619_),
    .Z(net1809));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1811 (.I(_08949_),
    .Z(net1810));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1812 (.I(_08711_),
    .Z(net1811));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2007 (.I(net2005),
    .Z(net2006));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1816 (.I(net1814),
    .Z(net1815));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1815 (.I(_08182_),
    .Z(net1814));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place2006 (.I(net2093),
    .Z(net2005));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2005 (.I(net2137),
    .Z(net2004));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2004 (.I(net2002),
    .Z(net2003));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1822 (.I(_08657_),
    .Z(net1821));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1819 (.I(net2483),
    .Z(net1818));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1818 (.I(_07555_),
    .Z(net1817));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1817 (.I(_07620_),
    .Z(net1816));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1820 (.I(_06473_),
    .Z(net1819));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1821 (.I(_08657_),
    .Z(net1820));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2003 (.I(net2055),
    .Z(net2002));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2002 (.I(net1999),
    .Z(net2001));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place2001 (.I(net1999),
    .Z(net2000));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1823 (.I(_08596_),
    .Z(net1822));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1824 (.I(_08199_),
    .Z(net1823));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1825 (.I(_08197_),
    .Z(net1824));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1826 (.I(_08181_),
    .Z(net1825));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1827 (.I(_07999_),
    .Z(net1826));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2000 (.I(net2093),
    .Z(net1999));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1828 (.I(_07842_),
    .Z(net1827));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1999 (.I(net1989),
    .Z(net1998));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1830 (.I(_07745_),
    .Z(net1829));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1829 (.I(_07745_),
    .Z(net1828));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1838 (.I(_09753_),
    .Z(net1837));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1831 (.I(_07684_),
    .Z(net1830));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1837 (.I(_09753_),
    .Z(net1836));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1832 (.I(_07596_),
    .Z(net1831));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1833 (.I(_07547_),
    .Z(net1832));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1834 (.I(_04560_),
    .Z(net1833));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1835 (.I(_10016_),
    .Z(net1834));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1836 (.I(_09930_),
    .Z(net1835));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place1998 (.I(net1996),
    .Z(net1997));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1839 (.I(_09749_),
    .Z(net1838));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1989 (.I(net1983),
    .Z(net1988));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1840 (.I(_09745_),
    .Z(net1839));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1988 (.I(net1983),
    .Z(net1987));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1841 (.I(_09650_),
    .Z(net1840));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1987 (.I(net1983),
    .Z(net1986));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1842 (.I(_08192_),
    .Z(net1841));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1845 (.I(_08010_),
    .Z(net1844));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1844 (.I(net1842),
    .Z(net1843));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1843 (.I(_08010_),
    .Z(net1842));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1986 (.I(net1983),
    .Z(net1985));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1984 (.I(net1972),
    .Z(net1983));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1983 (.I(net1976),
    .Z(net1982));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1852 (.I(net1847),
    .Z(net1851));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1982 (.I(net1980),
    .Z(net1981));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1853 (.I(net1847),
    .Z(net1852));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1985 (.I(net1983),
    .Z(net1984));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1846 (.I(_07947_),
    .Z(net1845));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1851 (.I(net1847),
    .Z(net1850));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1850 (.I(net1847),
    .Z(net1849));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1847 (.I(_07689_),
    .Z(net1846));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1849 (.I(net1847),
    .Z(net1848));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1848 (.I(_07681_),
    .Z(net1847));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1958 (.I(net2058),
    .Z(net1957));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1855 (.I(_07666_),
    .Z(net1854));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1854 (.I(_07666_),
    .Z(net1853));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1957 (.I(net2128),
    .Z(net1956));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1956 (.I(net2128),
    .Z(net1955));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1931 (.I(net1927),
    .Z(net1930));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1930 (.I(net1927),
    .Z(net1929));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1929 (.I(net1927),
    .Z(net1928));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1928 (.I(net1913),
    .Z(net1927));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1858 (.I(_07666_),
    .Z(net1857));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1857 (.I(_07666_),
    .Z(net1856));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1856 (.I(net1854),
    .Z(net1855));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1926 (.I(net1922),
    .Z(net1925));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1860 (.I(_07665_),
    .Z(net1859));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1859 (.I(_07665_),
    .Z(net1858));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1925 (.I(net1922),
    .Z(net1924));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1884 (.I(net1882),
    .Z(net1883));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1885 (.I(_07518_),
    .Z(net1884));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1861 (.I(_07657_),
    .Z(net1860));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1863 (.I(net1861),
    .Z(net1862));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1862 (.I(_07657_),
    .Z(net1861));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1883 (.I(_07518_),
    .Z(net1882));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1882 (.I(_07518_),
    .Z(net1881));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1880 (.I(net1877),
    .Z(net1879));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1876 (.I(net1874),
    .Z(net1875));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1875 (.I(net1871),
    .Z(net1874));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1881 (.I(net1877),
    .Z(net1880));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1874 (.I(net1872),
    .Z(net1873));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1873 (.I(net1871),
    .Z(net1872));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1868 (.I(_07537_),
    .Z(net1867));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1867 (.I(_07537_),
    .Z(net1866));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1866 (.I(net1864),
    .Z(net1865));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1865 (.I(_07537_),
    .Z(net1864));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1872 (.I(_07534_),
    .Z(net1871));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1869 (.I(_07534_),
    .Z(net1868));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1871 (.I(net1869),
    .Z(net1870));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1870 (.I(_07534_),
    .Z(net1869));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1877 (.I(_07523_),
    .Z(net1876));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1878 (.I(_07518_),
    .Z(net1877));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1924 (.I(net1922),
    .Z(net1923));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1918 (.I(net1916),
    .Z(net1917));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1917 (.I(net1913),
    .Z(net1916));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1916 (.I(net2179),
    .Z(net1915));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1915 (.I(net1913),
    .Z(net1914));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1914 (.I(net2090),
    .Z(net1913));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1887 (.I(\load_store_unit_i.rdata_offset_q[1] ),
    .Z(net1886));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1886 (.I(_01354_),
    .Z(net1885));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1923 (.I(net1913),
    .Z(net1922));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1922 (.I(net1918),
    .Z(net1921));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1921 (.I(net1918),
    .Z(net1920));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1920 (.I(net1918),
    .Z(net1919));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1919 (.I(net1913),
    .Z(net1918));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1888 (.I(\load_store_unit_i.rdata_offset_q[0] ),
    .Z(net1887));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1903 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net1902));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1889 (.I(\id_stage_i.controller_i.instr_i[6] ),
    .Z(net1888));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1902 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net1901));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 place1890 (.I(\id_stage_i.controller_i.instr_i[4] ),
    .Z(net1889));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1891 (.I(\id_stage_i.controller_i.instr_i[3] ),
    .Z(net1890));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1892 (.I(\id_stage_i.controller_i.instr_i[31] ),
    .Z(net1891));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1893 (.I(\id_stage_i.controller_i.instr_i[30] ),
    .Z(net1892));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 place1894 (.I(\id_stage_i.controller_i.instr_i[2] ),
    .Z(net1893));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1895 (.I(\id_stage_i.controller_i.instr_i[29] ),
    .Z(net1894));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1896 (.I(\id_stage_i.controller_i.instr_i[28] ),
    .Z(net1895));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1897 (.I(\id_stage_i.controller_i.instr_i[27] ),
    .Z(net1896));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1898 (.I(\id_stage_i.controller_i.instr_i[26] ),
    .Z(net1897));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1899 (.I(\id_stage_i.controller_i.instr_i[25] ),
    .Z(net1898));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1900 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .Z(net1899));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1901 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .Z(net1900));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1906 (.I(net2101),
    .Z(net1905));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1905 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net1904));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1904 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .Z(net1903));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1913 (.I(net1909),
    .Z(net1912));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1907 (.I(net2090),
    .Z(net1906));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1912 (.I(net1909),
    .Z(net1911));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1911 (.I(net2089),
    .Z(net1910));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1908 (.I(net2090),
    .Z(net1907));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1910 (.I(net2090),
    .Z(net1909));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1909 (.I(net1907),
    .Z(net1908));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place1932 (.I(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .Z(net1931));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1954 (.I(net1944),
    .Z(net1953));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1948 (.I(net2128),
    .Z(net1947));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1947 (.I(net1944),
    .Z(net1946));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1937 (.I(net1933),
    .Z(net1936));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1933 (.I(net2104),
    .Z(net1932));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1936 (.I(net1933),
    .Z(net1935));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1935 (.I(net1933),
    .Z(net1934));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1934 (.I(net2154),
    .Z(net1933));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1946 (.I(net2114),
    .Z(net1945));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1945 (.I(net2058),
    .Z(net1944));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 place1944 (.I(net2139),
    .Z(net1943));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place1943 (.I(net2141),
    .Z(net1942));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1942 (.I(net2141),
    .Z(net1941));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1941 (.I(net2141),
    .Z(net1940));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1938 (.I(net2140),
    .Z(net1937));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1940 (.I(net2140),
    .Z(net1939));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1939 (.I(net2139),
    .Z(net1938));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1953 (.I(net1944),
    .Z(net1952));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1952 (.I(net2128),
    .Z(net1951));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1951 (.I(net1944),
    .Z(net1950));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1950 (.I(net1944),
    .Z(net1949));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1949 (.I(net2128),
    .Z(net1948));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1962 (.I(net1959),
    .Z(net1961));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1972 (.I(net1968),
    .Z(net1971));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1971 (.I(net1968),
    .Z(net1970));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1970 (.I(net1968),
    .Z(net1969));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1969 (.I(net1966),
    .Z(net1968));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1980 (.I(net1976),
    .Z(net1979));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1979 (.I(net1976),
    .Z(net1978));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1978 (.I(net1976),
    .Z(net1977));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1977 (.I(net1972),
    .Z(net1976));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1976 (.I(net1972),
    .Z(net1975));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1968 (.I(net1966),
    .Z(net1967));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1964 (.I(net1962),
    .Z(net1963));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1963 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .Z(net1962));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1967 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net1966));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1966 (.I(net1964),
    .Z(net1965));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1965 (.I(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .Z(net1964));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1997 (.I(net1989),
    .Z(net1996));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1992 (.I(net1990),
    .Z(net1991));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place1991 (.I(net1989),
    .Z(net1990));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 place1990 (.I(net2093),
    .Z(net1989));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1996 (.I(net1989),
    .Z(net1995));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1995 (.I(net1989),
    .Z(net1994));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1994 (.I(net1990),
    .Z(net1993));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1993 (.I(net1990),
    .Z(net1992));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2045 (.I(net144),
    .Z(net2044));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2038 (.I(net2036),
    .Z(net2037));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place2037 (.I(net153),
    .Z(net2036));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2036 (.I(net2034),
    .Z(net2035));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 place2023 (.I(net2021),
    .Z(net2022));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place2020 (.I(\id_stage_i.controller_i.instr_i[14] ),
    .Z(net2019));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_22_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_22_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_clk_i_regs (.I(clknet_2_0__leaf_clk_i_regs),
    .Z(clknet_leaf_0_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_1_0__f_clk_i (.I(clknet_0_clk_i),
    .Z(clknet_1_0__leaf_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2047 (.I(net142),
    .Z(net2046));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_0_clk_i (.I(clk_i),
    .Z(clknet_0_clk_i));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_regs_0_core_clock (.I(delaynet_4_core_clock),
    .Z(clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2051 (.I(net134),
    .Z(net2050));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2050 (.I(net137),
    .Z(net2049));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2049 (.I(net138),
    .Z(net2048));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2048 (.I(net141),
    .Z(net2047));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_21_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_21_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_20_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_20_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_15_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_14_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_13_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_12_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_1_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_11_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_10_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_2_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_9_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_4_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_3_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_8_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_clk_i_regs (.I(clknet_2_1__leaf_clk_i_regs),
    .Z(clknet_leaf_7_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_6_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_clk_i_regs (.I(clknet_2_3__leaf_clk_i_regs),
    .Z(clknet_leaf_5_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_19_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_18_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_16_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_clk_i_regs (.I(clknet_2_2__leaf_clk_i_regs),
    .Z(clknet_leaf_17_clk_i_regs));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2025 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Z(net2024));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2026 (.I(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Z(net2025));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2029 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Z(net2028));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2030 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Z(net2029));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2031 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Z(net2030));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2032 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Z(net2031));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2033 (.I(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Z(net2032));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 place2034 (.I(net153),
    .Z(net2033));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2044 (.I(net145),
    .Z(net2043));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2042 (.I(net147),
    .Z(net2041));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2041 (.I(net148),
    .Z(net2040));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2040 (.I(net149),
    .Z(net2039));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place2039 (.I(net150),
    .Z(net2038));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1363 (.I(_05009_),
    .Z(net1362));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 place1369 (.I(_05065_),
    .Z(net1368));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 place1374 (.I(_04981_),
    .Z(net1373));
endmodule
