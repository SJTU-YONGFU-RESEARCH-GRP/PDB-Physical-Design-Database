module parameterized_pwm (clk,
    enable,
    pwm_out,
    rst_n,
    div,
    duty);
 input clk;
 input enable;
 output pwm_out;
 input rst_n;
 input [15:0] div;
 input [7:0] duty;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \div_counter[0] ;
 wire \div_counter[10] ;
 wire \div_counter[11] ;
 wire \div_counter[12] ;
 wire \div_counter[13] ;
 wire \div_counter[14] ;
 wire \div_counter[15] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_counter[5] ;
 wire \div_counter[6] ;
 wire \div_counter[7] ;
 wire \div_counter[8] ;
 wire \div_counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _235_ (.I(net8),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _236_ (.I(net10),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _237_ (.I(net9),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _238_ (.I(net14),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _239_ (.I(net13),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _240_ (.I(net11),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _241_ (.I(net12),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _242_ (.I(net7),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _243_ (.I(net6),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _244_ (.I(net5),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _245_ (.I(net4),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _246_ (.I(net3),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _247_ (.I(net2),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _248_ (.I(net16),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _249_ (.I(net15),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _250_ (.I(\counter[7] ),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _251_ (.I(\counter[6] ),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _252_ (.I(\counter[5] ),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _253_ (.I(\counter[4] ),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _254_ (.I(\counter[3] ),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _255_ (.I(\counter[2] ),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _256_ (.I(\counter[1] ),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _257_ (.I(\div_counter[0] ),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _258_ (.I(net17),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _259_ (.I(net26),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _260_ (.A1(_025_),
    .A2(\counter[0] ),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _261_ (.I(net26),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _262_ (.A1(\counter[4] ),
    .A2(\counter[2] ),
    .A3(\counter[3] ),
    .A4(_207_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _263_ (.A1(\counter[7] ),
    .A2(\counter[6] ),
    .A3(\counter[5] ),
    .A4(_028_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _264_ (.A1(_027_),
    .A2(\counter[0] ),
    .A3(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _265_ (.A1(_167_),
    .A2(_170_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _266_ (.A1(_166_),
    .A2(_031_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _267_ (.I(_160_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _268_ (.A1(_164_),
    .A2(_033_),
    .B(_163_),
    .C(_166_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _269_ (.A1(_164_),
    .A2(_161_),
    .A3(_170_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _270_ (.A1(_169_),
    .A2(_035_),
    .B(_167_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _271_ (.A1(_032_),
    .A2(_034_),
    .B(_036_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _272_ (.A1(_185_),
    .A2(_194_),
    .A3(_191_),
    .A4(_188_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _273_ (.A1(_197_),
    .A2(_206_),
    .A3(_203_),
    .A4(_200_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _274_ (.A1(_038_),
    .A2(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _275_ (.A1(_173_),
    .A2(_176_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _276_ (.A1(_182_),
    .A2(_179_),
    .A3(_040_),
    .A4(_041_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _277_ (.A1(_173_),
    .A2(_176_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _278_ (.A1(_182_),
    .A2(_178_),
    .B(_181_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _279_ (.A1(_173_),
    .A2(_175_),
    .B(_172_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _280_ (.A1(_043_),
    .A2(_044_),
    .B(_045_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _281_ (.A1(_037_),
    .A2(_042_),
    .B1(_046_),
    .B2(_040_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _282_ (.A1(_197_),
    .A2(_200_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _283_ (.A1(_203_),
    .A2(_205_),
    .B(_202_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _284_ (.A1(_197_),
    .A2(_199_),
    .B(_196_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _285_ (.A1(_048_),
    .A2(_049_),
    .B(_050_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _286_ (.A1(net16),
    .A2(net15),
    .A3(net3),
    .A4(net6),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _287_ (.A1(net2),
    .A2(net5),
    .A3(net4),
    .A4(net7),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _288_ (.A1(net8),
    .A2(net1),
    .A3(net10),
    .A4(net13),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _289_ (.A1(net9),
    .A2(net12),
    .A3(net11),
    .A4(net14),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _290_ (.A1(_052_),
    .A2(_053_),
    .A3(_054_),
    .A4(_055_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _291_ (.A1(_191_),
    .A2(_193_),
    .B(_190_),
    .C(_187_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _292_ (.A1(_188_),
    .A2(_187_),
    .B(_185_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _293_ (.A1(_057_),
    .A2(_058_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _294_ (.A1(_184_),
    .A2(_056_),
    .A3(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _295_ (.A1(_038_),
    .A2(_051_),
    .B(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _296_ (.I(net25),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _297_ (.I(_062_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _298_ (.A1(_047_),
    .A2(_061_),
    .B(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _299_ (.I0(_026_),
    .I1(_030_),
    .S(_064_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _300_ (.A1(net26),
    .A2(\counter[1] ),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _301_ (.A1(net26),
    .A2(_208_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _302_ (.I0(_065_),
    .I1(_066_),
    .S(_064_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _303_ (.A1(net26),
    .A2(_226_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _304_ (.A1(net26),
    .A2(\counter[2] ),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _305_ (.I(_164_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _306_ (.I(_163_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _307_ (.A1(_069_),
    .A2(_160_),
    .B(_070_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _308_ (.A1(_169_),
    .A2(_035_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _309_ (.A1(_031_),
    .A2(_071_),
    .B1(_072_),
    .B2(_167_),
    .C(_166_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _310_ (.A1(_182_),
    .A2(_179_),
    .A3(_040_),
    .A4(_041_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _311_ (.A1(_040_),
    .A2(_046_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _312_ (.A1(_038_),
    .A2(_051_),
    .B(_059_),
    .C(_184_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _313_ (.A1(_073_),
    .A2(_074_),
    .B(_075_),
    .C(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _314_ (.A1(_056_),
    .A2(_077_),
    .B(_062_),
    .C(_207_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _315_ (.I0(_067_),
    .I1(_068_),
    .S(_078_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _316_ (.A1(\counter[2] ),
    .A2(\counter[0] ),
    .A3(\counter[1] ),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _317_ (.A1(_029_),
    .A2(_079_),
    .B(_062_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _318_ (.A1(_047_),
    .A2(_061_),
    .B(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _319_ (.A1(_025_),
    .A2(_223_),
    .A3(_079_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _320_ (.A1(_056_),
    .A2(_077_),
    .B(_062_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _321_ (.A1(_027_),
    .A2(_223_),
    .A3(_081_),
    .B1(_082_),
    .B2(_083_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _322_ (.A1(net26),
    .A2(_220_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _323_ (.A1(net26),
    .A2(\counter[4] ),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _324_ (.A1(_062_),
    .A2(\counter[2] ),
    .A3(\counter[3] ),
    .A4(_207_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _325_ (.A1(_056_),
    .A2(_077_),
    .B(_086_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _326_ (.I0(_084_),
    .I1(_085_),
    .S(_087_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _327_ (.A1(\counter[4] ),
    .A2(\counter[3] ),
    .A3(_079_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _328_ (.A1(_029_),
    .A2(_088_),
    .B(_062_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _329_ (.A1(_047_),
    .A2(_061_),
    .B(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _330_ (.A1(_025_),
    .A2(_217_),
    .A3(_088_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _331_ (.A1(_027_),
    .A2(_217_),
    .A3(_090_),
    .B1(_091_),
    .B2(_083_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _332_ (.A1(net26),
    .A2(_214_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _333_ (.A1(net26),
    .A2(\counter[6] ),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _334_ (.A1(_062_),
    .A2(\counter[5] ),
    .A3(_028_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _335_ (.A1(_056_),
    .A2(_077_),
    .B(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _336_ (.I0(_092_),
    .I1(_093_),
    .S(_095_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _337_ (.A1(\counter[6] ),
    .A2(\counter[5] ),
    .A3(_088_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _338_ (.A1(_029_),
    .A2(_096_),
    .B(_062_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _339_ (.A1(_047_),
    .A2(_061_),
    .B(_097_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _340_ (.A1(_025_),
    .A2(_211_),
    .A3(_096_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _341_ (.A1(_027_),
    .A2(_211_),
    .A3(_098_),
    .B1(_099_),
    .B2(_083_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _342_ (.A1(_063_),
    .A2(\div_counter[0] ),
    .A3(_077_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _343_ (.A1(_063_),
    .A2(\div_counter[0] ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _344_ (.A1(_100_),
    .A2(_101_),
    .B(_027_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _345_ (.I(_025_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _346_ (.A1(_062_),
    .A2(_077_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _347_ (.I(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _348_ (.A1(net25),
    .A2(_209_),
    .A3(\div_counter[2] ),
    .A4(\div_counter[3] ),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _349_ (.A1(\div_counter[4] ),
    .A2(_105_),
    .Z(_106_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _350_ (.A1(\div_counter[5] ),
    .A2(\div_counter[6] ),
    .A3(\div_counter[7] ),
    .A4(_106_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _351_ (.A1(\div_counter[8] ),
    .A2(\div_counter[9] ),
    .A3(_107_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _352_ (.A1(\div_counter[10] ),
    .A2(_108_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _353_ (.A1(_102_),
    .A2(_104_),
    .A3(_109_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _354_ (.A1(net25),
    .A2(\div_counter[0] ),
    .A3(\div_counter[1] ),
    .Z(_110_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _355_ (.A1(\div_counter[2] ),
    .A2(\div_counter[3] ),
    .A3(\div_counter[4] ),
    .A4(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _356_ (.A1(\div_counter[5] ),
    .A2(\div_counter[6] ),
    .A3(\div_counter[7] ),
    .A4(_111_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _357_ (.A1(\div_counter[8] ),
    .A2(\div_counter[9] ),
    .A3(\div_counter[10] ),
    .A4(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _358_ (.A1(\div_counter[11] ),
    .A2(_113_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _359_ (.A1(_102_),
    .A2(_104_),
    .A3(_114_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _360_ (.A1(\div_counter[8] ),
    .A2(\div_counter[9] ),
    .A3(\div_counter[10] ),
    .A4(\div_counter[11] ),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _361_ (.A1(_107_),
    .A2(_115_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _362_ (.A1(\div_counter[12] ),
    .A2(_116_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _363_ (.A1(_102_),
    .A2(_104_),
    .A3(_117_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _364_ (.A1(\div_counter[12] ),
    .A2(_115_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _365_ (.A1(_112_),
    .A2(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _366_ (.A1(\div_counter[13] ),
    .A2(_119_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _367_ (.A1(_102_),
    .A2(_104_),
    .A3(_120_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _368_ (.A1(\div_counter[13] ),
    .A2(_118_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _369_ (.A1(_107_),
    .A2(_121_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _370_ (.A1(\div_counter[14] ),
    .A2(_122_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _371_ (.A1(_102_),
    .A2(_104_),
    .A3(_123_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _372_ (.A1(\div_counter[14] ),
    .A2(_112_),
    .A3(_121_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _373_ (.A1(\div_counter[15] ),
    .A2(_124_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _374_ (.A1(_102_),
    .A2(_104_),
    .A3(_125_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _375_ (.A1(_062_),
    .A2(_210_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _376_ (.A1(_063_),
    .A2(\div_counter[1] ),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _377_ (.A1(_077_),
    .A2(_126_),
    .B(_127_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _378_ (.A1(_102_),
    .A2(_128_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _379_ (.A1(net25),
    .A2(_209_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _380_ (.A1(\div_counter[2] ),
    .A2(_129_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _381_ (.A1(_102_),
    .A2(_104_),
    .A3(_130_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _382_ (.A1(\div_counter[2] ),
    .A2(_110_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _383_ (.A1(\div_counter[3] ),
    .A2(_131_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _384_ (.A1(_102_),
    .A2(_104_),
    .A3(_132_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _385_ (.A1(\div_counter[4] ),
    .A2(_105_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _386_ (.A1(_102_),
    .A2(_104_),
    .A3(_133_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _387_ (.A1(\div_counter[5] ),
    .A2(_111_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _388_ (.A1(_025_),
    .A2(_104_),
    .A3(_134_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _389_ (.A1(\div_counter[5] ),
    .A2(_106_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _390_ (.A1(\div_counter[6] ),
    .A2(_135_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _391_ (.A1(_025_),
    .A2(_103_),
    .A3(_136_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _392_ (.A1(\div_counter[5] ),
    .A2(\div_counter[6] ),
    .A3(_111_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _393_ (.A1(\div_counter[7] ),
    .A2(_137_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _394_ (.A1(_025_),
    .A2(_103_),
    .A3(_138_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _395_ (.A1(\div_counter[8] ),
    .A2(_107_),
    .Z(_139_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _396_ (.A1(_025_),
    .A2(_103_),
    .A3(_139_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _397_ (.A1(\div_counter[8] ),
    .A2(_112_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _398_ (.A1(\div_counter[9] ),
    .A2(_140_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _399_ (.A1(_025_),
    .A2(_103_),
    .A3(_141_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _400_ (.A1(_213_),
    .A2(_216_),
    .A3(_219_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _401_ (.A1(_225_),
    .A2(_231_),
    .A3(_234_),
    .A4(_222_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _402_ (.A1(_228_),
    .A2(_142_),
    .A3(_143_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _403_ (.A1(_027_),
    .A2(_063_),
    .A3(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _404_ (.I(_222_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _405_ (.I(_228_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _406_ (.I(_233_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _407_ (.A1(_231_),
    .A2(_148_),
    .B(_230_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _408_ (.I(_227_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _409_ (.A1(_147_),
    .A2(_149_),
    .B(_150_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _410_ (.A1(_225_),
    .A2(_151_),
    .B(_224_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _411_ (.A1(_216_),
    .A2(_218_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _412_ (.A1(_215_),
    .A2(_153_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _413_ (.A1(_213_),
    .A2(_154_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _414_ (.A1(_212_),
    .A2(_221_),
    .A3(_155_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _415_ (.A1(_146_),
    .A2(_152_),
    .B(_156_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _416_ (.A1(_212_),
    .A2(_142_),
    .A3(_155_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _417_ (.A1(_145_),
    .A2(_157_),
    .A3(_158_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _418_ (.A(net1),
    .B(_159_),
    .CO(_160_),
    .S(_161_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _419_ (.A(_162_),
    .B(\div_counter[1] ),
    .CO(_163_),
    .S(_164_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _420_ (.A(_165_),
    .B(\div_counter[3] ),
    .CO(_166_),
    .S(_167_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _421_ (.A(_168_),
    .B(\div_counter[2] ),
    .CO(_169_),
    .S(_170_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _422_ (.A(_171_),
    .B(\div_counter[7] ),
    .CO(_172_),
    .S(_173_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _423_ (.A(_174_),
    .B(\div_counter[6] ),
    .CO(_175_),
    .S(_176_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _424_ (.A(_177_),
    .B(\div_counter[4] ),
    .CO(_178_),
    .S(_179_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _425_ (.A(_180_),
    .B(\div_counter[5] ),
    .CO(_181_),
    .S(_182_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _426_ (.A(_183_),
    .B(\div_counter[15] ),
    .CO(_184_),
    .S(_185_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _427_ (.A(_186_),
    .B(\div_counter[14] ),
    .CO(_187_),
    .S(_188_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _428_ (.A(_189_),
    .B(\div_counter[13] ),
    .CO(_190_),
    .S(_191_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _429_ (.A(_192_),
    .B(\div_counter[12] ),
    .CO(_193_),
    .S(_194_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _430_ (.A(_195_),
    .B(\div_counter[11] ),
    .CO(_196_),
    .S(_197_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _431_ (.A(_198_),
    .B(\div_counter[10] ),
    .CO(_199_),
    .S(_200_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _432_ (.A(_201_),
    .B(\div_counter[9] ),
    .CO(_202_),
    .S(_203_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _433_ (.A(_204_),
    .B(\div_counter[8] ),
    .CO(_205_),
    .S(_206_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _434_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_207_),
    .S(_208_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _435_ (.A(\div_counter[0] ),
    .B(\div_counter[1] ),
    .CO(_209_),
    .S(_210_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _436_ (.A(_211_),
    .B(net24),
    .CO(_212_),
    .S(_213_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _437_ (.A(_214_),
    .B(net23),
    .CO(_215_),
    .S(_216_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _438_ (.A(_217_),
    .B(net22),
    .CO(_218_),
    .S(_219_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _439_ (.A(_220_),
    .B(net21),
    .CO(_221_),
    .S(_222_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _440_ (.A(_223_),
    .B(net20),
    .CO(_224_),
    .S(_225_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _441_ (.A(_226_),
    .B(net19),
    .CO(_227_),
    .S(_228_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _442_ (.A(_229_),
    .B(net18),
    .CO(_230_),
    .S(_231_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _443_ (.A(\counter[0] ),
    .B(_232_),
    .CO(_233_),
    .S(_234_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[0]$_SDFFE_PN0P_  (.D(_008_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\div_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[10]$_SDFFE_PN0P_  (.D(_009_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[11]$_SDFFE_PN0P_  (.D(_010_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[12]$_SDFFE_PN0P_  (.D(_011_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[13]$_SDFFE_PN0P_  (.D(_012_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[14]$_SDFFE_PN0P_  (.D(_013_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[15]$_SDFFE_PN0P_  (.D(_014_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[1]$_SDFFE_PN0P_  (.D(_015_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[2]$_SDFFE_PN0P_  (.D(_016_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[3]$_SDFFE_PN0P_  (.D(_017_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[4]$_SDFFE_PN0P_  (.D(_018_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[5]$_SDFFE_PN0P_  (.D(_019_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[6]$_SDFFE_PN0P_  (.D(_020_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[7]$_SDFFE_PN0P_  (.D(_021_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[8]$_SDFFE_PN0P_  (.D(_022_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \div_counter[9]$_SDFFE_PN0P_  (.D(_023_),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\div_counter[9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \pwm_reg$_SDFF_PN0_  (.D(_024_),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_84 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_127 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(div[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(div[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(div[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(div[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(div[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(div[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(div[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(div[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(div[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(div[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(div[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(div[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(div[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(div[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(div[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(div[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(duty[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(duty[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(duty[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(duty[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(duty[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(duty[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(duty[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(duty[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input25 (.I(enable),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input26 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net27),
    .Z(pwm_out));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_390 ();
endmodule
