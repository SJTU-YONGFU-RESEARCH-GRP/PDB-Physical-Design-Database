module riscv (clk,
    memread,
    memwrite,
    reset,
    suspend,
    aluout,
    instr,
    pc,
    readdata,
    writedata);
 input clk;
 output memread;
 output memwrite;
 input reset;
 output suspend;
 output [31:0] aluout;
 input [31:0] instr;
 output [31:0] pc;
 input [31:0] readdata;
 output [31:0] writedata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire net250;
 wire _0035_;
 wire net249;
 wire _0037_;
 wire net248;
 wire net247;
 wire net246;
 wire _0041_;
 wire _0042_;
 wire clknet_3_7__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire _0046_;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire _0051_;
 wire clknet_3_0__leaf_clk;
 wire clknet_0_clk;
 wire _0054_;
 wire _0055_;
 wire clknet_leaf_103_clk;
 wire _0057_;
 wire _0058_;
 wire clknet_leaf_102_clk;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire clknet_leaf_101_clk;
 wire _0066_;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_97_clk;
 wire _0071_;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_95_clk;
 wire _0074_;
 wire clknet_leaf_94_clk;
 wire _0076_;
 wire _0077_;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_92_clk;
 wire _0080_;
 wire _0081_;
 wire clknet_leaf_91_clk;
 wire _0083_;
 wire _0084_;
 wire clknet_leaf_90_clk;
 wire _0086_;
 wire clknet_leaf_89_clk;
 wire _0088_;
 wire _0089_;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_87_clk;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire clknet_leaf_86_clk;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire clknet_leaf_85_clk;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire clknet_leaf_84_clk;
 wire _0117_;
 wire clknet_leaf_83_clk;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_81_clk;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire clknet_leaf_80_clk;
 wire _0132_;
 wire _0133_;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_78_clk;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_74_clk;
 wire _0145_;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_72_clk;
 wire _0148_;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_64_clk;
 wire _0157_;
 wire _0158_;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_60_clk;
 wire _0163_;
 wire _0164_;
 wire clknet_leaf_59_clk;
 wire _0166_;
 wire clknet_leaf_58_clk;
 wire _0168_;
 wire clknet_leaf_57_clk;
 wire _0170_;
 wire clknet_leaf_56_clk;
 wire _0172_;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_53_clk;
 wire _0176_;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_49_clk;
 wire _0181_;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_46_clk;
 wire _0185_;
 wire _0186_;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_43_clk;
 wire _0190_;
 wire clknet_leaf_42_clk;
 wire _0192_;
 wire clknet_leaf_41_clk;
 wire _0194_;
 wire _0195_;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_36_clk;
 wire _0201_;
 wire _0202_;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_34_clk;
 wire _0205_;
 wire clknet_leaf_33_clk;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire _0217_;
 wire _0218_;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_27_clk;
 wire _0221_;
 wire clknet_leaf_26_clk;
 wire _0223_;
 wire _0224_;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire _0237_;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire clknet_leaf_17_clk;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire clknet_leaf_16_clk;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire _0266_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire clknet_leaf_11_clk;
 wire _0273_;
 wire _0274_;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire clknet_leaf_4_clk;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire clknet_leaf_1_clk;
 wire net245;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire net244;
 wire net243;
 wire net242;
 wire _0304_;
 wire net241;
 wire net240;
 wire net239;
 wire net238;
 wire _0309_;
 wire net237;
 wire _0311_;
 wire net236;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire net235;
 wire net234;
 wire net233;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire net232;
 wire _0336_;
 wire _0337_;
 wire net231;
 wire _0339_;
 wire _0340_;
 wire net230;
 wire _0342_;
 wire net229;
 wire _0344_;
 wire net228;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire net227;
 wire _0350_;
 wire _0351_;
 wire net226;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire net225;
 wire _0360_;
 wire net224;
 wire net223;
 wire net222;
 wire _0364_;
 wire net221;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire net219;
 wire net218;
 wire net217;
 wire _0376_;
 wire net216;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire net215;
 wire _0382_;
 wire _0383_;
 wire net214;
 wire net213;
 wire net212;
 wire net211;
 wire _0388_;
 wire _0389_;
 wire net210;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire net209;
 wire net208;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire net207;
 wire net206;
 wire net205;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire net204;
 wire _0421_;
 wire _0422_;
 wire net203;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire net202;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire net201;
 wire net200;
 wire _0442_;
 wire net199;
 wire _0444_;
 wire _0445_;
 wire net198;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire net197;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire net196;
 wire _0470_;
 wire _0471_;
 wire net195;
 wire _0473_;
 wire net194;
 wire _0475_;
 wire _0476_;
 wire net193;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire net192;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire net191;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire net190;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire net189;
 wire _0495_;
 wire net188;
 wire net187;
 wire net186;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire net185;
 wire _0503_;
 wire net184;
 wire net183;
 wire _0506_;
 wire _0507_;
 wire net182;
 wire _0509_;
 wire _0510_;
 wire net181;
 wire net180;
 wire _0513_;
 wire _0514_;
 wire net179;
 wire _0516_;
 wire net178;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire net177;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire net176;
 wire _0534_;
 wire _0535_;
 wire net175;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire net174;
 wire _0542_;
 wire net173;
 wire net172;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire net171;
 wire net170;
 wire net169;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire net168;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire net167;
 wire net166;
 wire _0576_;
 wire net165;
 wire _0578_;
 wire net164;
 wire net163;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire net162;
 wire _0585_;
 wire _0586_;
 wire net161;
 wire net160;
 wire net159;
 wire _0590_;
 wire _0591_;
 wire net158;
 wire _0593_;
 wire net157;
 wire _0595_;
 wire net156;
 wire net155;
 wire _0598_;
 wire _0599_;
 wire net154;
 wire _0601_;
 wire _0602_;
 wire net153;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire net152;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire net151;
 wire net150;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire net149;
 wire net148;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire net146;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire net145;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire net144;
 wire _0659_;
 wire _0660_;
 wire net143;
 wire net142;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire net141;
 wire net140;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire net139;
 wire _0673_;
 wire _0674_;
 wire net138;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire net137;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire net136;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire net135;
 wire _0716_;
 wire _0717_;
 wire net134;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire net133;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire net132;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire net131;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire net130;
 wire net129;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire net128;
 wire _0916_;
 wire _0917_;
 wire net127;
 wire _0919_;
 wire _0920_;
 wire net126;
 wire net125;
 wire _0923_;
 wire net124;
 wire net123;
 wire net122;
 wire net121;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire net120;
 wire net119;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire net118;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire net117;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire net116;
 wire net115;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire net114;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire net112;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire net111;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire net110;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire net109;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire net108;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire net107;
 wire net106;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire net105;
 wire _1257_;
 wire net104;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire net103;
 wire net102;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire net101;
 wire net100;
 wire net99;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire net97;
 wire net96;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire net91;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire net90;
 wire _1805_;
 wire _1806_;
 wire net89;
 wire _1808_;
 wire _1809_;
 wire net88;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire net87;
 wire _1820_;
 wire net86;
 wire net85;
 wire _1823_;
 wire _1824_;
 wire net84;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire net83;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire net82;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire net81;
 wire _1859_;
 wire net80;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire net79;
 wire net78;
 wire _1893_;
 wire net77;
 wire net76;
 wire _1896_;
 wire net75;
 wire net74;
 wire net73;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire net72;
 wire net71;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire net70;
 wire net69;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire net68;
 wire net67;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire net66;
 wire net65;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire net64;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire net63;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire net62;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire net61;
 wire net60;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire net59;
 wire net58;
 wire _1959_;
 wire _1960_;
 wire net57;
 wire net55;
 wire net56;
 wire net54;
 wire net53;
 wire _1966_;
 wire _1967_;
 wire net52;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire net51;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire net50;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire net49;
 wire net48;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire net47;
 wire _2005_;
 wire net46;
 wire net45;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire net44;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire net43;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire net42;
 wire _2045_;
 wire _2046_;
 wire net41;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire net40;
 wire net39;
 wire _2071_;
 wire net38;
 wire _2073_;
 wire net37;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire net36;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire net35;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire net34;
 wire _2109_;
 wire _2110_;
 wire net33;
 wire net32;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire net31;
 wire net30;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire net29;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire net28;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire net27;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire net26;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire net25;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire net24;
 wire _2743_;
 wire net23;
 wire net22;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire net21;
 wire _2756_;
 wire net20;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire net19;
 wire _2768_;
 wire net18;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire net17;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire net16;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire net15;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire net14;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire net13;
 wire _3130_;
 wire net12;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire net11;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire net10;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire net9;
 wire net8;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire net7;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire net6;
 wire _3162_;
 wire _3163_;
 wire net5;
 wire net4;
 wire _3166_;
 wire net3;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire net2;
 wire _3173_;
 wire _3174_;
 wire net1;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire clknet_leaf_9_clk;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire net220;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire net147;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire net113;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire net98;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire clknet_leaf_0_clk;
 wire \dp.ISRmux.d0[10] ;
 wire \dp.ISRmux.d0[11] ;
 wire \dp.ISRmux.d0[12] ;
 wire \dp.ISRmux.d0[13] ;
 wire \dp.ISRmux.d0[14] ;
 wire \dp.ISRmux.d0[15] ;
 wire \dp.ISRmux.d0[16] ;
 wire \dp.ISRmux.d0[17] ;
 wire \dp.ISRmux.d0[18] ;
 wire \dp.ISRmux.d0[19] ;
 wire \dp.ISRmux.d0[20] ;
 wire \dp.ISRmux.d0[21] ;
 wire \dp.ISRmux.d0[22] ;
 wire \dp.ISRmux.d0[23] ;
 wire \dp.ISRmux.d0[24] ;
 wire \dp.ISRmux.d0[25] ;
 wire \dp.ISRmux.d0[26] ;
 wire \dp.ISRmux.d0[27] ;
 wire \dp.ISRmux.d0[28] ;
 wire \dp.ISRmux.d0[29] ;
 wire \dp.ISRmux.d0[2] ;
 wire \dp.ISRmux.d0[30] ;
 wire \dp.ISRmux.d0[31] ;
 wire \dp.ISRmux.d0[3] ;
 wire \dp.ISRmux.d0[4] ;
 wire \dp.ISRmux.d0[5] ;
 wire \dp.ISRmux.d0[6] ;
 wire \dp.ISRmux.d0[7] ;
 wire \dp.ISRmux.d0[8] ;
 wire \dp.ISRmux.d0[9] ;
 wire \dp.result2[0] ;
 wire \dp.result2[10] ;
 wire \dp.result2[11] ;
 wire \dp.result2[12] ;
 wire \dp.result2[13] ;
 wire \dp.result2[14] ;
 wire \dp.result2[15] ;
 wire \dp.result2[16] ;
 wire \dp.result2[17] ;
 wire \dp.result2[18] ;
 wire \dp.result2[19] ;
 wire \dp.result2[1] ;
 wire \dp.result2[20] ;
 wire \dp.result2[21] ;
 wire \dp.result2[22] ;
 wire \dp.result2[23] ;
 wire \dp.result2[24] ;
 wire \dp.result2[25] ;
 wire \dp.result2[26] ;
 wire \dp.result2[27] ;
 wire \dp.result2[28] ;
 wire \dp.result2[29] ;
 wire \dp.result2[2] ;
 wire \dp.result2[30] ;
 wire \dp.result2[31] ;
 wire \dp.result2[3] ;
 wire \dp.result2[4] ;
 wire \dp.result2[5] ;
 wire \dp.result2[6] ;
 wire \dp.result2[7] ;
 wire \dp.result2[8] ;
 wire \dp.result2[9] ;
 wire \dp.rf.rf[0][0] ;
 wire \dp.rf.rf[0][10] ;
 wire \dp.rf.rf[0][11] ;
 wire \dp.rf.rf[0][12] ;
 wire \dp.rf.rf[0][13] ;
 wire \dp.rf.rf[0][14] ;
 wire \dp.rf.rf[0][15] ;
 wire \dp.rf.rf[0][18] ;
 wire \dp.rf.rf[0][19] ;
 wire \dp.rf.rf[0][1] ;
 wire \dp.rf.rf[0][20] ;
 wire \dp.rf.rf[0][21] ;
 wire \dp.rf.rf[0][22] ;
 wire \dp.rf.rf[0][23] ;
 wire \dp.rf.rf[0][24] ;
 wire \dp.rf.rf[0][25] ;
 wire \dp.rf.rf[0][26] ;
 wire \dp.rf.rf[0][27] ;
 wire \dp.rf.rf[0][28] ;
 wire \dp.rf.rf[0][29] ;
 wire \dp.rf.rf[0][2] ;
 wire \dp.rf.rf[0][30] ;
 wire \dp.rf.rf[0][31] ;
 wire \dp.rf.rf[0][3] ;
 wire \dp.rf.rf[0][4] ;
 wire \dp.rf.rf[0][5] ;
 wire \dp.rf.rf[0][6] ;
 wire \dp.rf.rf[0][7] ;
 wire \dp.rf.rf[0][8] ;
 wire \dp.rf.rf[0][9] ;
 wire \dp.rf.rf[10][0] ;
 wire \dp.rf.rf[10][10] ;
 wire \dp.rf.rf[10][11] ;
 wire \dp.rf.rf[10][12] ;
 wire \dp.rf.rf[10][13] ;
 wire \dp.rf.rf[10][14] ;
 wire \dp.rf.rf[10][15] ;
 wire \dp.rf.rf[10][16] ;
 wire \dp.rf.rf[10][17] ;
 wire \dp.rf.rf[10][18] ;
 wire \dp.rf.rf[10][19] ;
 wire \dp.rf.rf[10][1] ;
 wire \dp.rf.rf[10][20] ;
 wire \dp.rf.rf[10][21] ;
 wire \dp.rf.rf[10][22] ;
 wire \dp.rf.rf[10][23] ;
 wire \dp.rf.rf[10][24] ;
 wire \dp.rf.rf[10][25] ;
 wire \dp.rf.rf[10][26] ;
 wire \dp.rf.rf[10][27] ;
 wire \dp.rf.rf[10][28] ;
 wire \dp.rf.rf[10][29] ;
 wire \dp.rf.rf[10][2] ;
 wire \dp.rf.rf[10][30] ;
 wire \dp.rf.rf[10][31] ;
 wire \dp.rf.rf[10][3] ;
 wire \dp.rf.rf[10][4] ;
 wire \dp.rf.rf[10][5] ;
 wire \dp.rf.rf[10][6] ;
 wire \dp.rf.rf[10][7] ;
 wire \dp.rf.rf[10][8] ;
 wire \dp.rf.rf[10][9] ;
 wire \dp.rf.rf[11][0] ;
 wire \dp.rf.rf[11][10] ;
 wire \dp.rf.rf[11][11] ;
 wire \dp.rf.rf[11][12] ;
 wire \dp.rf.rf[11][13] ;
 wire \dp.rf.rf[11][14] ;
 wire \dp.rf.rf[11][15] ;
 wire \dp.rf.rf[11][16] ;
 wire \dp.rf.rf[11][17] ;
 wire \dp.rf.rf[11][18] ;
 wire \dp.rf.rf[11][19] ;
 wire \dp.rf.rf[11][1] ;
 wire \dp.rf.rf[11][20] ;
 wire \dp.rf.rf[11][21] ;
 wire \dp.rf.rf[11][22] ;
 wire \dp.rf.rf[11][23] ;
 wire \dp.rf.rf[11][24] ;
 wire \dp.rf.rf[11][25] ;
 wire \dp.rf.rf[11][26] ;
 wire \dp.rf.rf[11][27] ;
 wire \dp.rf.rf[11][28] ;
 wire \dp.rf.rf[11][29] ;
 wire \dp.rf.rf[11][2] ;
 wire \dp.rf.rf[11][30] ;
 wire \dp.rf.rf[11][31] ;
 wire \dp.rf.rf[11][3] ;
 wire \dp.rf.rf[11][4] ;
 wire \dp.rf.rf[11][5] ;
 wire \dp.rf.rf[11][6] ;
 wire \dp.rf.rf[11][7] ;
 wire \dp.rf.rf[11][8] ;
 wire \dp.rf.rf[11][9] ;
 wire \dp.rf.rf[12][0] ;
 wire \dp.rf.rf[12][10] ;
 wire \dp.rf.rf[12][11] ;
 wire \dp.rf.rf[12][12] ;
 wire \dp.rf.rf[12][13] ;
 wire \dp.rf.rf[12][14] ;
 wire \dp.rf.rf[12][15] ;
 wire \dp.rf.rf[12][16] ;
 wire \dp.rf.rf[12][17] ;
 wire \dp.rf.rf[12][18] ;
 wire \dp.rf.rf[12][19] ;
 wire \dp.rf.rf[12][1] ;
 wire \dp.rf.rf[12][20] ;
 wire \dp.rf.rf[12][21] ;
 wire \dp.rf.rf[12][22] ;
 wire \dp.rf.rf[12][23] ;
 wire \dp.rf.rf[12][24] ;
 wire \dp.rf.rf[12][25] ;
 wire \dp.rf.rf[12][26] ;
 wire \dp.rf.rf[12][27] ;
 wire \dp.rf.rf[12][28] ;
 wire \dp.rf.rf[12][29] ;
 wire \dp.rf.rf[12][2] ;
 wire \dp.rf.rf[12][30] ;
 wire \dp.rf.rf[12][31] ;
 wire \dp.rf.rf[12][3] ;
 wire \dp.rf.rf[12][4] ;
 wire \dp.rf.rf[12][5] ;
 wire \dp.rf.rf[12][6] ;
 wire \dp.rf.rf[12][7] ;
 wire \dp.rf.rf[12][8] ;
 wire \dp.rf.rf[12][9] ;
 wire \dp.rf.rf[13][0] ;
 wire \dp.rf.rf[13][10] ;
 wire \dp.rf.rf[13][11] ;
 wire \dp.rf.rf[13][12] ;
 wire \dp.rf.rf[13][13] ;
 wire \dp.rf.rf[13][14] ;
 wire \dp.rf.rf[13][15] ;
 wire \dp.rf.rf[13][16] ;
 wire \dp.rf.rf[13][17] ;
 wire \dp.rf.rf[13][18] ;
 wire \dp.rf.rf[13][19] ;
 wire \dp.rf.rf[13][1] ;
 wire \dp.rf.rf[13][20] ;
 wire \dp.rf.rf[13][21] ;
 wire \dp.rf.rf[13][22] ;
 wire \dp.rf.rf[13][23] ;
 wire \dp.rf.rf[13][24] ;
 wire \dp.rf.rf[13][25] ;
 wire \dp.rf.rf[13][26] ;
 wire \dp.rf.rf[13][27] ;
 wire \dp.rf.rf[13][28] ;
 wire \dp.rf.rf[13][29] ;
 wire \dp.rf.rf[13][2] ;
 wire \dp.rf.rf[13][30] ;
 wire \dp.rf.rf[13][31] ;
 wire \dp.rf.rf[13][3] ;
 wire \dp.rf.rf[13][4] ;
 wire \dp.rf.rf[13][5] ;
 wire \dp.rf.rf[13][6] ;
 wire \dp.rf.rf[13][7] ;
 wire \dp.rf.rf[13][8] ;
 wire \dp.rf.rf[13][9] ;
 wire \dp.rf.rf[14][0] ;
 wire \dp.rf.rf[14][10] ;
 wire \dp.rf.rf[14][11] ;
 wire \dp.rf.rf[14][12] ;
 wire \dp.rf.rf[14][13] ;
 wire \dp.rf.rf[14][14] ;
 wire \dp.rf.rf[14][15] ;
 wire \dp.rf.rf[14][16] ;
 wire \dp.rf.rf[14][17] ;
 wire \dp.rf.rf[14][18] ;
 wire \dp.rf.rf[14][19] ;
 wire \dp.rf.rf[14][1] ;
 wire \dp.rf.rf[14][20] ;
 wire \dp.rf.rf[14][21] ;
 wire \dp.rf.rf[14][22] ;
 wire \dp.rf.rf[14][23] ;
 wire \dp.rf.rf[14][24] ;
 wire \dp.rf.rf[14][25] ;
 wire \dp.rf.rf[14][26] ;
 wire \dp.rf.rf[14][27] ;
 wire \dp.rf.rf[14][28] ;
 wire \dp.rf.rf[14][29] ;
 wire \dp.rf.rf[14][2] ;
 wire \dp.rf.rf[14][30] ;
 wire \dp.rf.rf[14][31] ;
 wire \dp.rf.rf[14][3] ;
 wire \dp.rf.rf[14][4] ;
 wire \dp.rf.rf[14][5] ;
 wire \dp.rf.rf[14][6] ;
 wire \dp.rf.rf[14][7] ;
 wire \dp.rf.rf[14][8] ;
 wire \dp.rf.rf[14][9] ;
 wire \dp.rf.rf[15][0] ;
 wire \dp.rf.rf[15][10] ;
 wire \dp.rf.rf[15][11] ;
 wire \dp.rf.rf[15][12] ;
 wire \dp.rf.rf[15][13] ;
 wire \dp.rf.rf[15][14] ;
 wire \dp.rf.rf[15][15] ;
 wire \dp.rf.rf[15][16] ;
 wire \dp.rf.rf[15][17] ;
 wire \dp.rf.rf[15][18] ;
 wire \dp.rf.rf[15][19] ;
 wire \dp.rf.rf[15][1] ;
 wire \dp.rf.rf[15][20] ;
 wire \dp.rf.rf[15][21] ;
 wire \dp.rf.rf[15][22] ;
 wire \dp.rf.rf[15][23] ;
 wire \dp.rf.rf[15][24] ;
 wire \dp.rf.rf[15][25] ;
 wire \dp.rf.rf[15][26] ;
 wire \dp.rf.rf[15][27] ;
 wire \dp.rf.rf[15][28] ;
 wire \dp.rf.rf[15][29] ;
 wire \dp.rf.rf[15][2] ;
 wire \dp.rf.rf[15][30] ;
 wire \dp.rf.rf[15][31] ;
 wire \dp.rf.rf[15][3] ;
 wire \dp.rf.rf[15][4] ;
 wire \dp.rf.rf[15][5] ;
 wire \dp.rf.rf[15][6] ;
 wire \dp.rf.rf[15][7] ;
 wire \dp.rf.rf[15][8] ;
 wire \dp.rf.rf[15][9] ;
 wire \dp.rf.rf[16][0] ;
 wire \dp.rf.rf[16][10] ;
 wire \dp.rf.rf[16][11] ;
 wire \dp.rf.rf[16][12] ;
 wire \dp.rf.rf[16][13] ;
 wire \dp.rf.rf[16][14] ;
 wire \dp.rf.rf[16][15] ;
 wire \dp.rf.rf[16][16] ;
 wire \dp.rf.rf[16][17] ;
 wire \dp.rf.rf[16][18] ;
 wire \dp.rf.rf[16][19] ;
 wire \dp.rf.rf[16][1] ;
 wire \dp.rf.rf[16][20] ;
 wire \dp.rf.rf[16][21] ;
 wire \dp.rf.rf[16][22] ;
 wire \dp.rf.rf[16][23] ;
 wire \dp.rf.rf[16][24] ;
 wire \dp.rf.rf[16][25] ;
 wire \dp.rf.rf[16][26] ;
 wire \dp.rf.rf[16][27] ;
 wire \dp.rf.rf[16][28] ;
 wire \dp.rf.rf[16][29] ;
 wire \dp.rf.rf[16][2] ;
 wire \dp.rf.rf[16][30] ;
 wire \dp.rf.rf[16][31] ;
 wire \dp.rf.rf[16][3] ;
 wire \dp.rf.rf[16][4] ;
 wire \dp.rf.rf[16][5] ;
 wire \dp.rf.rf[16][6] ;
 wire \dp.rf.rf[16][7] ;
 wire \dp.rf.rf[16][8] ;
 wire \dp.rf.rf[16][9] ;
 wire \dp.rf.rf[17][0] ;
 wire \dp.rf.rf[17][10] ;
 wire \dp.rf.rf[17][11] ;
 wire \dp.rf.rf[17][12] ;
 wire \dp.rf.rf[17][13] ;
 wire \dp.rf.rf[17][14] ;
 wire \dp.rf.rf[17][15] ;
 wire \dp.rf.rf[17][16] ;
 wire \dp.rf.rf[17][17] ;
 wire \dp.rf.rf[17][18] ;
 wire \dp.rf.rf[17][19] ;
 wire \dp.rf.rf[17][1] ;
 wire \dp.rf.rf[17][20] ;
 wire \dp.rf.rf[17][21] ;
 wire \dp.rf.rf[17][22] ;
 wire \dp.rf.rf[17][23] ;
 wire \dp.rf.rf[17][24] ;
 wire \dp.rf.rf[17][25] ;
 wire \dp.rf.rf[17][26] ;
 wire \dp.rf.rf[17][27] ;
 wire \dp.rf.rf[17][28] ;
 wire \dp.rf.rf[17][29] ;
 wire \dp.rf.rf[17][2] ;
 wire \dp.rf.rf[17][30] ;
 wire \dp.rf.rf[17][31] ;
 wire \dp.rf.rf[17][3] ;
 wire \dp.rf.rf[17][4] ;
 wire \dp.rf.rf[17][5] ;
 wire \dp.rf.rf[17][6] ;
 wire \dp.rf.rf[17][7] ;
 wire \dp.rf.rf[17][8] ;
 wire \dp.rf.rf[17][9] ;
 wire \dp.rf.rf[18][0] ;
 wire \dp.rf.rf[18][10] ;
 wire \dp.rf.rf[18][11] ;
 wire \dp.rf.rf[18][12] ;
 wire \dp.rf.rf[18][13] ;
 wire \dp.rf.rf[18][14] ;
 wire \dp.rf.rf[18][15] ;
 wire \dp.rf.rf[18][16] ;
 wire \dp.rf.rf[18][17] ;
 wire \dp.rf.rf[18][18] ;
 wire \dp.rf.rf[18][19] ;
 wire \dp.rf.rf[18][1] ;
 wire \dp.rf.rf[18][20] ;
 wire \dp.rf.rf[18][21] ;
 wire \dp.rf.rf[18][22] ;
 wire \dp.rf.rf[18][23] ;
 wire \dp.rf.rf[18][24] ;
 wire \dp.rf.rf[18][25] ;
 wire \dp.rf.rf[18][26] ;
 wire \dp.rf.rf[18][27] ;
 wire \dp.rf.rf[18][28] ;
 wire \dp.rf.rf[18][29] ;
 wire \dp.rf.rf[18][2] ;
 wire \dp.rf.rf[18][30] ;
 wire \dp.rf.rf[18][31] ;
 wire \dp.rf.rf[18][3] ;
 wire \dp.rf.rf[18][4] ;
 wire \dp.rf.rf[18][5] ;
 wire \dp.rf.rf[18][6] ;
 wire \dp.rf.rf[18][7] ;
 wire \dp.rf.rf[18][8] ;
 wire \dp.rf.rf[18][9] ;
 wire \dp.rf.rf[19][0] ;
 wire \dp.rf.rf[19][10] ;
 wire \dp.rf.rf[19][11] ;
 wire \dp.rf.rf[19][12] ;
 wire \dp.rf.rf[19][13] ;
 wire \dp.rf.rf[19][14] ;
 wire \dp.rf.rf[19][15] ;
 wire \dp.rf.rf[19][16] ;
 wire \dp.rf.rf[19][17] ;
 wire \dp.rf.rf[19][18] ;
 wire \dp.rf.rf[19][19] ;
 wire \dp.rf.rf[19][1] ;
 wire \dp.rf.rf[19][20] ;
 wire \dp.rf.rf[19][21] ;
 wire \dp.rf.rf[19][22] ;
 wire \dp.rf.rf[19][23] ;
 wire \dp.rf.rf[19][24] ;
 wire \dp.rf.rf[19][25] ;
 wire \dp.rf.rf[19][26] ;
 wire \dp.rf.rf[19][27] ;
 wire \dp.rf.rf[19][28] ;
 wire \dp.rf.rf[19][29] ;
 wire \dp.rf.rf[19][2] ;
 wire \dp.rf.rf[19][30] ;
 wire \dp.rf.rf[19][31] ;
 wire \dp.rf.rf[19][3] ;
 wire \dp.rf.rf[19][4] ;
 wire \dp.rf.rf[19][5] ;
 wire \dp.rf.rf[19][6] ;
 wire \dp.rf.rf[19][7] ;
 wire \dp.rf.rf[19][8] ;
 wire \dp.rf.rf[19][9] ;
 wire \dp.rf.rf[1][0] ;
 wire \dp.rf.rf[1][10] ;
 wire \dp.rf.rf[1][11] ;
 wire \dp.rf.rf[1][12] ;
 wire \dp.rf.rf[1][13] ;
 wire \dp.rf.rf[1][14] ;
 wire \dp.rf.rf[1][15] ;
 wire \dp.rf.rf[1][16] ;
 wire \dp.rf.rf[1][17] ;
 wire \dp.rf.rf[1][18] ;
 wire \dp.rf.rf[1][19] ;
 wire \dp.rf.rf[1][1] ;
 wire \dp.rf.rf[1][20] ;
 wire \dp.rf.rf[1][21] ;
 wire \dp.rf.rf[1][22] ;
 wire \dp.rf.rf[1][23] ;
 wire \dp.rf.rf[1][24] ;
 wire \dp.rf.rf[1][25] ;
 wire \dp.rf.rf[1][26] ;
 wire \dp.rf.rf[1][27] ;
 wire \dp.rf.rf[1][28] ;
 wire \dp.rf.rf[1][29] ;
 wire \dp.rf.rf[1][2] ;
 wire \dp.rf.rf[1][30] ;
 wire \dp.rf.rf[1][31] ;
 wire \dp.rf.rf[1][3] ;
 wire \dp.rf.rf[1][4] ;
 wire \dp.rf.rf[1][5] ;
 wire \dp.rf.rf[1][6] ;
 wire \dp.rf.rf[1][7] ;
 wire \dp.rf.rf[1][8] ;
 wire \dp.rf.rf[1][9] ;
 wire \dp.rf.rf[20][0] ;
 wire \dp.rf.rf[20][10] ;
 wire \dp.rf.rf[20][11] ;
 wire \dp.rf.rf[20][12] ;
 wire \dp.rf.rf[20][13] ;
 wire \dp.rf.rf[20][14] ;
 wire \dp.rf.rf[20][15] ;
 wire \dp.rf.rf[20][16] ;
 wire \dp.rf.rf[20][17] ;
 wire \dp.rf.rf[20][18] ;
 wire \dp.rf.rf[20][19] ;
 wire \dp.rf.rf[20][1] ;
 wire \dp.rf.rf[20][20] ;
 wire \dp.rf.rf[20][21] ;
 wire \dp.rf.rf[20][22] ;
 wire \dp.rf.rf[20][23] ;
 wire \dp.rf.rf[20][24] ;
 wire \dp.rf.rf[20][25] ;
 wire \dp.rf.rf[20][26] ;
 wire \dp.rf.rf[20][27] ;
 wire \dp.rf.rf[20][28] ;
 wire \dp.rf.rf[20][29] ;
 wire \dp.rf.rf[20][2] ;
 wire \dp.rf.rf[20][30] ;
 wire \dp.rf.rf[20][31] ;
 wire \dp.rf.rf[20][3] ;
 wire \dp.rf.rf[20][4] ;
 wire \dp.rf.rf[20][5] ;
 wire \dp.rf.rf[20][6] ;
 wire \dp.rf.rf[20][7] ;
 wire \dp.rf.rf[20][8] ;
 wire \dp.rf.rf[20][9] ;
 wire \dp.rf.rf[21][0] ;
 wire \dp.rf.rf[21][10] ;
 wire \dp.rf.rf[21][11] ;
 wire \dp.rf.rf[21][12] ;
 wire \dp.rf.rf[21][13] ;
 wire \dp.rf.rf[21][14] ;
 wire \dp.rf.rf[21][15] ;
 wire \dp.rf.rf[21][16] ;
 wire \dp.rf.rf[21][17] ;
 wire \dp.rf.rf[21][18] ;
 wire \dp.rf.rf[21][19] ;
 wire \dp.rf.rf[21][1] ;
 wire \dp.rf.rf[21][20] ;
 wire \dp.rf.rf[21][21] ;
 wire \dp.rf.rf[21][22] ;
 wire \dp.rf.rf[21][23] ;
 wire \dp.rf.rf[21][24] ;
 wire \dp.rf.rf[21][25] ;
 wire \dp.rf.rf[21][26] ;
 wire \dp.rf.rf[21][27] ;
 wire \dp.rf.rf[21][28] ;
 wire \dp.rf.rf[21][29] ;
 wire \dp.rf.rf[21][2] ;
 wire \dp.rf.rf[21][30] ;
 wire \dp.rf.rf[21][31] ;
 wire \dp.rf.rf[21][3] ;
 wire \dp.rf.rf[21][4] ;
 wire \dp.rf.rf[21][5] ;
 wire \dp.rf.rf[21][6] ;
 wire \dp.rf.rf[21][7] ;
 wire \dp.rf.rf[21][8] ;
 wire \dp.rf.rf[21][9] ;
 wire \dp.rf.rf[22][0] ;
 wire \dp.rf.rf[22][10] ;
 wire \dp.rf.rf[22][11] ;
 wire \dp.rf.rf[22][12] ;
 wire \dp.rf.rf[22][13] ;
 wire \dp.rf.rf[22][14] ;
 wire \dp.rf.rf[22][15] ;
 wire \dp.rf.rf[22][16] ;
 wire \dp.rf.rf[22][17] ;
 wire \dp.rf.rf[22][18] ;
 wire \dp.rf.rf[22][19] ;
 wire \dp.rf.rf[22][1] ;
 wire \dp.rf.rf[22][20] ;
 wire \dp.rf.rf[22][21] ;
 wire \dp.rf.rf[22][22] ;
 wire \dp.rf.rf[22][23] ;
 wire \dp.rf.rf[22][24] ;
 wire \dp.rf.rf[22][25] ;
 wire \dp.rf.rf[22][26] ;
 wire \dp.rf.rf[22][27] ;
 wire \dp.rf.rf[22][28] ;
 wire \dp.rf.rf[22][29] ;
 wire \dp.rf.rf[22][2] ;
 wire \dp.rf.rf[22][30] ;
 wire \dp.rf.rf[22][31] ;
 wire \dp.rf.rf[22][3] ;
 wire \dp.rf.rf[22][4] ;
 wire \dp.rf.rf[22][5] ;
 wire \dp.rf.rf[22][6] ;
 wire \dp.rf.rf[22][7] ;
 wire \dp.rf.rf[22][8] ;
 wire \dp.rf.rf[22][9] ;
 wire \dp.rf.rf[23][0] ;
 wire \dp.rf.rf[23][10] ;
 wire \dp.rf.rf[23][11] ;
 wire \dp.rf.rf[23][12] ;
 wire \dp.rf.rf[23][13] ;
 wire \dp.rf.rf[23][14] ;
 wire \dp.rf.rf[23][15] ;
 wire \dp.rf.rf[23][16] ;
 wire \dp.rf.rf[23][17] ;
 wire \dp.rf.rf[23][18] ;
 wire \dp.rf.rf[23][19] ;
 wire \dp.rf.rf[23][1] ;
 wire \dp.rf.rf[23][20] ;
 wire \dp.rf.rf[23][21] ;
 wire \dp.rf.rf[23][22] ;
 wire \dp.rf.rf[23][23] ;
 wire \dp.rf.rf[23][24] ;
 wire \dp.rf.rf[23][25] ;
 wire \dp.rf.rf[23][26] ;
 wire \dp.rf.rf[23][27] ;
 wire \dp.rf.rf[23][28] ;
 wire \dp.rf.rf[23][29] ;
 wire \dp.rf.rf[23][2] ;
 wire \dp.rf.rf[23][30] ;
 wire \dp.rf.rf[23][31] ;
 wire \dp.rf.rf[23][3] ;
 wire \dp.rf.rf[23][4] ;
 wire \dp.rf.rf[23][5] ;
 wire \dp.rf.rf[23][6] ;
 wire \dp.rf.rf[23][7] ;
 wire \dp.rf.rf[23][8] ;
 wire \dp.rf.rf[23][9] ;
 wire \dp.rf.rf[24][0] ;
 wire \dp.rf.rf[24][10] ;
 wire \dp.rf.rf[24][11] ;
 wire \dp.rf.rf[24][12] ;
 wire \dp.rf.rf[24][13] ;
 wire \dp.rf.rf[24][14] ;
 wire \dp.rf.rf[24][15] ;
 wire \dp.rf.rf[24][16] ;
 wire \dp.rf.rf[24][17] ;
 wire \dp.rf.rf[24][18] ;
 wire \dp.rf.rf[24][19] ;
 wire \dp.rf.rf[24][1] ;
 wire \dp.rf.rf[24][20] ;
 wire \dp.rf.rf[24][21] ;
 wire \dp.rf.rf[24][22] ;
 wire \dp.rf.rf[24][23] ;
 wire \dp.rf.rf[24][24] ;
 wire \dp.rf.rf[24][25] ;
 wire \dp.rf.rf[24][26] ;
 wire \dp.rf.rf[24][27] ;
 wire \dp.rf.rf[24][28] ;
 wire \dp.rf.rf[24][29] ;
 wire \dp.rf.rf[24][2] ;
 wire \dp.rf.rf[24][30] ;
 wire \dp.rf.rf[24][31] ;
 wire \dp.rf.rf[24][3] ;
 wire \dp.rf.rf[24][4] ;
 wire \dp.rf.rf[24][5] ;
 wire \dp.rf.rf[24][6] ;
 wire \dp.rf.rf[24][7] ;
 wire \dp.rf.rf[24][8] ;
 wire \dp.rf.rf[24][9] ;
 wire \dp.rf.rf[25][0] ;
 wire \dp.rf.rf[25][10] ;
 wire \dp.rf.rf[25][11] ;
 wire \dp.rf.rf[25][12] ;
 wire \dp.rf.rf[25][13] ;
 wire \dp.rf.rf[25][14] ;
 wire \dp.rf.rf[25][15] ;
 wire \dp.rf.rf[25][16] ;
 wire \dp.rf.rf[25][17] ;
 wire \dp.rf.rf[25][18] ;
 wire \dp.rf.rf[25][19] ;
 wire \dp.rf.rf[25][1] ;
 wire \dp.rf.rf[25][20] ;
 wire \dp.rf.rf[25][21] ;
 wire \dp.rf.rf[25][22] ;
 wire \dp.rf.rf[25][23] ;
 wire \dp.rf.rf[25][24] ;
 wire \dp.rf.rf[25][25] ;
 wire \dp.rf.rf[25][26] ;
 wire \dp.rf.rf[25][27] ;
 wire \dp.rf.rf[25][28] ;
 wire \dp.rf.rf[25][29] ;
 wire \dp.rf.rf[25][2] ;
 wire \dp.rf.rf[25][30] ;
 wire \dp.rf.rf[25][31] ;
 wire \dp.rf.rf[25][3] ;
 wire \dp.rf.rf[25][4] ;
 wire \dp.rf.rf[25][5] ;
 wire \dp.rf.rf[25][6] ;
 wire \dp.rf.rf[25][7] ;
 wire \dp.rf.rf[25][8] ;
 wire \dp.rf.rf[25][9] ;
 wire \dp.rf.rf[26][0] ;
 wire \dp.rf.rf[26][10] ;
 wire \dp.rf.rf[26][11] ;
 wire \dp.rf.rf[26][12] ;
 wire \dp.rf.rf[26][13] ;
 wire \dp.rf.rf[26][14] ;
 wire \dp.rf.rf[26][15] ;
 wire \dp.rf.rf[26][16] ;
 wire \dp.rf.rf[26][17] ;
 wire \dp.rf.rf[26][18] ;
 wire \dp.rf.rf[26][19] ;
 wire \dp.rf.rf[26][1] ;
 wire \dp.rf.rf[26][20] ;
 wire \dp.rf.rf[26][21] ;
 wire \dp.rf.rf[26][22] ;
 wire \dp.rf.rf[26][23] ;
 wire \dp.rf.rf[26][24] ;
 wire \dp.rf.rf[26][25] ;
 wire \dp.rf.rf[26][26] ;
 wire \dp.rf.rf[26][27] ;
 wire \dp.rf.rf[26][28] ;
 wire \dp.rf.rf[26][29] ;
 wire \dp.rf.rf[26][2] ;
 wire \dp.rf.rf[26][30] ;
 wire \dp.rf.rf[26][31] ;
 wire \dp.rf.rf[26][3] ;
 wire \dp.rf.rf[26][4] ;
 wire \dp.rf.rf[26][5] ;
 wire \dp.rf.rf[26][6] ;
 wire \dp.rf.rf[26][7] ;
 wire \dp.rf.rf[26][8] ;
 wire \dp.rf.rf[26][9] ;
 wire \dp.rf.rf[27][0] ;
 wire \dp.rf.rf[27][10] ;
 wire \dp.rf.rf[27][11] ;
 wire \dp.rf.rf[27][12] ;
 wire \dp.rf.rf[27][13] ;
 wire \dp.rf.rf[27][14] ;
 wire \dp.rf.rf[27][15] ;
 wire \dp.rf.rf[27][16] ;
 wire \dp.rf.rf[27][17] ;
 wire \dp.rf.rf[27][18] ;
 wire \dp.rf.rf[27][19] ;
 wire \dp.rf.rf[27][1] ;
 wire \dp.rf.rf[27][20] ;
 wire \dp.rf.rf[27][21] ;
 wire \dp.rf.rf[27][22] ;
 wire \dp.rf.rf[27][23] ;
 wire \dp.rf.rf[27][24] ;
 wire \dp.rf.rf[27][25] ;
 wire \dp.rf.rf[27][26] ;
 wire \dp.rf.rf[27][27] ;
 wire \dp.rf.rf[27][28] ;
 wire \dp.rf.rf[27][29] ;
 wire \dp.rf.rf[27][2] ;
 wire \dp.rf.rf[27][30] ;
 wire \dp.rf.rf[27][31] ;
 wire \dp.rf.rf[27][3] ;
 wire \dp.rf.rf[27][4] ;
 wire \dp.rf.rf[27][5] ;
 wire \dp.rf.rf[27][6] ;
 wire \dp.rf.rf[27][7] ;
 wire \dp.rf.rf[27][8] ;
 wire \dp.rf.rf[27][9] ;
 wire \dp.rf.rf[28][0] ;
 wire \dp.rf.rf[28][10] ;
 wire \dp.rf.rf[28][11] ;
 wire \dp.rf.rf[28][12] ;
 wire \dp.rf.rf[28][13] ;
 wire \dp.rf.rf[28][14] ;
 wire \dp.rf.rf[28][15] ;
 wire \dp.rf.rf[28][16] ;
 wire \dp.rf.rf[28][17] ;
 wire \dp.rf.rf[28][18] ;
 wire \dp.rf.rf[28][19] ;
 wire \dp.rf.rf[28][1] ;
 wire \dp.rf.rf[28][20] ;
 wire \dp.rf.rf[28][21] ;
 wire \dp.rf.rf[28][22] ;
 wire \dp.rf.rf[28][23] ;
 wire \dp.rf.rf[28][24] ;
 wire \dp.rf.rf[28][25] ;
 wire \dp.rf.rf[28][26] ;
 wire \dp.rf.rf[28][27] ;
 wire \dp.rf.rf[28][28] ;
 wire \dp.rf.rf[28][29] ;
 wire \dp.rf.rf[28][2] ;
 wire \dp.rf.rf[28][30] ;
 wire \dp.rf.rf[28][31] ;
 wire \dp.rf.rf[28][3] ;
 wire \dp.rf.rf[28][4] ;
 wire \dp.rf.rf[28][5] ;
 wire \dp.rf.rf[28][6] ;
 wire \dp.rf.rf[28][7] ;
 wire \dp.rf.rf[28][8] ;
 wire \dp.rf.rf[28][9] ;
 wire \dp.rf.rf[29][0] ;
 wire \dp.rf.rf[29][10] ;
 wire \dp.rf.rf[29][11] ;
 wire \dp.rf.rf[29][12] ;
 wire \dp.rf.rf[29][13] ;
 wire \dp.rf.rf[29][14] ;
 wire \dp.rf.rf[29][15] ;
 wire \dp.rf.rf[29][16] ;
 wire \dp.rf.rf[29][17] ;
 wire \dp.rf.rf[29][18] ;
 wire \dp.rf.rf[29][19] ;
 wire \dp.rf.rf[29][1] ;
 wire \dp.rf.rf[29][20] ;
 wire \dp.rf.rf[29][21] ;
 wire \dp.rf.rf[29][22] ;
 wire \dp.rf.rf[29][23] ;
 wire \dp.rf.rf[29][24] ;
 wire \dp.rf.rf[29][25] ;
 wire \dp.rf.rf[29][26] ;
 wire \dp.rf.rf[29][27] ;
 wire \dp.rf.rf[29][28] ;
 wire \dp.rf.rf[29][29] ;
 wire \dp.rf.rf[29][2] ;
 wire \dp.rf.rf[29][30] ;
 wire \dp.rf.rf[29][31] ;
 wire \dp.rf.rf[29][3] ;
 wire \dp.rf.rf[29][4] ;
 wire \dp.rf.rf[29][5] ;
 wire \dp.rf.rf[29][6] ;
 wire \dp.rf.rf[29][7] ;
 wire \dp.rf.rf[29][8] ;
 wire \dp.rf.rf[29][9] ;
 wire \dp.rf.rf[2][0] ;
 wire \dp.rf.rf[2][10] ;
 wire \dp.rf.rf[2][11] ;
 wire \dp.rf.rf[2][12] ;
 wire \dp.rf.rf[2][13] ;
 wire \dp.rf.rf[2][14] ;
 wire \dp.rf.rf[2][15] ;
 wire \dp.rf.rf[2][16] ;
 wire \dp.rf.rf[2][17] ;
 wire \dp.rf.rf[2][18] ;
 wire \dp.rf.rf[2][19] ;
 wire \dp.rf.rf[2][1] ;
 wire \dp.rf.rf[2][20] ;
 wire \dp.rf.rf[2][21] ;
 wire \dp.rf.rf[2][22] ;
 wire \dp.rf.rf[2][23] ;
 wire \dp.rf.rf[2][24] ;
 wire \dp.rf.rf[2][25] ;
 wire \dp.rf.rf[2][26] ;
 wire \dp.rf.rf[2][27] ;
 wire \dp.rf.rf[2][28] ;
 wire \dp.rf.rf[2][29] ;
 wire \dp.rf.rf[2][2] ;
 wire \dp.rf.rf[2][30] ;
 wire \dp.rf.rf[2][31] ;
 wire \dp.rf.rf[2][3] ;
 wire \dp.rf.rf[2][4] ;
 wire \dp.rf.rf[2][5] ;
 wire \dp.rf.rf[2][6] ;
 wire \dp.rf.rf[2][7] ;
 wire \dp.rf.rf[2][8] ;
 wire \dp.rf.rf[2][9] ;
 wire \dp.rf.rf[30][0] ;
 wire \dp.rf.rf[30][10] ;
 wire \dp.rf.rf[30][11] ;
 wire \dp.rf.rf[30][12] ;
 wire \dp.rf.rf[30][13] ;
 wire \dp.rf.rf[30][14] ;
 wire \dp.rf.rf[30][15] ;
 wire \dp.rf.rf[30][16] ;
 wire \dp.rf.rf[30][17] ;
 wire \dp.rf.rf[30][18] ;
 wire \dp.rf.rf[30][19] ;
 wire \dp.rf.rf[30][1] ;
 wire \dp.rf.rf[30][20] ;
 wire \dp.rf.rf[30][21] ;
 wire \dp.rf.rf[30][22] ;
 wire \dp.rf.rf[30][23] ;
 wire \dp.rf.rf[30][24] ;
 wire \dp.rf.rf[30][25] ;
 wire \dp.rf.rf[30][26] ;
 wire \dp.rf.rf[30][27] ;
 wire \dp.rf.rf[30][28] ;
 wire \dp.rf.rf[30][29] ;
 wire \dp.rf.rf[30][2] ;
 wire \dp.rf.rf[30][30] ;
 wire \dp.rf.rf[30][31] ;
 wire \dp.rf.rf[30][3] ;
 wire \dp.rf.rf[30][4] ;
 wire \dp.rf.rf[30][5] ;
 wire \dp.rf.rf[30][6] ;
 wire \dp.rf.rf[30][7] ;
 wire \dp.rf.rf[30][8] ;
 wire \dp.rf.rf[30][9] ;
 wire \dp.rf.rf[31][0] ;
 wire \dp.rf.rf[31][10] ;
 wire \dp.rf.rf[31][11] ;
 wire \dp.rf.rf[31][12] ;
 wire \dp.rf.rf[31][13] ;
 wire \dp.rf.rf[31][14] ;
 wire \dp.rf.rf[31][15] ;
 wire \dp.rf.rf[31][16] ;
 wire \dp.rf.rf[31][17] ;
 wire \dp.rf.rf[31][18] ;
 wire \dp.rf.rf[31][19] ;
 wire \dp.rf.rf[31][1] ;
 wire \dp.rf.rf[31][20] ;
 wire \dp.rf.rf[31][21] ;
 wire \dp.rf.rf[31][22] ;
 wire \dp.rf.rf[31][23] ;
 wire \dp.rf.rf[31][24] ;
 wire \dp.rf.rf[31][25] ;
 wire \dp.rf.rf[31][26] ;
 wire \dp.rf.rf[31][27] ;
 wire \dp.rf.rf[31][28] ;
 wire \dp.rf.rf[31][29] ;
 wire \dp.rf.rf[31][2] ;
 wire \dp.rf.rf[31][30] ;
 wire \dp.rf.rf[31][31] ;
 wire \dp.rf.rf[31][3] ;
 wire \dp.rf.rf[31][4] ;
 wire \dp.rf.rf[31][5] ;
 wire \dp.rf.rf[31][6] ;
 wire \dp.rf.rf[31][7] ;
 wire \dp.rf.rf[31][8] ;
 wire \dp.rf.rf[31][9] ;
 wire \dp.rf.rf[3][0] ;
 wire \dp.rf.rf[3][10] ;
 wire \dp.rf.rf[3][11] ;
 wire \dp.rf.rf[3][12] ;
 wire \dp.rf.rf[3][13] ;
 wire \dp.rf.rf[3][14] ;
 wire \dp.rf.rf[3][15] ;
 wire \dp.rf.rf[3][16] ;
 wire \dp.rf.rf[3][17] ;
 wire \dp.rf.rf[3][18] ;
 wire \dp.rf.rf[3][19] ;
 wire \dp.rf.rf[3][1] ;
 wire \dp.rf.rf[3][20] ;
 wire \dp.rf.rf[3][21] ;
 wire \dp.rf.rf[3][22] ;
 wire \dp.rf.rf[3][23] ;
 wire \dp.rf.rf[3][24] ;
 wire \dp.rf.rf[3][25] ;
 wire \dp.rf.rf[3][26] ;
 wire \dp.rf.rf[3][27] ;
 wire \dp.rf.rf[3][28] ;
 wire \dp.rf.rf[3][29] ;
 wire \dp.rf.rf[3][2] ;
 wire \dp.rf.rf[3][30] ;
 wire \dp.rf.rf[3][31] ;
 wire \dp.rf.rf[3][3] ;
 wire \dp.rf.rf[3][4] ;
 wire \dp.rf.rf[3][5] ;
 wire \dp.rf.rf[3][6] ;
 wire \dp.rf.rf[3][7] ;
 wire \dp.rf.rf[3][8] ;
 wire \dp.rf.rf[3][9] ;
 wire \dp.rf.rf[4][0] ;
 wire \dp.rf.rf[4][10] ;
 wire \dp.rf.rf[4][11] ;
 wire \dp.rf.rf[4][12] ;
 wire \dp.rf.rf[4][13] ;
 wire \dp.rf.rf[4][14] ;
 wire \dp.rf.rf[4][15] ;
 wire \dp.rf.rf[4][16] ;
 wire \dp.rf.rf[4][17] ;
 wire \dp.rf.rf[4][18] ;
 wire \dp.rf.rf[4][19] ;
 wire \dp.rf.rf[4][1] ;
 wire \dp.rf.rf[4][20] ;
 wire \dp.rf.rf[4][21] ;
 wire \dp.rf.rf[4][22] ;
 wire \dp.rf.rf[4][23] ;
 wire \dp.rf.rf[4][24] ;
 wire \dp.rf.rf[4][25] ;
 wire \dp.rf.rf[4][26] ;
 wire \dp.rf.rf[4][27] ;
 wire \dp.rf.rf[4][28] ;
 wire \dp.rf.rf[4][29] ;
 wire \dp.rf.rf[4][2] ;
 wire \dp.rf.rf[4][30] ;
 wire \dp.rf.rf[4][31] ;
 wire \dp.rf.rf[4][3] ;
 wire \dp.rf.rf[4][4] ;
 wire \dp.rf.rf[4][5] ;
 wire \dp.rf.rf[4][6] ;
 wire \dp.rf.rf[4][7] ;
 wire \dp.rf.rf[4][8] ;
 wire \dp.rf.rf[4][9] ;
 wire \dp.rf.rf[5][0] ;
 wire \dp.rf.rf[5][10] ;
 wire \dp.rf.rf[5][11] ;
 wire \dp.rf.rf[5][12] ;
 wire \dp.rf.rf[5][13] ;
 wire \dp.rf.rf[5][14] ;
 wire \dp.rf.rf[5][15] ;
 wire \dp.rf.rf[5][16] ;
 wire \dp.rf.rf[5][17] ;
 wire \dp.rf.rf[5][18] ;
 wire \dp.rf.rf[5][19] ;
 wire \dp.rf.rf[5][1] ;
 wire \dp.rf.rf[5][20] ;
 wire \dp.rf.rf[5][21] ;
 wire \dp.rf.rf[5][22] ;
 wire \dp.rf.rf[5][23] ;
 wire \dp.rf.rf[5][24] ;
 wire \dp.rf.rf[5][25] ;
 wire \dp.rf.rf[5][26] ;
 wire \dp.rf.rf[5][27] ;
 wire \dp.rf.rf[5][28] ;
 wire \dp.rf.rf[5][29] ;
 wire \dp.rf.rf[5][2] ;
 wire \dp.rf.rf[5][30] ;
 wire \dp.rf.rf[5][31] ;
 wire \dp.rf.rf[5][3] ;
 wire \dp.rf.rf[5][4] ;
 wire \dp.rf.rf[5][5] ;
 wire \dp.rf.rf[5][6] ;
 wire \dp.rf.rf[5][7] ;
 wire \dp.rf.rf[5][8] ;
 wire \dp.rf.rf[5][9] ;
 wire \dp.rf.rf[6][0] ;
 wire \dp.rf.rf[6][10] ;
 wire \dp.rf.rf[6][11] ;
 wire \dp.rf.rf[6][12] ;
 wire \dp.rf.rf[6][13] ;
 wire \dp.rf.rf[6][14] ;
 wire \dp.rf.rf[6][15] ;
 wire \dp.rf.rf[6][16] ;
 wire \dp.rf.rf[6][17] ;
 wire \dp.rf.rf[6][18] ;
 wire \dp.rf.rf[6][19] ;
 wire \dp.rf.rf[6][1] ;
 wire \dp.rf.rf[6][20] ;
 wire \dp.rf.rf[6][21] ;
 wire \dp.rf.rf[6][22] ;
 wire \dp.rf.rf[6][23] ;
 wire \dp.rf.rf[6][24] ;
 wire \dp.rf.rf[6][25] ;
 wire \dp.rf.rf[6][26] ;
 wire \dp.rf.rf[6][27] ;
 wire \dp.rf.rf[6][28] ;
 wire \dp.rf.rf[6][29] ;
 wire \dp.rf.rf[6][2] ;
 wire \dp.rf.rf[6][30] ;
 wire \dp.rf.rf[6][31] ;
 wire \dp.rf.rf[6][3] ;
 wire \dp.rf.rf[6][4] ;
 wire \dp.rf.rf[6][5] ;
 wire \dp.rf.rf[6][6] ;
 wire \dp.rf.rf[6][7] ;
 wire \dp.rf.rf[6][8] ;
 wire \dp.rf.rf[6][9] ;
 wire \dp.rf.rf[7][0] ;
 wire \dp.rf.rf[7][10] ;
 wire \dp.rf.rf[7][11] ;
 wire \dp.rf.rf[7][12] ;
 wire \dp.rf.rf[7][13] ;
 wire \dp.rf.rf[7][14] ;
 wire \dp.rf.rf[7][15] ;
 wire \dp.rf.rf[7][16] ;
 wire \dp.rf.rf[7][17] ;
 wire \dp.rf.rf[7][18] ;
 wire \dp.rf.rf[7][19] ;
 wire \dp.rf.rf[7][1] ;
 wire \dp.rf.rf[7][20] ;
 wire \dp.rf.rf[7][21] ;
 wire \dp.rf.rf[7][22] ;
 wire \dp.rf.rf[7][23] ;
 wire \dp.rf.rf[7][24] ;
 wire \dp.rf.rf[7][25] ;
 wire \dp.rf.rf[7][26] ;
 wire \dp.rf.rf[7][27] ;
 wire \dp.rf.rf[7][28] ;
 wire \dp.rf.rf[7][29] ;
 wire \dp.rf.rf[7][2] ;
 wire \dp.rf.rf[7][30] ;
 wire \dp.rf.rf[7][31] ;
 wire \dp.rf.rf[7][3] ;
 wire \dp.rf.rf[7][4] ;
 wire \dp.rf.rf[7][5] ;
 wire \dp.rf.rf[7][6] ;
 wire \dp.rf.rf[7][7] ;
 wire \dp.rf.rf[7][8] ;
 wire \dp.rf.rf[7][9] ;
 wire \dp.rf.rf[8][0] ;
 wire \dp.rf.rf[8][10] ;
 wire \dp.rf.rf[8][11] ;
 wire \dp.rf.rf[8][12] ;
 wire \dp.rf.rf[8][13] ;
 wire \dp.rf.rf[8][14] ;
 wire \dp.rf.rf[8][15] ;
 wire \dp.rf.rf[8][16] ;
 wire \dp.rf.rf[8][17] ;
 wire \dp.rf.rf[8][18] ;
 wire \dp.rf.rf[8][19] ;
 wire \dp.rf.rf[8][1] ;
 wire \dp.rf.rf[8][20] ;
 wire \dp.rf.rf[8][21] ;
 wire \dp.rf.rf[8][22] ;
 wire \dp.rf.rf[8][23] ;
 wire \dp.rf.rf[8][24] ;
 wire \dp.rf.rf[8][25] ;
 wire \dp.rf.rf[8][26] ;
 wire \dp.rf.rf[8][27] ;
 wire \dp.rf.rf[8][28] ;
 wire \dp.rf.rf[8][29] ;
 wire \dp.rf.rf[8][2] ;
 wire \dp.rf.rf[8][30] ;
 wire \dp.rf.rf[8][31] ;
 wire \dp.rf.rf[8][3] ;
 wire \dp.rf.rf[8][4] ;
 wire \dp.rf.rf[8][5] ;
 wire \dp.rf.rf[8][6] ;
 wire \dp.rf.rf[8][7] ;
 wire \dp.rf.rf[8][8] ;
 wire \dp.rf.rf[8][9] ;
 wire \dp.rf.rf[9][0] ;
 wire \dp.rf.rf[9][10] ;
 wire \dp.rf.rf[9][11] ;
 wire \dp.rf.rf[9][12] ;
 wire \dp.rf.rf[9][13] ;
 wire \dp.rf.rf[9][14] ;
 wire \dp.rf.rf[9][15] ;
 wire \dp.rf.rf[9][16] ;
 wire \dp.rf.rf[9][17] ;
 wire \dp.rf.rf[9][18] ;
 wire \dp.rf.rf[9][19] ;
 wire \dp.rf.rf[9][1] ;
 wire \dp.rf.rf[9][20] ;
 wire \dp.rf.rf[9][21] ;
 wire \dp.rf.rf[9][22] ;
 wire \dp.rf.rf[9][23] ;
 wire \dp.rf.rf[9][24] ;
 wire \dp.rf.rf[9][25] ;
 wire \dp.rf.rf[9][26] ;
 wire \dp.rf.rf[9][27] ;
 wire \dp.rf.rf[9][28] ;
 wire \dp.rf.rf[9][29] ;
 wire \dp.rf.rf[9][2] ;
 wire \dp.rf.rf[9][30] ;
 wire \dp.rf.rf[9][31] ;
 wire \dp.rf.rf[9][3] ;
 wire \dp.rf.rf[9][4] ;
 wire \dp.rf.rf[9][5] ;
 wire \dp.rf.rf[9][6] ;
 wire \dp.rf.rf[9][7] ;
 wire \dp.rf.rf[9][8] ;
 wire \dp.rf.rf[9][9] ;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net275;
 wire net276;
 wire net280;
 wire net284;
 wire net288;
 wire net301;
 wire net308;
 wire net309;
 wire net358;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net465;
 wire net466;
 wire net474;
 wire net475;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net530;
 wire net531;
 wire net587;
 wire net588;
 wire net304;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net617;
 wire net625;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net648;
 wire net649;
 wire net650;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net678;
 wire net686;
 wire net687;
 wire net688;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net272;
 wire net273;
 wire net274;
 wire net277;
 wire net278;
 wire net279;
 wire net305;
 wire net321;
 wire net492;
 wire net493;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net613;
 wire net614;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net742;
 wire net814;
 wire net815;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net906;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;

 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_363 ();
 sky130_fd_sc_hd__inv_1 _3654_ (.A(net29),
    .Y(_0035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_362 ();
 sky130_fd_sc_hd__nand2b_2 _3656_ (.A_N(net27),
    .B(net28),
    .Y(_0037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_359 ();
 sky130_fd_sc_hd__and4bb_4 _3660_ (.A_N(net26),
    .B_N(net23),
    .C(net1),
    .D(net12),
    .X(_0041_));
 sky130_fd_sc_hd__nor2b_4 _3661_ (.A(_0037_),
    .B_N(_0041_),
    .Y(_0042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_358 ();
 sky130_fd_sc_hd__and2_4 _3663_ (.A(_0035_),
    .B(_0042_),
    .X(net99));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_356 ();
 sky130_fd_sc_hd__nor2_8 _3666_ (.A(net17),
    .B(net15),
    .Y(_0046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_352 ();
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(\dp.rf.rf[1][0] ),
    .B(net212),
    .Y(_0051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_350 ();
 sky130_fd_sc_hd__nor2_8 _3674_ (.A(net274),
    .B(net16),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _3675_ (.A(_0051_),
    .B(_0054_),
    .Y(_0055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_349 ();
 sky130_fd_sc_hd__clkinvlp_4 _3677_ (.A(net274),
    .Y(_0057_));
 sky130_fd_sc_hd__mux4_2 _3678_ (.A0(\dp.rf.rf[2][0] ),
    .A1(\dp.rf.rf[3][0] ),
    .A2(\dp.rf.rf[10][0] ),
    .A3(\dp.rf.rf[11][0] ),
    .S0(net212),
    .S1(net16),
    .X(_0058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_348 ();
 sky130_fd_sc_hd__mux2i_1 _3680_ (.A0(\dp.rf.rf[8][0] ),
    .A1(\dp.rf.rf[9][0] ),
    .S(net212),
    .Y(_0060_));
 sky130_fd_sc_hd__nor2b_4 _3681_ (.A(net274),
    .B_N(net16),
    .Y(_0061_));
 sky130_fd_sc_hd__a2bb2oi_2 _3682_ (.A1_N(_0057_),
    .A2_N(_0058_),
    .B1(_0060_),
    .B2(_0061_),
    .Y(_0062_));
 sky130_fd_sc_hd__and3_4 _3683_ (.A(_0046_),
    .B(_0055_),
    .C(_0062_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2b_4 _3684_ (.A_N(net17),
    .B(net15),
    .Y(_0064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_347 ();
 sky130_fd_sc_hd__and2_4 _3686_ (.A(net274),
    .B(net16),
    .X(_0066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_343 ();
 sky130_fd_sc_hd__mux2i_1 _3691_ (.A0(\dp.rf.rf[14][0] ),
    .A1(\dp.rf.rf[15][0] ),
    .S(net212),
    .Y(_0071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_341 ();
 sky130_fd_sc_hd__mux2i_1 _3694_ (.A0(\dp.rf.rf[12][0] ),
    .A1(\dp.rf.rf[13][0] ),
    .S(net212),
    .Y(_0074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_340 ();
 sky130_fd_sc_hd__a22oi_1 _3696_ (.A1(_0066_),
    .A2(_0071_),
    .B1(_0074_),
    .B2(_0061_),
    .Y(_0076_));
 sky130_fd_sc_hd__mux2i_1 _3697_ (.A0(\dp.rf.rf[4][0] ),
    .A1(\dp.rf.rf[5][0] ),
    .S(net212),
    .Y(_0077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_338 ();
 sky130_fd_sc_hd__mux2i_1 _3700_ (.A0(\dp.rf.rf[6][0] ),
    .A1(\dp.rf.rf[7][0] ),
    .S(net212),
    .Y(_0080_));
 sky130_fd_sc_hd__nor2b_4 _3701_ (.A(net16),
    .B_N(net274),
    .Y(_0081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_337 ();
 sky130_fd_sc_hd__a22oi_1 _3703_ (.A1(_0054_),
    .A2(_0077_),
    .B1(_0080_),
    .B2(_0081_),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _3704_ (.A(_0076_),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_336 ();
 sky130_fd_sc_hd__clkinv_16 _3706_ (.A(net17),
    .Y(_0086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_335 ();
 sky130_fd_sc_hd__nor2_4 _3708_ (.A(_0086_),
    .B(net15),
    .Y(_0088_));
 sky130_fd_sc_hd__mux2i_1 _3709_ (.A0(\dp.rf.rf[26][0] ),
    .A1(\dp.rf.rf[27][0] ),
    .S(net212),
    .Y(_0089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_333 ();
 sky130_fd_sc_hd__mux2i_1 _3712_ (.A0(\dp.rf.rf[24][0] ),
    .A1(\dp.rf.rf[25][0] ),
    .S(net212),
    .Y(_0092_));
 sky130_fd_sc_hd__a22oi_1 _3713_ (.A1(_0066_),
    .A2(_0089_),
    .B1(_0092_),
    .B2(_0061_),
    .Y(_0093_));
 sky130_fd_sc_hd__mux2i_1 _3714_ (.A0(\dp.rf.rf[18][0] ),
    .A1(\dp.rf.rf[19][0] ),
    .S(net212),
    .Y(_0094_));
 sky130_fd_sc_hd__mux2i_1 _3715_ (.A0(\dp.rf.rf[16][0] ),
    .A1(\dp.rf.rf[17][0] ),
    .S(net212),
    .Y(_0095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_332 ();
 sky130_fd_sc_hd__a22oi_1 _3717_ (.A1(_0081_),
    .A2(_0094_),
    .B1(_0095_),
    .B2(_0054_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand3_1 _3718_ (.A(_0088_),
    .B(_0093_),
    .C(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__o21ai_2 _3719_ (.A1(_0064_),
    .A2(_0084_),
    .B1(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__mux4_2 _3720_ (.A0(\dp.rf.rf[20][0] ),
    .A1(\dp.rf.rf[21][0] ),
    .A2(\dp.rf.rf[22][0] ),
    .A3(\dp.rf.rf[23][0] ),
    .S0(net212),
    .S1(net274),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_2 _3721_ (.A(net17),
    .B(net15),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_4 _3722_ (.A(net16),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__clkinv_16 _3723_ (.A(net16),
    .Y(_0103_));
 sky130_fd_sc_hd__nor2_4 _3724_ (.A(_0103_),
    .B(_0101_),
    .Y(_0104_));
 sky130_fd_sc_hd__mux4_2 _3725_ (.A0(\dp.rf.rf[28][0] ),
    .A1(\dp.rf.rf[29][0] ),
    .A2(\dp.rf.rf[30][0] ),
    .A3(\dp.rf.rf[31][0] ),
    .S0(net212),
    .S1(net274),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _3726_ (.A1(_0100_),
    .A2(_0102_),
    .B1(_0104_),
    .B2(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__or3_4 _3727_ (.A(_0063_),
    .B(_0099_),
    .C(_0106_),
    .X(net133));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_331 ();
 sky130_fd_sc_hd__nand2_4 _3729_ (.A(_0035_),
    .B(_0041_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_2 _3730_ (.A(net4),
    .B(net5),
    .Y(_0109_));
 sky130_fd_sc_hd__nand3_1 _3731_ (.A(net28),
    .B(net24),
    .C(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _3732_ (.A(net28),
    .B(net24),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _3733_ (.A(net5),
    .B(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__o21ai_0 _3734_ (.A1(_0108_),
    .A2(_0110_),
    .B1(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hd__a22oi_1 _3735_ (.A1(net5),
    .A2(_0108_),
    .B1(_0113_),
    .B2(net27),
    .Y(_0114_));
 sky130_fd_sc_hd__and3_4 _3736_ (.A(net1),
    .B(net12),
    .C(net23),
    .X(_0115_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_330 ();
 sky130_fd_sc_hd__nor3b_4 _3738_ (.A(net26),
    .B(net29),
    .C_N(net27),
    .Y(_0117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_329 ();
 sky130_fd_sc_hd__nand2_8 _3740_ (.A(_0115_),
    .B(_0117_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_8 _3741_ (.A(net29),
    .B(_0042_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2_4 _3742_ (.A(_0119_),
    .B(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__or3_4 _3743_ (.A(net6),
    .B(_0114_),
    .C(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_327 ();
 sky130_fd_sc_hd__o21ai_2 _3746_ (.A1(net28),
    .A2(net29),
    .B1(_0037_),
    .Y(_0125_));
 sky130_fd_sc_hd__nand3_4 _3747_ (.A(net1),
    .B(net12),
    .C(net23),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _3748_ (.A(net28),
    .B(net29),
    .Y(_0127_));
 sky130_fd_sc_hd__nor3_4 _3749_ (.A(net27),
    .B(_0126_),
    .C(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__or3b_4 _3750_ (.A(net26),
    .B(net29),
    .C_N(net27),
    .X(_0129_));
 sky130_fd_sc_hd__nor2_8 _3751_ (.A(_0126_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_326 ();
 sky130_fd_sc_hd__a211oi_4 _3753_ (.A1(_0041_),
    .A2(_0125_),
    .B1(net202),
    .C1(_0130_),
    .Y(_0132_));
 sky130_fd_sc_hd__and2_4 _3754_ (.A(net26),
    .B(_0128_),
    .X(_0133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_324 ();
 sky130_fd_sc_hd__nor2b_1 _3757_ (.A(net29),
    .B_N(net30),
    .Y(_0136_));
 sky130_fd_sc_hd__mux2i_2 _3758_ (.A0(net13),
    .A1(_0136_),
    .S(_0042_),
    .Y(_0137_));
 sky130_fd_sc_hd__nor3_4 _3759_ (.A(_0130_),
    .B(_0133_),
    .C(_0137_),
    .Y(_3530_));
 sky130_fd_sc_hd__a211o_4 _3760_ (.A1(_0041_),
    .A2(_0125_),
    .B1(net202),
    .C1(_0130_),
    .X(_0138_));
 sky130_fd_sc_hd__or3_4 _3761_ (.A(_0106_),
    .B(_0063_),
    .C(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__o22a_4 _3762_ (.A1(net179),
    .A2(_3530_),
    .B1(_0139_),
    .B2(_0099_),
    .X(_0140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_321 ();
 sky130_fd_sc_hd__xnor2_1 _3766_ (.A(_0122_),
    .B(_0140_),
    .Y(_3276_));
 sky130_fd_sc_hd__inv_1 _3767_ (.A(_3276_),
    .Y(_3280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_320 ();
 sky130_fd_sc_hd__inv_8 _3769_ (.A(net10),
    .Y(_0145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_318 ();
 sky130_fd_sc_hd__clkinv_16 _3772_ (.A(net208),
    .Y(_0148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_310 ();
 sky130_fd_sc_hd__mux4_1 _3781_ (.A0(\dp.rf.rf[16][0] ),
    .A1(\dp.rf.rf[17][0] ),
    .A2(\dp.rf.rf[18][0] ),
    .A3(\dp.rf.rf[19][0] ),
    .S0(net209),
    .S1(net8),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _3782_ (.A(_0148_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_306 ();
 sky130_fd_sc_hd__mux4_1 _3787_ (.A0(\dp.rf.rf[20][0] ),
    .A1(\dp.rf.rf[21][0] ),
    .A2(\dp.rf.rf[22][0] ),
    .A3(\dp.rf.rf[23][0] ),
    .S0(net209),
    .S1(net8),
    .X(_0163_));
 sky130_fd_sc_hd__nand2_1 _3788_ (.A(net206),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_305 ();
 sky130_fd_sc_hd__nand2_8 _3790_ (.A(net11),
    .B(_0119_),
    .Y(_0166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_304 ();
 sky130_fd_sc_hd__a31oi_2 _3792_ (.A1(_0145_),
    .A2(_0158_),
    .A3(_0164_),
    .B1(_0166_),
    .Y(_0168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_303 ();
 sky130_fd_sc_hd__or2_4 _3794_ (.A(net211),
    .B(net8),
    .X(_0170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_302 ();
 sky130_fd_sc_hd__a21oi_1 _3796_ (.A1(_0119_),
    .A2(_0170_),
    .B1(\dp.rf.rf[24][0] ),
    .Y(_0172_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_299 ();
 sky130_fd_sc_hd__o21ai_4 _3800_ (.A1(_0126_),
    .A2(_0129_),
    .B1(net210),
    .Y(_0176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_295 ();
 sky130_fd_sc_hd__mux2i_1 _3805_ (.A0(\dp.rf.rf[26][0] ),
    .A1(\dp.rf.rf[27][0] ),
    .S(net209),
    .Y(_0181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_292 ();
 sky130_fd_sc_hd__a21oi_1 _3809_ (.A1(net8),
    .A2(_0181_),
    .B1(net206),
    .Y(_0185_));
 sky130_fd_sc_hd__o31ai_1 _3810_ (.A1(\dp.rf.rf[25][0] ),
    .A2(net8),
    .A3(_0176_),
    .B1(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_289 ();
 sky130_fd_sc_hd__mux4_1 _3814_ (.A0(\dp.rf.rf[28][0] ),
    .A1(\dp.rf.rf[29][0] ),
    .A2(\dp.rf.rf[30][0] ),
    .A3(\dp.rf.rf[31][0] ),
    .S0(net209),
    .S1(net8),
    .X(_0190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_288 ();
 sky130_fd_sc_hd__o21ai_4 _3816_ (.A1(_0126_),
    .A2(_0129_),
    .B1(net10),
    .Y(_0192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__a21oi_1 _3818_ (.A1(net206),
    .A2(_0190_),
    .B1(net199),
    .Y(_0194_));
 sky130_fd_sc_hd__o21ai_1 _3819_ (.A1(_0172_),
    .A2(_0186_),
    .B1(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__mux4_1 _3825_ (.A0(\dp.rf.rf[2][0] ),
    .A1(\dp.rf.rf[3][0] ),
    .A2(\dp.rf.rf[6][0] ),
    .A3(\dp.rf.rf[7][0] ),
    .S0(net209),
    .S1(net206),
    .X(_0201_));
 sky130_fd_sc_hd__o21ai_4 _3826_ (.A1(_0126_),
    .A2(_0129_),
    .B1(_0145_),
    .Y(_0202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__nor2_1 _3829_ (.A(_0201_),
    .B(net196),
    .Y(_0205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__mux4_1 _3831_ (.A0(\dp.rf.rf[0][0] ),
    .A1(\dp.rf.rf[1][0] ),
    .A2(\dp.rf.rf[4][0] ),
    .A3(\dp.rf.rf[5][0] ),
    .S0(net209),
    .S1(net206),
    .X(_0207_));
 sky130_fd_sc_hd__nor4_2 _3832_ (.A(net210),
    .B(net8),
    .C(net208),
    .D(net10),
    .Y(_0208_));
 sky130_fd_sc_hd__a211oi_4 _3833_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0208_),
    .C1(net11),
    .Y(_0209_));
 sky130_fd_sc_hd__o31ai_2 _3834_ (.A1(net8),
    .A2(net10),
    .A3(_0207_),
    .B1(net194),
    .Y(_0210_));
 sky130_fd_sc_hd__a21oi_2 _3835_ (.A1(net8),
    .A2(_0205_),
    .B1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__o21ai_4 _3836_ (.A1(_0126_),
    .A2(_0129_),
    .B1(net8),
    .Y(_0212_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__nor2b_1 _3841_ (.A(net209),
    .B_N(\dp.rf.rf[14][0] ),
    .Y(_0217_));
 sky130_fd_sc_hd__a211oi_1 _3842_ (.A1(\dp.rf.rf[15][0] ),
    .A2(net209),
    .B1(_0148_),
    .C1(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__a21oi_4 _3845_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0148_),
    .Y(_0221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__a221oi_2 _3847_ (.A1(net268),
    .A2(net209),
    .B1(_0176_),
    .B2(net269),
    .C1(_0221_),
    .Y(_0223_));
 sky130_fd_sc_hd__clkinv_16 _3848_ (.A(net8),
    .Y(_0224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__mux4_1 _3852_ (.A0(\dp.rf.rf[8][0] ),
    .A1(\dp.rf.rf[9][0] ),
    .A2(\dp.rf.rf[12][0] ),
    .A3(\dp.rf.rf[13][0] ),
    .S0(net209),
    .S1(net206),
    .X(_0228_));
 sky130_fd_sc_hd__a21oi_1 _3853_ (.A1(net205),
    .A2(_0228_),
    .B1(net199),
    .Y(_0229_));
 sky130_fd_sc_hd__o31ai_2 _3854_ (.A1(_0212_),
    .A2(_0218_),
    .A3(_0223_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a22oi_4 _3855_ (.A1(_0168_),
    .A2(_0195_),
    .B1(_0230_),
    .B2(_0211_),
    .Y(_3279_));
 sky130_fd_sc_hd__inv_6 _3856_ (.A(net11),
    .Y(_0231_));
 sky130_fd_sc_hd__a21oi_4 _3857_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__a21oi_1 _3858_ (.A1(_0119_),
    .A2(_0170_),
    .B1(\dp.rf.rf[24][31] ),
    .Y(_0233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_266 ();
 sky130_fd_sc_hd__mux2i_1 _3862_ (.A0(\dp.rf.rf[26][31] ),
    .A1(\dp.rf.rf[27][31] ),
    .S(net211),
    .Y(_0237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_264 ();
 sky130_fd_sc_hd__a21oi_1 _3865_ (.A1(net8),
    .A2(_0237_),
    .B1(net207),
    .Y(_0240_));
 sky130_fd_sc_hd__o31ai_1 _3866_ (.A1(\dp.rf.rf[25][31] ),
    .A2(net8),
    .A3(net201),
    .B1(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__mux4_1 _3867_ (.A0(\dp.rf.rf[28][31] ),
    .A1(\dp.rf.rf[29][31] ),
    .A2(\dp.rf.rf[30][31] ),
    .A3(\dp.rf.rf[31][31] ),
    .S0(net211),
    .S1(net8),
    .X(_0242_));
 sky130_fd_sc_hd__a21oi_1 _3868_ (.A1(net207),
    .A2(_0242_),
    .B1(net198),
    .Y(_0243_));
 sky130_fd_sc_hd__o21ai_1 _3869_ (.A1(_0233_),
    .A2(_0241_),
    .B1(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__clkinv_16 _3870_ (.A(net211),
    .Y(_0245_));
 sky130_fd_sc_hd__mux2_1 _3871_ (.A0(\dp.rf.rf[17][31] ),
    .A1(\dp.rf.rf[19][31] ),
    .S(net8),
    .X(_0246_));
 sky130_fd_sc_hd__nand2b_4 _3872_ (.A_N(net211),
    .B(net8),
    .Y(_0247_));
 sky130_fd_sc_hd__o221a_1 _3873_ (.A1(_0245_),
    .A2(_0246_),
    .B1(_0247_),
    .B2(\dp.rf.rf[18][31] ),
    .C1(_0148_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _3874_ (.A(net196),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_263 ();
 sky130_fd_sc_hd__nand3_1 _3876_ (.A(_0245_),
    .B(net205),
    .C(_0145_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21oi_1 _3877_ (.A1(_0119_),
    .A2(_0251_),
    .B1(\dp.rf.rf[16][31] ),
    .Y(_0252_));
 sky130_fd_sc_hd__mux4_1 _3878_ (.A0(\dp.rf.rf[20][31] ),
    .A1(\dp.rf.rf[21][31] ),
    .A2(\dp.rf.rf[22][31] ),
    .A3(\dp.rf.rf[23][31] ),
    .S0(net211),
    .S1(net8),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_1 _3879_ (.A(net190),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__o21ai_1 _3880_ (.A1(_0249_),
    .A2(_0252_),
    .B1(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21oi_4 _3881_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0145_),
    .Y(_0256_));
 sky130_fd_sc_hd__mux4_1 _3882_ (.A0(\dp.rf.rf[10][31] ),
    .A1(\dp.rf.rf[11][31] ),
    .A2(\dp.rf.rf[14][31] ),
    .A3(\dp.rf.rf[15][31] ),
    .S0(net211),
    .S1(net207),
    .X(_0257_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_262 ();
 sky130_fd_sc_hd__mux4_1 _3884_ (.A0(\dp.rf.rf[8][31] ),
    .A1(\dp.rf.rf[9][31] ),
    .A2(\dp.rf.rf[12][31] ),
    .A3(\dp.rf.rf[13][31] ),
    .S0(net211),
    .S1(net207),
    .X(_0259_));
 sky130_fd_sc_hd__mux2i_2 _3885_ (.A0(_0257_),
    .A1(_0259_),
    .S(_0224_),
    .Y(_0260_));
 sky130_fd_sc_hd__mux4_1 _3886_ (.A0(\dp.rf.rf[2][31] ),
    .A1(\dp.rf.rf[3][31] ),
    .A2(\dp.rf.rf[6][31] ),
    .A3(\dp.rf.rf[7][31] ),
    .S0(net211),
    .S1(net207),
    .X(_0261_));
 sky130_fd_sc_hd__inv_1 _3887_ (.A(\dp.rf.rf[4][31] ),
    .Y(_0262_));
 sky130_fd_sc_hd__nor2b_4 _3888_ (.A(net211),
    .B_N(net208),
    .Y(_0263_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_260 ();
 sky130_fd_sc_hd__mux2i_1 _3891_ (.A0(\dp.rf.rf[1][31] ),
    .A1(\dp.rf.rf[5][31] ),
    .S(net207),
    .Y(_0266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_258 ();
 sky130_fd_sc_hd__a221oi_1 _3894_ (.A1(_0262_),
    .A2(net203),
    .B1(_0266_),
    .B2(net211),
    .C1(net8),
    .Y(_0269_));
 sky130_fd_sc_hd__a211oi_1 _3895_ (.A1(net8),
    .A2(_0261_),
    .B1(_0269_),
    .C1(net196),
    .Y(_0270_));
 sky130_fd_sc_hd__or3_4 _3896_ (.A(net11),
    .B(_0130_),
    .C(_0208_),
    .X(_0271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_257 ();
 sky130_fd_sc_hd__a211oi_2 _3898_ (.A1(net185),
    .A2(_0260_),
    .B1(_0270_),
    .C1(_0271_),
    .Y(_0273_));
 sky130_fd_sc_hd__a31oi_4 _3899_ (.A1(net187),
    .A2(_0244_),
    .A3(_0255_),
    .B1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_251 ();
 sky130_fd_sc_hd__mux4_1 _3906_ (.A0(\dp.rf.rf[24][31] ),
    .A1(\dp.rf.rf[25][31] ),
    .A2(\dp.rf.rf[26][31] ),
    .A3(\dp.rf.rf[27][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0280_));
 sky130_fd_sc_hd__mux4_1 _3907_ (.A0(\dp.rf.rf[16][31] ),
    .A1(\dp.rf.rf[17][31] ),
    .A2(\dp.rf.rf[18][31] ),
    .A3(\dp.rf.rf[19][31] ),
    .S0(net212),
    .S1(net274),
    .X(_0281_));
 sky130_fd_sc_hd__mux4_1 _3908_ (.A0(\dp.rf.rf[28][31] ),
    .A1(\dp.rf.rf[29][31] ),
    .A2(\dp.rf.rf[30][31] ),
    .A3(\dp.rf.rf[31][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0282_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_250 ();
 sky130_fd_sc_hd__mux4_1 _3910_ (.A0(\dp.rf.rf[20][31] ),
    .A1(\dp.rf.rf[21][31] ),
    .A2(\dp.rf.rf[22][31] ),
    .A3(\dp.rf.rf[23][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0284_));
 sky130_fd_sc_hd__mux4_1 _3911_ (.A0(_0280_),
    .A1(_0281_),
    .A2(_0282_),
    .A3(_0284_),
    .S0(_0103_),
    .S1(net15),
    .X(_0285_));
 sky130_fd_sc_hd__clkinv_16 _3912_ (.A(net15),
    .Y(_0286_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_248 ();
 sky130_fd_sc_hd__nor3_4 _3915_ (.A(net274),
    .B(net212),
    .C(net16),
    .Y(_0289_));
 sky130_fd_sc_hd__a21oi_4 _3916_ (.A1(_0286_),
    .A2(_0289_),
    .B1(net17),
    .Y(_0290_));
 sky130_fd_sc_hd__mux4_1 _3917_ (.A0(\dp.rf.rf[8][31] ),
    .A1(\dp.rf.rf[9][31] ),
    .A2(\dp.rf.rf[10][31] ),
    .A3(\dp.rf.rf[11][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0291_));
 sky130_fd_sc_hd__mux4_1 _3918_ (.A0(\dp.rf.rf[0][31] ),
    .A1(\dp.rf.rf[1][31] ),
    .A2(\dp.rf.rf[2][31] ),
    .A3(\dp.rf.rf[3][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0292_));
 sky130_fd_sc_hd__mux4_1 _3919_ (.A0(\dp.rf.rf[12][31] ),
    .A1(\dp.rf.rf[13][31] ),
    .A2(\dp.rf.rf[14][31] ),
    .A3(\dp.rf.rf[15][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0293_));
 sky130_fd_sc_hd__mux4_1 _3920_ (.A0(\dp.rf.rf[4][31] ),
    .A1(\dp.rf.rf[5][31] ),
    .A2(\dp.rf.rf[6][31] ),
    .A3(\dp.rf.rf[7][31] ),
    .S0(net213),
    .S1(net274),
    .X(_0294_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_246 ();
 sky130_fd_sc_hd__mux4_2 _3923_ (.A0(_0291_),
    .A1(_0292_),
    .A2(_0293_),
    .A3(_0294_),
    .S0(_0103_),
    .S1(net15),
    .X(_0297_));
 sky130_fd_sc_hd__a22oi_4 _3924_ (.A1(net17),
    .A2(_0285_),
    .B1(_0290_),
    .B2(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(net179),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__o21ai_1 _3926_ (.A1(net25),
    .A2(net179),
    .B1(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__xor2_1 _3927_ (.A(_0122_),
    .B(_0300_),
    .X(_3283_));
 sky130_fd_sc_hd__inv_1 _3928_ (.A(_3283_),
    .Y(_3287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_243 ();
 sky130_fd_sc_hd__nand2_4 _3932_ (.A(net25),
    .B(_0119_),
    .Y(_0304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_239 ();
 sky130_fd_sc_hd__nand2_1 _3937_ (.A(net24),
    .B(_0130_),
    .Y(_0309_));
 sky130_fd_sc_hd__nand2_1 _3938_ (.A(_0304_),
    .B(_0309_),
    .Y(_3649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_238 ();
 sky130_fd_sc_hd__nand2_8 _3940_ (.A(_0046_),
    .B(_0289_),
    .Y(_0311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_237 ();
 sky130_fd_sc_hd__mux4_1 _3942_ (.A0(\dp.rf.rf[24][30] ),
    .A1(\dp.rf.rf[25][30] ),
    .A2(\dp.rf.rf[26][30] ),
    .A3(\dp.rf.rf[27][30] ),
    .S0(net212),
    .S1(net274),
    .X(_0313_));
 sky130_fd_sc_hd__mux4_1 _3943_ (.A0(\dp.rf.rf[16][30] ),
    .A1(\dp.rf.rf[17][30] ),
    .A2(\dp.rf.rf[18][30] ),
    .A3(\dp.rf.rf[19][30] ),
    .S0(net212),
    .S1(net274),
    .X(_0314_));
 sky130_fd_sc_hd__mux4_1 _3944_ (.A0(\dp.rf.rf[28][30] ),
    .A1(\dp.rf.rf[29][30] ),
    .A2(\dp.rf.rf[30][30] ),
    .A3(\dp.rf.rf[31][30] ),
    .S0(net212),
    .S1(net274),
    .X(_0315_));
 sky130_fd_sc_hd__mux4_1 _3945_ (.A0(\dp.rf.rf[20][30] ),
    .A1(\dp.rf.rf[21][30] ),
    .A2(\dp.rf.rf[22][30] ),
    .A3(\dp.rf.rf[23][30] ),
    .S0(net212),
    .S1(net274),
    .X(_0316_));
 sky130_fd_sc_hd__mux4_1 _3946_ (.A0(_0313_),
    .A1(_0314_),
    .A2(_0315_),
    .A3(_0316_),
    .S0(_0103_),
    .S1(net15),
    .X(_0317_));
 sky130_fd_sc_hd__mux4_1 _3947_ (.A0(\dp.rf.rf[8][30] ),
    .A1(\dp.rf.rf[9][30] ),
    .A2(\dp.rf.rf[10][30] ),
    .A3(\dp.rf.rf[11][30] ),
    .S0(net213),
    .S1(net274),
    .X(_0318_));
 sky130_fd_sc_hd__mux4_1 _3948_ (.A0(\dp.rf.rf[0][30] ),
    .A1(\dp.rf.rf[1][30] ),
    .A2(\dp.rf.rf[2][30] ),
    .A3(\dp.rf.rf[3][30] ),
    .S0(net213),
    .S1(net274),
    .X(_0319_));
 sky130_fd_sc_hd__mux4_1 _3949_ (.A0(\dp.rf.rf[12][30] ),
    .A1(\dp.rf.rf[13][30] ),
    .A2(\dp.rf.rf[14][30] ),
    .A3(\dp.rf.rf[15][30] ),
    .S0(net213),
    .S1(net274),
    .X(_0320_));
 sky130_fd_sc_hd__mux4_1 _3950_ (.A0(\dp.rf.rf[4][30] ),
    .A1(\dp.rf.rf[5][30] ),
    .A2(\dp.rf.rf[6][30] ),
    .A3(\dp.rf.rf[7][30] ),
    .S0(net213),
    .S1(net274),
    .X(_0321_));
 sky130_fd_sc_hd__mux4_1 _3951_ (.A0(_0318_),
    .A1(_0319_),
    .A2(_0320_),
    .A3(_0321_),
    .S0(_0103_),
    .S1(net15),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(_0317_),
    .A1(_0322_),
    .S(_0086_),
    .X(_0323_));
 sky130_fd_sc_hd__nand2_4 _3953_ (.A(_0311_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_1 _3954_ (.A(_0138_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__a21oi_1 _3955_ (.A1(_0138_),
    .A2(_3649_),
    .B1(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__xor2_1 _3956_ (.A(_0122_),
    .B(_0326_),
    .X(_3292_));
 sky130_fd_sc_hd__inv_1 _3957_ (.A(_3292_),
    .Y(_3296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_234 ();
 sky130_fd_sc_hd__mux4_1 _3961_ (.A0(\dp.rf.rf[10][30] ),
    .A1(\dp.rf.rf[11][30] ),
    .A2(\dp.rf.rf[14][30] ),
    .A3(\dp.rf.rf[15][30] ),
    .S0(net209),
    .S1(net207),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _3962_ (.A(net8),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__mux4_1 _3963_ (.A0(\dp.rf.rf[8][30] ),
    .A1(\dp.rf.rf[9][30] ),
    .A2(\dp.rf.rf[12][30] ),
    .A3(\dp.rf.rf[13][30] ),
    .S0(net209),
    .S1(net207),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(net205),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand3_2 _3965_ (.A(net185),
    .B(_0331_),
    .C(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_233 ();
 sky130_fd_sc_hd__mux2_1 _3967_ (.A0(\dp.rf.rf[6][30] ),
    .A1(\dp.rf.rf[7][30] ),
    .S(net209),
    .X(_0336_));
 sky130_fd_sc_hd__a21oi_4 _3968_ (.A1(_0115_),
    .A2(_0117_),
    .B1(net205),
    .Y(_0337_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_232 ();
 sky130_fd_sc_hd__o21ai_0 _3970_ (.A1(_0148_),
    .A2(_0336_),
    .B1(net182),
    .Y(_0339_));
 sky130_fd_sc_hd__a221oi_1 _3971_ (.A1(\dp.rf.rf[3][30] ),
    .A2(net209),
    .B1(net201),
    .B2(\dp.rf.rf[2][30] ),
    .C1(net190),
    .Y(_0340_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_231 ();
 sky130_fd_sc_hd__inv_1 _3973_ (.A(\dp.rf.rf[4][30] ),
    .Y(_0342_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_230 ();
 sky130_fd_sc_hd__mux2i_1 _3975_ (.A0(\dp.rf.rf[1][30] ),
    .A1(\dp.rf.rf[5][30] ),
    .S(net207),
    .Y(_0344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_229 ();
 sky130_fd_sc_hd__a221oi_1 _3977_ (.A1(_0342_),
    .A2(net203),
    .B1(_0344_),
    .B2(net209),
    .C1(net8),
    .Y(_0346_));
 sky130_fd_sc_hd__nor2_2 _3978_ (.A(net210),
    .B(net208),
    .Y(_0347_));
 sky130_fd_sc_hd__a22oi_4 _3979_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0347_),
    .B2(_0145_),
    .Y(_0348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_228 ();
 sky130_fd_sc_hd__o22ai_1 _3981_ (.A1(net196),
    .A2(_0346_),
    .B1(net181),
    .B2(\dp.rf.rf[0][30] ),
    .Y(_0350_));
 sky130_fd_sc_hd__o21ai_2 _3982_ (.A1(_0339_),
    .A2(_0340_),
    .B1(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_227 ();
 sky130_fd_sc_hd__mux4_1 _3984_ (.A0(\dp.rf.rf[26][30] ),
    .A1(\dp.rf.rf[27][30] ),
    .A2(\dp.rf.rf[30][30] ),
    .A3(\dp.rf.rf[31][30] ),
    .S0(net209),
    .S1(net206),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _3985_ (.A(net8),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__mux4_1 _3986_ (.A0(\dp.rf.rf[24][30] ),
    .A1(\dp.rf.rf[25][30] ),
    .A2(\dp.rf.rf[28][30] ),
    .A3(\dp.rf.rf[29][30] ),
    .S0(net209),
    .S1(net206),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(net205),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__a31oi_2 _3988_ (.A1(net10),
    .A2(_0354_),
    .A3(_0356_),
    .B1(_0166_),
    .Y(_0357_));
 sky130_fd_sc_hd__mux2_1 _3989_ (.A0(\dp.rf.rf[22][30] ),
    .A1(\dp.rf.rf[23][30] ),
    .S(net209),
    .X(_0358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_226 ();
 sky130_fd_sc_hd__o21ai_0 _3991_ (.A1(_0148_),
    .A2(_0358_),
    .B1(net182),
    .Y(_0360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_223 ();
 sky130_fd_sc_hd__a221oi_1 _3995_ (.A1(\dp.rf.rf[19][30] ),
    .A2(net209),
    .B1(net201),
    .B2(\dp.rf.rf[18][30] ),
    .C1(net190),
    .Y(_0364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_222 ();
 sky130_fd_sc_hd__inv_1 _3997_ (.A(\dp.rf.rf[20][30] ),
    .Y(_0366_));
 sky130_fd_sc_hd__mux2i_1 _3998_ (.A0(\dp.rf.rf[17][30] ),
    .A1(\dp.rf.rf[21][30] ),
    .S(net206),
    .Y(_0367_));
 sky130_fd_sc_hd__a221oi_1 _3999_ (.A1(_0366_),
    .A2(net203),
    .B1(_0367_),
    .B2(net209),
    .C1(net8),
    .Y(_0368_));
 sky130_fd_sc_hd__o22ai_1 _4000_ (.A1(\dp.rf.rf[16][30] ),
    .A2(net181),
    .B1(_0368_),
    .B2(net196),
    .Y(_0369_));
 sky130_fd_sc_hd__o21ai_1 _4001_ (.A1(_0360_),
    .A2(_0364_),
    .B1(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a32oi_4 _4002_ (.A1(net194),
    .A2(_0334_),
    .A3(_0351_),
    .B1(_0357_),
    .B2(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_221 ();
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(net22),
    .B(_0130_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _4005_ (.A(_0304_),
    .B(_0372_),
    .Y(_3645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_218 ();
 sky130_fd_sc_hd__mux4_1 _4009_ (.A0(\dp.rf.rf[28][29] ),
    .A1(\dp.rf.rf[29][29] ),
    .A2(\dp.rf.rf[30][29] ),
    .A3(\dp.rf.rf[31][29] ),
    .S0(net213),
    .S1(net274),
    .X(_0376_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_217 ();
 sky130_fd_sc_hd__mux4_1 _4011_ (.A0(\dp.rf.rf[20][29] ),
    .A1(\dp.rf.rf[21][29] ),
    .A2(\dp.rf.rf[22][29] ),
    .A3(\dp.rf.rf[23][29] ),
    .S0(net215),
    .S1(net274),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _4012_ (.A0(\dp.rf.rf[24][29] ),
    .A1(\dp.rf.rf[25][29] ),
    .A2(\dp.rf.rf[26][29] ),
    .A3(\dp.rf.rf[27][29] ),
    .S0(net213),
    .S1(net274),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _4013_ (.A0(\dp.rf.rf[16][29] ),
    .A1(\dp.rf.rf[17][29] ),
    .A2(\dp.rf.rf[18][29] ),
    .A3(\dp.rf.rf[19][29] ),
    .S0(net215),
    .S1(net274),
    .X(_0380_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_216 ();
 sky130_fd_sc_hd__mux4_1 _4015_ (.A0(_0376_),
    .A1(_0378_),
    .A2(_0379_),
    .A3(_0380_),
    .S0(_0103_),
    .S1(_0286_),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _4016_ (.A(_0086_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_212 ();
 sky130_fd_sc_hd__mux4_1 _4021_ (.A0(\dp.rf.rf[12][29] ),
    .A1(\dp.rf.rf[13][29] ),
    .A2(\dp.rf.rf[14][29] ),
    .A3(\dp.rf.rf[15][29] ),
    .S0(net215),
    .S1(net14),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_1 _4022_ (.A(_0286_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_211 ();
 sky130_fd_sc_hd__mux4_1 _4024_ (.A0(\dp.rf.rf[8][29] ),
    .A1(\dp.rf.rf[9][29] ),
    .A2(\dp.rf.rf[10][29] ),
    .A3(\dp.rf.rf[11][29] ),
    .S0(net215),
    .S1(net14),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_1 _4025_ (.A(net15),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _4026_ (.A(_0389_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_2 _4027_ (.A(net17),
    .B(net16),
    .Y(_0394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_209 ();
 sky130_fd_sc_hd__mux4_1 _4030_ (.A0(\dp.rf.rf[4][29] ),
    .A1(\dp.rf.rf[5][29] ),
    .A2(\dp.rf.rf[6][29] ),
    .A3(\dp.rf.rf[7][29] ),
    .S0(net215),
    .S1(net14),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _4031_ (.A(net15),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__mux4_1 _4032_ (.A0(\dp.rf.rf[0][29] ),
    .A1(\dp.rf.rf[1][29] ),
    .A2(\dp.rf.rf[2][29] ),
    .A3(\dp.rf.rf[3][29] ),
    .S0(net215),
    .S1(net14),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _4033_ (.A(_0286_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__and2_4 _4034_ (.A(_0046_),
    .B(_0289_),
    .X(_0401_));
 sky130_fd_sc_hd__a31oi_1 _4035_ (.A1(_0394_),
    .A2(_0398_),
    .A3(_0400_),
    .B1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__o31ai_2 _4036_ (.A1(net17),
    .A2(_0103_),
    .A3(_0393_),
    .B1(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nor2_4 _4037_ (.A(_0383_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__mux2i_1 _4038_ (.A0(_3645_),
    .A1(_0404_),
    .S(net179),
    .Y(_0405_));
 sky130_fd_sc_hd__xor2_1 _4039_ (.A(_0122_),
    .B(_0405_),
    .X(_3300_));
 sky130_fd_sc_hd__inv_1 _4040_ (.A(_3300_),
    .Y(_3304_));
 sky130_fd_sc_hd__a211oi_4 _4041_ (.A1(_0115_),
    .A2(_0117_),
    .B1(net205),
    .C1(_0231_),
    .Y(_0406_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_206 ();
 sky130_fd_sc_hd__mux2i_1 _4045_ (.A0(\dp.rf.rf[30][29] ),
    .A1(\dp.rf.rf[31][29] ),
    .S(net211),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(net207),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a221o_1 _4047_ (.A1(\dp.rf.rf[27][29] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[26][29] ),
    .C1(net190),
    .X(_0412_));
 sky130_fd_sc_hd__mux2i_1 _4048_ (.A0(\dp.rf.rf[24][29] ),
    .A1(\dp.rf.rf[28][29] ),
    .S(net207),
    .Y(_0413_));
 sky130_fd_sc_hd__mux2i_1 _4049_ (.A0(\dp.rf.rf[25][29] ),
    .A1(\dp.rf.rf[29][29] ),
    .S(net207),
    .Y(_0414_));
 sky130_fd_sc_hd__nand2b_4 _4050_ (.A_N(net8),
    .B(net209),
    .Y(_0415_));
 sky130_fd_sc_hd__o221ai_1 _4051_ (.A1(_0170_),
    .A2(_0413_),
    .B1(_0414_),
    .B2(_0415_),
    .C1(net10),
    .Y(_0416_));
 sky130_fd_sc_hd__a32o_1 _4052_ (.A1(_0406_),
    .A2(_0411_),
    .A3(_0412_),
    .B1(_0416_),
    .B2(net188),
    .X(_0417_));
 sky130_fd_sc_hd__nor2b_1 _4053_ (.A(net211),
    .B_N(\dp.rf.rf[22][29] ),
    .Y(_0418_));
 sky130_fd_sc_hd__a211oi_1 _4054_ (.A1(\dp.rf.rf[23][29] ),
    .A2(net211),
    .B1(_0148_),
    .C1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_205 ();
 sky130_fd_sc_hd__a221oi_1 _4056_ (.A1(\dp.rf.rf[19][29] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[18][29] ),
    .C1(net190),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_1 _4057_ (.A(\dp.rf.rf[20][29] ),
    .Y(_0422_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_204 ();
 sky130_fd_sc_hd__mux2i_1 _4059_ (.A0(\dp.rf.rf[17][29] ),
    .A1(\dp.rf.rf[21][29] ),
    .S(net207),
    .Y(_0424_));
 sky130_fd_sc_hd__a221oi_1 _4060_ (.A1(_0422_),
    .A2(net203),
    .B1(_0424_),
    .B2(net211),
    .C1(net8),
    .Y(_0425_));
 sky130_fd_sc_hd__o22ai_1 _4061_ (.A1(\dp.rf.rf[16][29] ),
    .A2(net180),
    .B1(_0425_),
    .B2(net195),
    .Y(_0426_));
 sky130_fd_sc_hd__o31ai_2 _4062_ (.A1(net192),
    .A2(_0419_),
    .A3(_0421_),
    .B1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__mux4_1 _4063_ (.A0(\dp.rf.rf[2][29] ),
    .A1(\dp.rf.rf[3][29] ),
    .A2(\dp.rf.rf[6][29] ),
    .A3(\dp.rf.rf[7][29] ),
    .S0(net211),
    .S1(net207),
    .X(_0428_));
 sky130_fd_sc_hd__inv_1 _4064_ (.A(\dp.rf.rf[4][29] ),
    .Y(_0429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_203 ();
 sky130_fd_sc_hd__mux2i_1 _4066_ (.A0(\dp.rf.rf[1][29] ),
    .A1(\dp.rf.rf[5][29] ),
    .S(net207),
    .Y(_0431_));
 sky130_fd_sc_hd__a221oi_1 _4067_ (.A1(_0429_),
    .A2(net204),
    .B1(_0431_),
    .B2(net211),
    .C1(net8),
    .Y(_0432_));
 sky130_fd_sc_hd__a211oi_1 _4068_ (.A1(net8),
    .A2(_0428_),
    .B1(_0432_),
    .C1(net195),
    .Y(_0433_));
 sky130_fd_sc_hd__mux4_1 _4069_ (.A0(\dp.rf.rf[10][29] ),
    .A1(\dp.rf.rf[11][29] ),
    .A2(\dp.rf.rf[14][29] ),
    .A3(\dp.rf.rf[15][29] ),
    .S0(net211),
    .S1(net207),
    .X(_0434_));
 sky130_fd_sc_hd__mux4_1 _4070_ (.A0(\dp.rf.rf[8][29] ),
    .A1(\dp.rf.rf[9][29] ),
    .A2(\dp.rf.rf[12][29] ),
    .A3(\dp.rf.rf[13][29] ),
    .S0(net211),
    .S1(net207),
    .X(_0435_));
 sky130_fd_sc_hd__and2_0 _4071_ (.A(_0224_),
    .B(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a211oi_1 _4072_ (.A1(net182),
    .A2(_0434_),
    .B1(_0436_),
    .C1(net198),
    .Y(_0437_));
 sky130_fd_sc_hd__nor3_2 _4073_ (.A(_0271_),
    .B(_0433_),
    .C(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__a21oi_4 _4074_ (.A1(_0417_),
    .A2(_0427_),
    .B1(_0438_),
    .Y(_3303_));
 sky130_fd_sc_hd__nand2_1 _4075_ (.A(net21),
    .B(_0130_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _4076_ (.A(_0304_),
    .B(_0439_),
    .Y(_3641_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_201 ();
 sky130_fd_sc_hd__mux4_1 _4079_ (.A0(\dp.rf.rf[4][28] ),
    .A1(\dp.rf.rf[5][28] ),
    .A2(\dp.rf.rf[6][28] ),
    .A3(\dp.rf.rf[7][28] ),
    .S0(net215),
    .S1(net14),
    .X(_0442_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_200 ();
 sky130_fd_sc_hd__mux4_1 _4081_ (.A0(\dp.rf.rf[0][28] ),
    .A1(\dp.rf.rf[1][28] ),
    .A2(\dp.rf.rf[2][28] ),
    .A3(\dp.rf.rf[3][28] ),
    .S0(net215),
    .S1(net14),
    .X(_0444_));
 sky130_fd_sc_hd__mux2i_4 _4082_ (.A0(_0442_),
    .A1(_0444_),
    .S(_0286_),
    .Y(_0445_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_199 ();
 sky130_fd_sc_hd__mux4_1 _4084_ (.A0(\dp.rf.rf[8][28] ),
    .A1(\dp.rf.rf[9][28] ),
    .A2(\dp.rf.rf[10][28] ),
    .A3(\dp.rf.rf[11][28] ),
    .S0(net215),
    .S1(net274),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _4085_ (.A(net16),
    .B(_0046_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand3_1 _4086_ (.A(_0086_),
    .B(net15),
    .C(net16),
    .Y(_0449_));
 sky130_fd_sc_hd__mux4_1 _4087_ (.A0(\dp.rf.rf[12][28] ),
    .A1(\dp.rf.rf[13][28] ),
    .A2(\dp.rf.rf[14][28] ),
    .A3(\dp.rf.rf[15][28] ),
    .S0(net215),
    .S1(net14),
    .X(_0450_));
 sky130_fd_sc_hd__o221ai_2 _4088_ (.A1(_0447_),
    .A2(_0448_),
    .B1(_0449_),
    .B2(_0450_),
    .C1(_0311_),
    .Y(_0451_));
 sky130_fd_sc_hd__mux4_1 _4089_ (.A0(\dp.rf.rf[28][28] ),
    .A1(\dp.rf.rf[29][28] ),
    .A2(\dp.rf.rf[30][28] ),
    .A3(\dp.rf.rf[31][28] ),
    .S0(net213),
    .S1(net277),
    .X(_0452_));
 sky130_fd_sc_hd__mux4_1 _4090_ (.A0(\dp.rf.rf[20][28] ),
    .A1(\dp.rf.rf[21][28] ),
    .A2(\dp.rf.rf[22][28] ),
    .A3(\dp.rf.rf[23][28] ),
    .S0(net213),
    .S1(net277),
    .X(_0453_));
 sky130_fd_sc_hd__mux4_1 _4091_ (.A0(\dp.rf.rf[24][28] ),
    .A1(\dp.rf.rf[25][28] ),
    .A2(\dp.rf.rf[26][28] ),
    .A3(\dp.rf.rf[27][28] ),
    .S0(net213),
    .S1(net277),
    .X(_0454_));
 sky130_fd_sc_hd__mux4_1 _4092_ (.A0(\dp.rf.rf[16][28] ),
    .A1(\dp.rf.rf[17][28] ),
    .A2(\dp.rf.rf[18][28] ),
    .A3(\dp.rf.rf[19][28] ),
    .S0(net213),
    .S1(net277),
    .X(_0455_));
 sky130_fd_sc_hd__mux4_2 _4093_ (.A0(_0452_),
    .A1(_0453_),
    .A2(_0454_),
    .A3(_0455_),
    .S0(_0103_),
    .S1(_0286_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_1 _4094_ (.A(_0086_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__a211o_4 _4095_ (.A1(_0394_),
    .A2(_0445_),
    .B1(_0451_),
    .C1(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_1 _4096_ (.A(_0138_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _4097_ (.A1(_0138_),
    .A2(_3641_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__xor2_1 _4098_ (.A(_0122_),
    .B(_0460_),
    .X(_3308_));
 sky130_fd_sc_hd__inv_1 _4099_ (.A(_3308_),
    .Y(_3312_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_198 ();
 sky130_fd_sc_hd__mux4_1 _4101_ (.A0(\dp.rf.rf[18][28] ),
    .A1(\dp.rf.rf[19][28] ),
    .A2(\dp.rf.rf[22][28] ),
    .A3(\dp.rf.rf[23][28] ),
    .S0(net209),
    .S1(net206),
    .X(_0462_));
 sky130_fd_sc_hd__nand2_1 _4102_ (.A(_0406_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__mux2i_1 _4103_ (.A0(\dp.rf.rf[17][28] ),
    .A1(\dp.rf.rf[21][28] ),
    .S(net206),
    .Y(_0464_));
 sky130_fd_sc_hd__nor3b_1 _4104_ (.A(\dp.rf.rf[20][28] ),
    .B(net209),
    .C_N(net206),
    .Y(_0465_));
 sky130_fd_sc_hd__nor3_1 _4105_ (.A(\dp.rf.rf[16][28] ),
    .B(net209),
    .C(net206),
    .Y(_0466_));
 sky130_fd_sc_hd__a2111oi_0 _4106_ (.A1(net209),
    .A2(_0464_),
    .B1(_0465_),
    .C1(_0466_),
    .D1(net8),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_1 _4107_ (.A1(net10),
    .A2(_0467_),
    .B1(net187),
    .Y(_0468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_197 ();
 sky130_fd_sc_hd__nand4_1 _4109_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[26][28] ),
    .Y(_0470_));
 sky130_fd_sc_hd__o2bb2ai_1 _4110_ (.A1_N(\dp.rf.rf[26][28] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_196 ();
 sky130_fd_sc_hd__and2_0 _4112_ (.A(\dp.rf.rf[27][28] ),
    .B(net209),
    .X(_0473_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_195 ();
 sky130_fd_sc_hd__mux2i_1 _4114_ (.A0(\dp.rf.rf[30][28] ),
    .A1(\dp.rf.rf[31][28] ),
    .S(net209),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _4115_ (.A(net206),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_194 ();
 sky130_fd_sc_hd__o311ai_4 _4117_ (.A1(net190),
    .A2(_0471_),
    .A3(_0473_),
    .B1(_0476_),
    .C1(net182),
    .Y(_0478_));
 sky130_fd_sc_hd__mux4_1 _4118_ (.A0(\dp.rf.rf[24][28] ),
    .A1(\dp.rf.rf[25][28] ),
    .A2(\dp.rf.rf[28][28] ),
    .A3(\dp.rf.rf[29][28] ),
    .S0(net209),
    .S1(net206),
    .X(_0479_));
 sky130_fd_sc_hd__a21oi_1 _4119_ (.A1(net205),
    .A2(_0479_),
    .B1(net198),
    .Y(_0480_));
 sky130_fd_sc_hd__a22oi_4 _4120_ (.A1(_0463_),
    .A2(_0468_),
    .B1(_0478_),
    .B2(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_193 ();
 sky130_fd_sc_hd__mux4_1 _4122_ (.A0(\dp.rf.rf[10][28] ),
    .A1(\dp.rf.rf[11][28] ),
    .A2(\dp.rf.rf[14][28] ),
    .A3(\dp.rf.rf[15][28] ),
    .S0(net211),
    .S1(net207),
    .X(_0483_));
 sky130_fd_sc_hd__mux4_1 _4123_ (.A0(\dp.rf.rf[8][28] ),
    .A1(\dp.rf.rf[9][28] ),
    .A2(\dp.rf.rf[12][28] ),
    .A3(\dp.rf.rf[13][28] ),
    .S0(net211),
    .S1(net207),
    .X(_0484_));
 sky130_fd_sc_hd__mux2i_2 _4124_ (.A0(_0483_),
    .A1(_0484_),
    .S(_0224_),
    .Y(_0485_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_192 ();
 sky130_fd_sc_hd__mux4_1 _4126_ (.A0(\dp.rf.rf[2][28] ),
    .A1(\dp.rf.rf[3][28] ),
    .A2(\dp.rf.rf[6][28] ),
    .A3(\dp.rf.rf[7][28] ),
    .S0(net211),
    .S1(net207),
    .X(_0487_));
 sky130_fd_sc_hd__inv_1 _4127_ (.A(\dp.rf.rf[4][28] ),
    .Y(_0488_));
 sky130_fd_sc_hd__mux2i_1 _4128_ (.A0(\dp.rf.rf[1][28] ),
    .A1(\dp.rf.rf[5][28] ),
    .S(net207),
    .Y(_0489_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_191 ();
 sky130_fd_sc_hd__a221oi_1 _4130_ (.A1(_0488_),
    .A2(net204),
    .B1(_0489_),
    .B2(net211),
    .C1(net8),
    .Y(_0491_));
 sky130_fd_sc_hd__a21oi_2 _4131_ (.A1(net8),
    .A2(_0487_),
    .B1(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__a21oi_4 _4132_ (.A1(_0115_),
    .A2(_0117_),
    .B1(net10),
    .Y(_0493_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_190 ();
 sky130_fd_sc_hd__a221oi_4 _4134_ (.A1(net185),
    .A2(_0485_),
    .B1(_0492_),
    .B2(_0493_),
    .C1(_0271_),
    .Y(_0495_));
 sky130_fd_sc_hd__nor2_4 _4135_ (.A(_0481_),
    .B(_0495_),
    .Y(_3311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_187 ();
 sky130_fd_sc_hd__mux4_1 _4139_ (.A0(\dp.rf.rf[24][27] ),
    .A1(\dp.rf.rf[25][27] ),
    .A2(\dp.rf.rf[26][27] ),
    .A3(\dp.rf.rf[27][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0499_));
 sky130_fd_sc_hd__mux4_1 _4140_ (.A0(\dp.rf.rf[16][27] ),
    .A1(\dp.rf.rf[17][27] ),
    .A2(\dp.rf.rf[18][27] ),
    .A3(\dp.rf.rf[19][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0500_));
 sky130_fd_sc_hd__mux4_1 _4141_ (.A0(\dp.rf.rf[28][27] ),
    .A1(\dp.rf.rf[29][27] ),
    .A2(\dp.rf.rf[30][27] ),
    .A3(\dp.rf.rf[31][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_186 ();
 sky130_fd_sc_hd__mux4_1 _4143_ (.A0(\dp.rf.rf[20][27] ),
    .A1(\dp.rf.rf[21][27] ),
    .A2(\dp.rf.rf[22][27] ),
    .A3(\dp.rf.rf[23][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_184 ();
 sky130_fd_sc_hd__mux4_1 _4146_ (.A0(_0499_),
    .A1(_0500_),
    .A2(_0501_),
    .A3(_0503_),
    .S0(_0103_),
    .S1(net15),
    .X(_0506_));
 sky130_fd_sc_hd__mux4_1 _4147_ (.A0(\dp.rf.rf[8][27] ),
    .A1(\dp.rf.rf[9][27] ),
    .A2(\dp.rf.rf[10][27] ),
    .A3(\dp.rf.rf[11][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0507_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_183 ();
 sky130_fd_sc_hd__mux4_1 _4149_ (.A0(\dp.rf.rf[0][27] ),
    .A1(\dp.rf.rf[1][27] ),
    .A2(\dp.rf.rf[2][27] ),
    .A3(\dp.rf.rf[3][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0509_));
 sky130_fd_sc_hd__mux4_1 _4150_ (.A0(\dp.rf.rf[12][27] ),
    .A1(\dp.rf.rf[13][27] ),
    .A2(\dp.rf.rf[14][27] ),
    .A3(\dp.rf.rf[15][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0510_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_181 ();
 sky130_fd_sc_hd__mux4_1 _4153_ (.A0(\dp.rf.rf[4][27] ),
    .A1(\dp.rf.rf[5][27] ),
    .A2(\dp.rf.rf[6][27] ),
    .A3(\dp.rf.rf[7][27] ),
    .S0(net213),
    .S1(net14),
    .X(_0513_));
 sky130_fd_sc_hd__mux4_2 _4154_ (.A0(_0507_),
    .A1(_0509_),
    .A2(_0510_),
    .A3(_0513_),
    .S0(_0103_),
    .S1(net15),
    .X(_0514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_180 ();
 sky130_fd_sc_hd__a22oi_4 _4156_ (.A1(net17),
    .A2(_0506_),
    .B1(_0514_),
    .B2(_0290_),
    .Y(_0516_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_179 ();
 sky130_fd_sc_hd__nand2_1 _4158_ (.A(net20),
    .B(_0130_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _4159_ (.A(_0304_),
    .B(_0518_),
    .Y(_3637_));
 sky130_fd_sc_hd__nor2_1 _4160_ (.A(net179),
    .B(_3637_),
    .Y(_0519_));
 sky130_fd_sc_hd__a21oi_1 _4161_ (.A1(net179),
    .A2(_0516_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__xnor2_1 _4162_ (.A(_0122_),
    .B(_0520_),
    .Y(_3316_));
 sky130_fd_sc_hd__inv_1 _4163_ (.A(_3316_),
    .Y(_3320_));
 sky130_fd_sc_hd__mux4_1 _4164_ (.A0(\dp.rf.rf[10][27] ),
    .A1(\dp.rf.rf[11][27] ),
    .A2(\dp.rf.rf[14][27] ),
    .A3(\dp.rf.rf[15][27] ),
    .S0(net211),
    .S1(net207),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_1 _4165_ (.A(net8),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__mux4_1 _4166_ (.A0(\dp.rf.rf[8][27] ),
    .A1(\dp.rf.rf[9][27] ),
    .A2(\dp.rf.rf[12][27] ),
    .A3(\dp.rf.rf[13][27] ),
    .S0(net211),
    .S1(net207),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(_0224_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__and3_1 _4168_ (.A(net185),
    .B(_0522_),
    .C(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__mux4_1 _4169_ (.A0(\dp.rf.rf[2][27] ),
    .A1(\dp.rf.rf[3][27] ),
    .A2(\dp.rf.rf[6][27] ),
    .A3(\dp.rf.rf[7][27] ),
    .S0(net211),
    .S1(net207),
    .X(_0526_));
 sky130_fd_sc_hd__mux2i_1 _4170_ (.A0(\dp.rf.rf[1][27] ),
    .A1(\dp.rf.rf[5][27] ),
    .S(net207),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2b_4 _4171_ (.A_N(net211),
    .B(net207),
    .Y(_0528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_178 ();
 sky130_fd_sc_hd__nor2_1 _4173_ (.A(\dp.rf.rf[4][27] ),
    .B(_0528_),
    .Y(_0530_));
 sky130_fd_sc_hd__a211oi_1 _4174_ (.A1(net211),
    .A2(_0527_),
    .B1(_0530_),
    .C1(net8),
    .Y(_0531_));
 sky130_fd_sc_hd__a211oi_2 _4175_ (.A1(net8),
    .A2(_0526_),
    .B1(_0531_),
    .C1(net196),
    .Y(_0532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_177 ();
 sky130_fd_sc_hd__mux2i_1 _4177_ (.A0(\dp.rf.rf[30][27] ),
    .A1(\dp.rf.rf[31][27] ),
    .S(net211),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _4178_ (.A(net207),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_176 ();
 sky130_fd_sc_hd__a221o_1 _4180_ (.A1(\dp.rf.rf[27][27] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[26][27] ),
    .C1(net190),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_1 _4181_ (.A0(\dp.rf.rf[24][27] ),
    .A1(\dp.rf.rf[25][27] ),
    .A2(\dp.rf.rf[28][27] ),
    .A3(\dp.rf.rf[29][27] ),
    .S0(net211),
    .S1(net207),
    .X(_0538_));
 sky130_fd_sc_hd__nand2_1 _4182_ (.A(_0224_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _4183_ (.A(net185),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_175 ();
 sky130_fd_sc_hd__a32oi_2 _4185_ (.A1(_0406_),
    .A2(_0535_),
    .A3(_0537_),
    .B1(_0540_),
    .B2(net187),
    .Y(_0542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__mux2i_1 _4188_ (.A0(\dp.rf.rf[22][27] ),
    .A1(\dp.rf.rf[23][27] ),
    .S(net211),
    .Y(_0545_));
 sky130_fd_sc_hd__a21oi_1 _4189_ (.A1(net207),
    .A2(_0545_),
    .B1(net192),
    .Y(_0546_));
 sky130_fd_sc_hd__a221o_1 _4190_ (.A1(\dp.rf.rf[19][27] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[18][27] ),
    .C1(net190),
    .X(_0547_));
 sky130_fd_sc_hd__inv_1 _4191_ (.A(\dp.rf.rf[20][27] ),
    .Y(_0548_));
 sky130_fd_sc_hd__mux2i_1 _4192_ (.A0(\dp.rf.rf[17][27] ),
    .A1(\dp.rf.rf[21][27] ),
    .S(net207),
    .Y(_0549_));
 sky130_fd_sc_hd__a221oi_1 _4193_ (.A1(_0548_),
    .A2(net203),
    .B1(_0549_),
    .B2(net211),
    .C1(net8),
    .Y(_0550_));
 sky130_fd_sc_hd__o22a_1 _4194_ (.A1(\dp.rf.rf[16][27] ),
    .A2(net180),
    .B1(_0550_),
    .B2(net196),
    .X(_0551_));
 sky130_fd_sc_hd__a21oi_1 _4195_ (.A1(_0546_),
    .A2(_0547_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__o32ai_4 _4196_ (.A1(_0271_),
    .A2(_0525_),
    .A3(_0532_),
    .B1(_0542_),
    .B2(_0552_),
    .Y(_3315_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(_3315_),
    .Y(_3319_));
 sky130_fd_sc_hd__nand2_1 _4198_ (.A(net19),
    .B(_0130_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _4199_ (.A(_0304_),
    .B(_0553_),
    .Y(_3633_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_170 ();
 sky130_fd_sc_hd__mux4_1 _4203_ (.A0(\dp.rf.rf[24][26] ),
    .A1(\dp.rf.rf[25][26] ),
    .A2(\dp.rf.rf[26][26] ),
    .A3(\dp.rf.rf[27][26] ),
    .S0(net213),
    .S1(net278),
    .X(_0557_));
 sky130_fd_sc_hd__mux4_1 _4204_ (.A0(\dp.rf.rf[16][26] ),
    .A1(\dp.rf.rf[17][26] ),
    .A2(\dp.rf.rf[18][26] ),
    .A3(\dp.rf.rf[19][26] ),
    .S0(net213),
    .S1(net278),
    .X(_0558_));
 sky130_fd_sc_hd__mux4_1 _4205_ (.A0(\dp.rf.rf[28][26] ),
    .A1(\dp.rf.rf[29][26] ),
    .A2(\dp.rf.rf[30][26] ),
    .A3(\dp.rf.rf[31][26] ),
    .S0(net213),
    .S1(net278),
    .X(_0559_));
 sky130_fd_sc_hd__mux4_1 _4206_ (.A0(\dp.rf.rf[20][26] ),
    .A1(\dp.rf.rf[21][26] ),
    .A2(\dp.rf.rf[22][26] ),
    .A3(\dp.rf.rf[23][26] ),
    .S0(net213),
    .S1(net278),
    .X(_0560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__mux4_1 _4208_ (.A0(_0557_),
    .A1(_0558_),
    .A2(_0559_),
    .A3(_0560_),
    .S0(_0103_),
    .S1(net15),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_1 _4209_ (.A(net17),
    .B(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__mux4_1 _4210_ (.A0(\dp.rf.rf[8][26] ),
    .A1(\dp.rf.rf[9][26] ),
    .A2(\dp.rf.rf[10][26] ),
    .A3(\dp.rf.rf[11][26] ),
    .S0(net215),
    .S1(net14),
    .X(_0564_));
 sky130_fd_sc_hd__mux4_1 _4211_ (.A0(\dp.rf.rf[0][26] ),
    .A1(\dp.rf.rf[1][26] ),
    .A2(\dp.rf.rf[2][26] ),
    .A3(\dp.rf.rf[3][26] ),
    .S0(net215),
    .S1(net14),
    .X(_0565_));
 sky130_fd_sc_hd__mux4_1 _4212_ (.A0(\dp.rf.rf[12][26] ),
    .A1(\dp.rf.rf[13][26] ),
    .A2(\dp.rf.rf[14][26] ),
    .A3(\dp.rf.rf[15][26] ),
    .S0(net215),
    .S1(net14),
    .X(_0566_));
 sky130_fd_sc_hd__mux4_1 _4213_ (.A0(\dp.rf.rf[4][26] ),
    .A1(\dp.rf.rf[5][26] ),
    .A2(\dp.rf.rf[6][26] ),
    .A3(\dp.rf.rf[7][26] ),
    .S0(net215),
    .S1(net14),
    .X(_0567_));
 sky130_fd_sc_hd__mux4_1 _4214_ (.A0(_0564_),
    .A1(_0565_),
    .A2(_0566_),
    .A3(_0567_),
    .S0(_0103_),
    .S1(net15),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _4215_ (.A(_0086_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(_0563_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_4 _4217_ (.A(_0311_),
    .B(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor2_1 _4218_ (.A(_0138_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__a21oi_1 _4219_ (.A1(_0138_),
    .A2(_3633_),
    .B1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__xor2_1 _4220_ (.A(_0122_),
    .B(_0573_),
    .X(_3324_));
 sky130_fd_sc_hd__inv_1 _4221_ (.A(_3324_),
    .Y(_3328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(\dp.rf.rf[26][26] ),
    .A1(\dp.rf.rf[27][26] ),
    .S(net7),
    .X(_0576_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__mux2i_1 _4226_ (.A0(\dp.rf.rf[30][26] ),
    .A1(\dp.rf.rf[31][26] ),
    .S(net7),
    .Y(_0578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__a21oi_1 _4229_ (.A1(net206),
    .A2(_0578_),
    .B1(_0224_),
    .Y(_0581_));
 sky130_fd_sc_hd__o21ai_0 _4230_ (.A1(net189),
    .A2(_0576_),
    .B1(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__mux4_1 _4231_ (.A0(\dp.rf.rf[24][26] ),
    .A1(\dp.rf.rf[25][26] ),
    .A2(\dp.rf.rf[28][26] ),
    .A3(\dp.rf.rf[29][26] ),
    .S0(net7),
    .S1(net206),
    .X(_0583_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_163 ();
 sky130_fd_sc_hd__a21oi_1 _4233_ (.A1(_0224_),
    .A2(_0583_),
    .B1(net198),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _4234_ (.A(_0582_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__nor2b_1 _4238_ (.A(net7),
    .B_N(\dp.rf.rf[22][26] ),
    .Y(_0590_));
 sky130_fd_sc_hd__a211oi_1 _4239_ (.A1(\dp.rf.rf[23][26] ),
    .A2(net7),
    .B1(_0148_),
    .C1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__a221oi_1 _4241_ (.A1(\dp.rf.rf[19][26] ),
    .A2(net7),
    .B1(net201),
    .B2(\dp.rf.rf[18][26] ),
    .C1(net189),
    .Y(_0593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__inv_1 _4243_ (.A(\dp.rf.rf[20][26] ),
    .Y(_0595_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__mux2i_1 _4246_ (.A0(\dp.rf.rf[17][26] ),
    .A1(\dp.rf.rf[21][26] ),
    .S(net206),
    .Y(_0598_));
 sky130_fd_sc_hd__a221oi_1 _4247_ (.A1(_0595_),
    .A2(net204),
    .B1(_0598_),
    .B2(net7),
    .C1(net8),
    .Y(_0599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__o22ai_1 _4249_ (.A1(\dp.rf.rf[16][26] ),
    .A2(net180),
    .B1(_0599_),
    .B2(net195),
    .Y(_0601_));
 sky130_fd_sc_hd__o31ai_2 _4250_ (.A1(net192),
    .A2(_0591_),
    .A3(_0593_),
    .B1(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__mux4_1 _4252_ (.A0(\dp.rf.rf[2][26] ),
    .A1(\dp.rf.rf[3][26] ),
    .A2(\dp.rf.rf[6][26] ),
    .A3(\dp.rf.rf[7][26] ),
    .S0(net211),
    .S1(net207),
    .X(_0604_));
 sky130_fd_sc_hd__inv_1 _4253_ (.A(\dp.rf.rf[4][26] ),
    .Y(_0605_));
 sky130_fd_sc_hd__mux2i_1 _4254_ (.A0(\dp.rf.rf[1][26] ),
    .A1(\dp.rf.rf[5][26] ),
    .S(net207),
    .Y(_0606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__a221oi_1 _4256_ (.A1(_0605_),
    .A2(net204),
    .B1(_0606_),
    .B2(net211),
    .C1(net8),
    .Y(_0608_));
 sky130_fd_sc_hd__a21oi_1 _4257_ (.A1(net8),
    .A2(_0604_),
    .B1(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__a21oi_1 _4258_ (.A1(_0493_),
    .A2(_0609_),
    .B1(_0271_),
    .Y(_0610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__nor2b_1 _4261_ (.A(net211),
    .B_N(\dp.rf.rf[14][26] ),
    .Y(_0613_));
 sky130_fd_sc_hd__a211oi_1 _4262_ (.A1(\dp.rf.rf[15][26] ),
    .A2(net211),
    .B1(_0148_),
    .C1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__a221oi_1 _4263_ (.A1(\dp.rf.rf[11][26] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[10][26] ),
    .C1(net189),
    .Y(_0615_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__mux4_1 _4266_ (.A0(\dp.rf.rf[8][26] ),
    .A1(\dp.rf.rf[9][26] ),
    .A2(\dp.rf.rf[12][26] ),
    .A3(\dp.rf.rf[13][26] ),
    .S0(net211),
    .S1(net207),
    .X(_0618_));
 sky130_fd_sc_hd__a21oi_1 _4267_ (.A1(_0224_),
    .A2(_0618_),
    .B1(net198),
    .Y(_0619_));
 sky130_fd_sc_hd__o31ai_2 _4268_ (.A1(net192),
    .A2(_0614_),
    .A3(_0615_),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__a32oi_4 _4269_ (.A1(net188),
    .A2(_0586_),
    .A3(_0602_),
    .B1(_0610_),
    .B2(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_148 ();
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(net18),
    .B(_0130_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _4272_ (.A(_0304_),
    .B(_0622_),
    .Y(_3629_));
 sky130_fd_sc_hd__mux4_1 _4273_ (.A0(\dp.rf.rf[24][25] ),
    .A1(\dp.rf.rf[25][25] ),
    .A2(\dp.rf.rf[26][25] ),
    .A3(\dp.rf.rf[27][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0623_));
 sky130_fd_sc_hd__mux4_1 _4274_ (.A0(\dp.rf.rf[16][25] ),
    .A1(\dp.rf.rf[17][25] ),
    .A2(\dp.rf.rf[18][25] ),
    .A3(\dp.rf.rf[19][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_1 _4275_ (.A0(\dp.rf.rf[28][25] ),
    .A1(\dp.rf.rf[29][25] ),
    .A2(\dp.rf.rf[30][25] ),
    .A3(\dp.rf.rf[31][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_1 _4276_ (.A0(\dp.rf.rf[20][25] ),
    .A1(\dp.rf.rf[21][25] ),
    .A2(\dp.rf.rf[22][25] ),
    .A3(\dp.rf.rf[23][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0626_));
 sky130_fd_sc_hd__mux4_1 _4277_ (.A0(_0623_),
    .A1(_0624_),
    .A2(_0625_),
    .A3(_0626_),
    .S0(_0103_),
    .S1(net15),
    .X(_0627_));
 sky130_fd_sc_hd__nand2_1 _4278_ (.A(net17),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__mux4_1 _4279_ (.A0(\dp.rf.rf[8][25] ),
    .A1(\dp.rf.rf[9][25] ),
    .A2(\dp.rf.rf[10][25] ),
    .A3(\dp.rf.rf[11][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0629_));
 sky130_fd_sc_hd__mux4_1 _4280_ (.A0(\dp.rf.rf[0][25] ),
    .A1(\dp.rf.rf[1][25] ),
    .A2(\dp.rf.rf[2][25] ),
    .A3(\dp.rf.rf[3][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0630_));
 sky130_fd_sc_hd__mux4_1 _4281_ (.A0(\dp.rf.rf[12][25] ),
    .A1(\dp.rf.rf[13][25] ),
    .A2(\dp.rf.rf[14][25] ),
    .A3(\dp.rf.rf[15][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0631_));
 sky130_fd_sc_hd__mux4_1 _4282_ (.A0(\dp.rf.rf[4][25] ),
    .A1(\dp.rf.rf[5][25] ),
    .A2(\dp.rf.rf[6][25] ),
    .A3(\dp.rf.rf[7][25] ),
    .S0(net213),
    .S1(net277),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_1 _4283_ (.A0(_0629_),
    .A1(_0630_),
    .A2(_0631_),
    .A3(_0632_),
    .S0(_0103_),
    .S1(net15),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_0086_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_0628_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand2_2 _4286_ (.A(_0311_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__nor2_1 _4287_ (.A(_0138_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _4288_ (.A1(_0138_),
    .A2(_3629_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__xor2_1 _4289_ (.A(_0122_),
    .B(_0638_),
    .X(_3332_));
 sky130_fd_sc_hd__inv_1 _4290_ (.A(_3332_),
    .Y(_3336_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(\dp.rf.rf[22][25] ),
    .A1(\dp.rf.rf[23][25] ),
    .S(net210),
    .X(_0639_));
 sky130_fd_sc_hd__o21ai_0 _4292_ (.A1(_0148_),
    .A2(_0639_),
    .B1(_0337_),
    .Y(_0640_));
 sky130_fd_sc_hd__a221oi_1 _4293_ (.A1(\dp.rf.rf[19][25] ),
    .A2(net210),
    .B1(net201),
    .B2(\dp.rf.rf[18][25] ),
    .C1(net190),
    .Y(_0641_));
 sky130_fd_sc_hd__inv_1 _4294_ (.A(\dp.rf.rf[20][25] ),
    .Y(_0642_));
 sky130_fd_sc_hd__mux2i_1 _4295_ (.A0(\dp.rf.rf[17][25] ),
    .A1(\dp.rf.rf[21][25] ),
    .S(net208),
    .Y(_0643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_147 ();
 sky130_fd_sc_hd__a221oi_1 _4297_ (.A1(_0642_),
    .A2(net204),
    .B1(_0643_),
    .B2(net210),
    .C1(net8),
    .Y(_0645_));
 sky130_fd_sc_hd__o22ai_1 _4298_ (.A1(\dp.rf.rf[16][25] ),
    .A2(net181),
    .B1(_0645_),
    .B2(_0202_),
    .Y(_0646_));
 sky130_fd_sc_hd__o21ai_1 _4299_ (.A1(_0640_),
    .A2(_0641_),
    .B1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(\dp.rf.rf[30][25] ),
    .A1(\dp.rf.rf[31][25] ),
    .S(net209),
    .X(_0648_));
 sky130_fd_sc_hd__o21ai_0 _4301_ (.A1(_0148_),
    .A2(_0648_),
    .B1(net182),
    .Y(_0649_));
 sky130_fd_sc_hd__a221oi_1 _4302_ (.A1(\dp.rf.rf[27][25] ),
    .A2(net209),
    .B1(net201),
    .B2(\dp.rf.rf[26][25] ),
    .C1(net190),
    .Y(_0650_));
 sky130_fd_sc_hd__mux4_1 _4303_ (.A0(\dp.rf.rf[24][25] ),
    .A1(\dp.rf.rf[25][25] ),
    .A2(\dp.rf.rf[28][25] ),
    .A3(\dp.rf.rf[29][25] ),
    .S0(net209),
    .S1(net208),
    .X(_0651_));
 sky130_fd_sc_hd__a21oi_1 _4304_ (.A1(net205),
    .A2(_0651_),
    .B1(net198),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_1 _4305_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_146 ();
 sky130_fd_sc_hd__mux4_1 _4307_ (.A0(\dp.rf.rf[2][25] ),
    .A1(\dp.rf.rf[3][25] ),
    .A2(\dp.rf.rf[6][25] ),
    .A3(\dp.rf.rf[7][25] ),
    .S0(net209),
    .S1(net208),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_1 _4308_ (.A(net8),
    .B(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(\dp.rf.rf[1][25] ),
    .A1(\dp.rf.rf[5][25] ),
    .S(net208),
    .X(_0657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_145 ();
 sky130_fd_sc_hd__o221ai_1 _4311_ (.A1(\dp.rf.rf[4][25] ),
    .A2(_0528_),
    .B1(_0657_),
    .B2(_0245_),
    .C1(net205),
    .Y(_0659_));
 sky130_fd_sc_hd__a31oi_2 _4312_ (.A1(_0493_),
    .A2(_0656_),
    .A3(_0659_),
    .B1(_0271_),
    .Y(_0660_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__a221oi_1 _4315_ (.A1(\dp.rf.rf[11][25] ),
    .A2(net209),
    .B1(net201),
    .B2(\dp.rf.rf[10][25] ),
    .C1(net190),
    .Y(_0663_));
 sky130_fd_sc_hd__mux2i_1 _4316_ (.A0(\dp.rf.rf[14][25] ),
    .A1(\dp.rf.rf[15][25] ),
    .S(net209),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(net208),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand3_1 _4318_ (.A(net8),
    .B(_0119_),
    .C(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_141 ();
 sky130_fd_sc_hd__mux4_1 _4321_ (.A0(\dp.rf.rf[8][25] ),
    .A1(\dp.rf.rf[9][25] ),
    .A2(\dp.rf.rf[12][25] ),
    .A3(\dp.rf.rf[13][25] ),
    .S0(net209),
    .S1(net208),
    .X(_0669_));
 sky130_fd_sc_hd__a21oi_1 _4322_ (.A1(net205),
    .A2(_0669_),
    .B1(net198),
    .Y(_0670_));
 sky130_fd_sc_hd__o21ai_1 _4323_ (.A1(_0663_),
    .A2(_0666_),
    .B1(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a32oi_4 _4324_ (.A1(net188),
    .A2(_0647_),
    .A3(_0653_),
    .B1(_0660_),
    .B2(_0671_),
    .Y(_3335_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_140 ();
 sky130_fd_sc_hd__mux4_1 _4326_ (.A0(\dp.rf.rf[28][24] ),
    .A1(\dp.rf.rf[29][24] ),
    .A2(\dp.rf.rf[30][24] ),
    .A3(\dp.rf.rf[31][24] ),
    .S0(net212),
    .S1(net274),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(net16),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_139 ();
 sky130_fd_sc_hd__mux4_1 _4329_ (.A0(\dp.rf.rf[20][24] ),
    .A1(\dp.rf.rf[21][24] ),
    .A2(\dp.rf.rf[22][24] ),
    .A3(\dp.rf.rf[23][24] ),
    .S0(net212),
    .S1(net274),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_0103_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand3_1 _4331_ (.A(net15),
    .B(_0674_),
    .C(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__mux4_1 _4332_ (.A0(\dp.rf.rf[24][24] ),
    .A1(\dp.rf.rf[25][24] ),
    .A2(\dp.rf.rf[26][24] ),
    .A3(\dp.rf.rf[27][24] ),
    .S0(net212),
    .S1(net274),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(net16),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__mux4_1 _4334_ (.A0(\dp.rf.rf[16][24] ),
    .A1(\dp.rf.rf[17][24] ),
    .A2(\dp.rf.rf[18][24] ),
    .A3(\dp.rf.rf[19][24] ),
    .S0(net212),
    .S1(net274),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _4335_ (.A(_0103_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand3_1 _4336_ (.A(_0286_),
    .B(_0680_),
    .C(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_138 ();
 sky130_fd_sc_hd__mux4_1 _4338_ (.A0(\dp.rf.rf[12][24] ),
    .A1(\dp.rf.rf[13][24] ),
    .A2(\dp.rf.rf[14][24] ),
    .A3(\dp.rf.rf[15][24] ),
    .S0(net215),
    .S1(net14),
    .X(_0685_));
 sky130_fd_sc_hd__mux4_1 _4339_ (.A0(\dp.rf.rf[4][24] ),
    .A1(\dp.rf.rf[5][24] ),
    .A2(\dp.rf.rf[6][24] ),
    .A3(\dp.rf.rf[7][24] ),
    .S0(net215),
    .S1(net14),
    .X(_0686_));
 sky130_fd_sc_hd__mux2i_2 _4340_ (.A0(_0685_),
    .A1(_0686_),
    .S(_0103_),
    .Y(_0687_));
 sky130_fd_sc_hd__mux4_1 _4341_ (.A0(\dp.rf.rf[8][24] ),
    .A1(\dp.rf.rf[9][24] ),
    .A2(\dp.rf.rf[10][24] ),
    .A3(\dp.rf.rf[11][24] ),
    .S0(net215),
    .S1(net14),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _4342_ (.A(net16),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__mux4_1 _4343_ (.A0(\dp.rf.rf[0][24] ),
    .A1(\dp.rf.rf[1][24] ),
    .A2(\dp.rf.rf[2][24] ),
    .A3(\dp.rf.rf[3][24] ),
    .S0(net215),
    .S1(net14),
    .X(_0690_));
 sky130_fd_sc_hd__nand2_1 _4344_ (.A(_0103_),
    .B(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__and3_1 _4345_ (.A(_0286_),
    .B(_0689_),
    .C(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__a21oi_4 _4346_ (.A1(net15),
    .A2(_0687_),
    .B1(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__a32oi_4 _4347_ (.A1(net17),
    .A2(_0678_),
    .A3(_0683_),
    .B1(_0693_),
    .B2(_0290_),
    .Y(_0694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__o21ai_1 _4349_ (.A1(_0086_),
    .A2(_0119_),
    .B1(_0304_),
    .Y(_3625_));
 sky130_fd_sc_hd__nor2_1 _4350_ (.A(net179),
    .B(_3625_),
    .Y(_0696_));
 sky130_fd_sc_hd__a21oi_1 _4351_ (.A1(net179),
    .A2(_0694_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__xnor2_1 _4352_ (.A(_0122_),
    .B(_0697_),
    .Y(_3340_));
 sky130_fd_sc_hd__inv_1 _4353_ (.A(_3340_),
    .Y(_3344_));
 sky130_fd_sc_hd__mux2i_1 _4354_ (.A0(\dp.rf.rf[24][24] ),
    .A1(\dp.rf.rf[28][24] ),
    .S(net207),
    .Y(_0698_));
 sky130_fd_sc_hd__mux2i_1 _4355_ (.A0(\dp.rf.rf[25][24] ),
    .A1(\dp.rf.rf[29][24] ),
    .S(net207),
    .Y(_0699_));
 sky130_fd_sc_hd__o22ai_1 _4356_ (.A1(_0170_),
    .A2(_0698_),
    .B1(_0699_),
    .B2(_0415_),
    .Y(_0700_));
 sky130_fd_sc_hd__o21ai_1 _4357_ (.A1(_0145_),
    .A2(_0700_),
    .B1(net187),
    .Y(_0701_));
 sky130_fd_sc_hd__nand4_1 _4358_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[26][24] ),
    .Y(_0702_));
 sky130_fd_sc_hd__o2bb2ai_1 _4359_ (.A1_N(\dp.rf.rf[26][24] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__and2_0 _4360_ (.A(\dp.rf.rf[27][24] ),
    .B(net209),
    .X(_0704_));
 sky130_fd_sc_hd__mux2i_1 _4361_ (.A0(\dp.rf.rf[30][24] ),
    .A1(\dp.rf.rf[31][24] ),
    .S(net209),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_1 _4362_ (.A(net207),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__o311ai_4 _4363_ (.A1(net190),
    .A2(_0703_),
    .A3(_0704_),
    .B1(_0406_),
    .C1(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand4_1 _4364_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[18][24] ),
    .Y(_0708_));
 sky130_fd_sc_hd__o2bb2ai_1 _4365_ (.A1_N(\dp.rf.rf[18][24] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__and2_0 _4366_ (.A(\dp.rf.rf[19][24] ),
    .B(net209),
    .X(_0710_));
 sky130_fd_sc_hd__mux2i_1 _4367_ (.A0(\dp.rf.rf[22][24] ),
    .A1(\dp.rf.rf[23][24] ),
    .S(net209),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _4368_ (.A(net207),
    .B(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__o311ai_4 _4369_ (.A1(net190),
    .A2(_0709_),
    .A3(_0710_),
    .B1(_0712_),
    .C1(net182),
    .Y(_0713_));
 sky130_fd_sc_hd__inv_1 _4370_ (.A(\dp.rf.rf[20][24] ),
    .Y(_0714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__mux2i_1 _4372_ (.A0(\dp.rf.rf[17][24] ),
    .A1(\dp.rf.rf[21][24] ),
    .S(net207),
    .Y(_0716_));
 sky130_fd_sc_hd__a221oi_1 _4373_ (.A1(_0714_),
    .A2(net203),
    .B1(_0716_),
    .B2(net209),
    .C1(net8),
    .Y(_0717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__o22ai_2 _4375_ (.A1(\dp.rf.rf[16][24] ),
    .A2(net181),
    .B1(_0717_),
    .B2(net196),
    .Y(_0719_));
 sky130_fd_sc_hd__a22oi_4 _4376_ (.A1(_0701_),
    .A2(_0707_),
    .B1(_0713_),
    .B2(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand4_1 _4377_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[10][24] ),
    .Y(_0721_));
 sky130_fd_sc_hd__o2bb2ai_1 _4378_ (.A1_N(\dp.rf.rf[10][24] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__and2_0 _4379_ (.A(\dp.rf.rf[11][24] ),
    .B(net211),
    .X(_0723_));
 sky130_fd_sc_hd__mux2i_1 _4380_ (.A0(\dp.rf.rf[14][24] ),
    .A1(\dp.rf.rf[15][24] ),
    .S(net211),
    .Y(_0724_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(net207),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o311ai_2 _4382_ (.A1(net190),
    .A2(_0722_),
    .A3(_0723_),
    .B1(_0725_),
    .C1(net182),
    .Y(_0726_));
 sky130_fd_sc_hd__mux4_1 _4383_ (.A0(\dp.rf.rf[8][24] ),
    .A1(\dp.rf.rf[9][24] ),
    .A2(\dp.rf.rf[12][24] ),
    .A3(\dp.rf.rf[13][24] ),
    .S0(net211),
    .S1(net207),
    .X(_0727_));
 sky130_fd_sc_hd__a21oi_1 _4384_ (.A1(_0224_),
    .A2(_0727_),
    .B1(net198),
    .Y(_0728_));
 sky130_fd_sc_hd__mux4_1 _4385_ (.A0(\dp.rf.rf[2][24] ),
    .A1(\dp.rf.rf[3][24] ),
    .A2(\dp.rf.rf[6][24] ),
    .A3(\dp.rf.rf[7][24] ),
    .S0(net211),
    .S1(net207),
    .X(_0729_));
 sky130_fd_sc_hd__inv_1 _4386_ (.A(\dp.rf.rf[4][24] ),
    .Y(_0730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__mux2i_1 _4388_ (.A0(\dp.rf.rf[1][24] ),
    .A1(\dp.rf.rf[5][24] ),
    .S(net207),
    .Y(_0732_));
 sky130_fd_sc_hd__a221oi_1 _4389_ (.A1(_0730_),
    .A2(net204),
    .B1(_0732_),
    .B2(net211),
    .C1(net8),
    .Y(_0733_));
 sky130_fd_sc_hd__a211oi_2 _4390_ (.A1(net8),
    .A2(_0729_),
    .B1(_0733_),
    .C1(net195),
    .Y(_0734_));
 sky130_fd_sc_hd__a211oi_4 _4391_ (.A1(_0726_),
    .A2(_0728_),
    .B1(_0734_),
    .C1(_0271_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_8 _4392_ (.A(_0720_),
    .B(_0735_),
    .Y(_3343_));
 sky130_fd_sc_hd__o21ai_1 _4393_ (.A1(_0103_),
    .A2(_0119_),
    .B1(_0304_),
    .Y(_3621_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__mux4_1 _4395_ (.A0(\dp.rf.rf[24][23] ),
    .A1(\dp.rf.rf[25][23] ),
    .A2(\dp.rf.rf[26][23] ),
    .A3(\dp.rf.rf[27][23] ),
    .S0(net213),
    .S1(net274),
    .X(_0737_));
 sky130_fd_sc_hd__mux4_1 _4396_ (.A0(\dp.rf.rf[16][23] ),
    .A1(\dp.rf.rf[17][23] ),
    .A2(\dp.rf.rf[18][23] ),
    .A3(\dp.rf.rf[19][23] ),
    .S0(net215),
    .S1(net274),
    .X(_0738_));
 sky130_fd_sc_hd__mux4_1 _4397_ (.A0(\dp.rf.rf[28][23] ),
    .A1(\dp.rf.rf[29][23] ),
    .A2(\dp.rf.rf[30][23] ),
    .A3(\dp.rf.rf[31][23] ),
    .S0(net213),
    .S1(net274),
    .X(_0739_));
 sky130_fd_sc_hd__mux4_1 _4398_ (.A0(\dp.rf.rf[20][23] ),
    .A1(\dp.rf.rf[21][23] ),
    .A2(\dp.rf.rf[22][23] ),
    .A3(\dp.rf.rf[23][23] ),
    .S0(net215),
    .S1(net274),
    .X(_0740_));
 sky130_fd_sc_hd__mux4_1 _4399_ (.A0(_0737_),
    .A1(_0738_),
    .A2(_0739_),
    .A3(_0740_),
    .S0(_0103_),
    .S1(net15),
    .X(_0741_));
 sky130_fd_sc_hd__mux4_1 _4400_ (.A0(\dp.rf.rf[8][23] ),
    .A1(\dp.rf.rf[9][23] ),
    .A2(\dp.rf.rf[10][23] ),
    .A3(\dp.rf.rf[11][23] ),
    .S0(net215),
    .S1(net14),
    .X(_0742_));
 sky130_fd_sc_hd__mux4_1 _4401_ (.A0(\dp.rf.rf[0][23] ),
    .A1(\dp.rf.rf[1][23] ),
    .A2(\dp.rf.rf[2][23] ),
    .A3(\dp.rf.rf[3][23] ),
    .S0(net215),
    .S1(net14),
    .X(_0743_));
 sky130_fd_sc_hd__mux4_1 _4402_ (.A0(\dp.rf.rf[12][23] ),
    .A1(\dp.rf.rf[13][23] ),
    .A2(\dp.rf.rf[14][23] ),
    .A3(\dp.rf.rf[15][23] ),
    .S0(net215),
    .S1(net14),
    .X(_0744_));
 sky130_fd_sc_hd__mux4_1 _4403_ (.A0(\dp.rf.rf[4][23] ),
    .A1(\dp.rf.rf[5][23] ),
    .A2(\dp.rf.rf[6][23] ),
    .A3(\dp.rf.rf[7][23] ),
    .S0(net215),
    .S1(net14),
    .X(_0745_));
 sky130_fd_sc_hd__mux4_2 _4404_ (.A0(_0742_),
    .A1(_0743_),
    .A2(_0744_),
    .A3(_0745_),
    .S0(_0103_),
    .S1(net15),
    .X(_0746_));
 sky130_fd_sc_hd__mux2i_4 _4405_ (.A0(_0741_),
    .A1(_0746_),
    .S(_0086_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor3_1 _4406_ (.A(_0138_),
    .B(_0401_),
    .C(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__a21oi_1 _4407_ (.A1(_0138_),
    .A2(_3621_),
    .B1(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__xor2_1 _4408_ (.A(_0122_),
    .B(_0749_),
    .X(_3348_));
 sky130_fd_sc_hd__inv_1 _4409_ (.A(_3348_),
    .Y(_3352_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(\dp.rf.rf[22][23] ),
    .A1(\dp.rf.rf[23][23] ),
    .S(net211),
    .X(_0750_));
 sky130_fd_sc_hd__o21ai_0 _4411_ (.A1(_0148_),
    .A2(_0750_),
    .B1(net182),
    .Y(_0751_));
 sky130_fd_sc_hd__a221oi_1 _4412_ (.A1(\dp.rf.rf[19][23] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[18][23] ),
    .C1(net190),
    .Y(_0752_));
 sky130_fd_sc_hd__inv_1 _4413_ (.A(\dp.rf.rf[20][23] ),
    .Y(_0753_));
 sky130_fd_sc_hd__mux2i_1 _4414_ (.A0(\dp.rf.rf[17][23] ),
    .A1(\dp.rf.rf[21][23] ),
    .S(net207),
    .Y(_0754_));
 sky130_fd_sc_hd__a221oi_1 _4415_ (.A1(_0753_),
    .A2(net203),
    .B1(_0754_),
    .B2(net211),
    .C1(net8),
    .Y(_0755_));
 sky130_fd_sc_hd__o22ai_1 _4416_ (.A1(\dp.rf.rf[16][23] ),
    .A2(net180),
    .B1(_0755_),
    .B2(net195),
    .Y(_0756_));
 sky130_fd_sc_hd__o21ai_1 _4417_ (.A1(_0751_),
    .A2(_0752_),
    .B1(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__mux4_1 _4418_ (.A0(\dp.rf.rf[26][23] ),
    .A1(\dp.rf.rf[27][23] ),
    .A2(\dp.rf.rf[30][23] ),
    .A3(\dp.rf.rf[31][23] ),
    .S0(net211),
    .S1(net207),
    .X(_0758_));
 sky130_fd_sc_hd__mux2i_1 _4419_ (.A0(\dp.rf.rf[25][23] ),
    .A1(\dp.rf.rf[29][23] ),
    .S(net207),
    .Y(_0759_));
 sky130_fd_sc_hd__mux2i_1 _4420_ (.A0(\dp.rf.rf[24][23] ),
    .A1(\dp.rf.rf[28][23] ),
    .S(net207),
    .Y(_0760_));
 sky130_fd_sc_hd__o22ai_1 _4421_ (.A1(_0415_),
    .A2(_0759_),
    .B1(_0760_),
    .B2(_0170_),
    .Y(_0761_));
 sky130_fd_sc_hd__a211o_1 _4422_ (.A1(net8),
    .A2(_0758_),
    .B1(_0761_),
    .C1(net198),
    .X(_0762_));
 sky130_fd_sc_hd__nor2b_1 _4423_ (.A(net211),
    .B_N(\dp.rf.rf[14][23] ),
    .Y(_0763_));
 sky130_fd_sc_hd__a211oi_1 _4424_ (.A1(\dp.rf.rf[15][23] ),
    .A2(net211),
    .B1(_0148_),
    .C1(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__a221oi_1 _4425_ (.A1(\dp.rf.rf[11][23] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[10][23] ),
    .C1(net190),
    .Y(_0765_));
 sky130_fd_sc_hd__mux4_1 _4426_ (.A0(\dp.rf.rf[8][23] ),
    .A1(\dp.rf.rf[9][23] ),
    .A2(\dp.rf.rf[12][23] ),
    .A3(\dp.rf.rf[13][23] ),
    .S0(net211),
    .S1(net207),
    .X(_0766_));
 sky130_fd_sc_hd__a21oi_1 _4427_ (.A1(_0224_),
    .A2(_0766_),
    .B1(net198),
    .Y(_0767_));
 sky130_fd_sc_hd__o31ai_2 _4428_ (.A1(net192),
    .A2(_0764_),
    .A3(_0765_),
    .B1(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__mux4_1 _4429_ (.A0(\dp.rf.rf[2][23] ),
    .A1(\dp.rf.rf[3][23] ),
    .A2(\dp.rf.rf[6][23] ),
    .A3(\dp.rf.rf[7][23] ),
    .S0(net211),
    .S1(net207),
    .X(_0769_));
 sky130_fd_sc_hd__inv_1 _4430_ (.A(\dp.rf.rf[4][23] ),
    .Y(_0770_));
 sky130_fd_sc_hd__mux2i_1 _4431_ (.A0(\dp.rf.rf[1][23] ),
    .A1(\dp.rf.rf[5][23] ),
    .S(net207),
    .Y(_0771_));
 sky130_fd_sc_hd__a221oi_1 _4432_ (.A1(_0770_),
    .A2(net203),
    .B1(_0771_),
    .B2(net211),
    .C1(net8),
    .Y(_0772_));
 sky130_fd_sc_hd__a211oi_1 _4433_ (.A1(net8),
    .A2(_0769_),
    .B1(_0772_),
    .C1(net196),
    .Y(_0773_));
 sky130_fd_sc_hd__nor2_1 _4434_ (.A(_0271_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__a32oi_4 _4435_ (.A1(net188),
    .A2(_0757_),
    .A3(_0762_),
    .B1(_0768_),
    .B2(_0774_),
    .Y(_3351_));
 sky130_fd_sc_hd__mux4_1 _4436_ (.A0(\dp.rf.rf[28][22] ),
    .A1(\dp.rf.rf[29][22] ),
    .A2(\dp.rf.rf[30][22] ),
    .A3(\dp.rf.rf[31][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0775_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(net16),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__mux4_1 _4438_ (.A0(\dp.rf.rf[20][22] ),
    .A1(\dp.rf.rf[21][22] ),
    .A2(\dp.rf.rf[22][22] ),
    .A3(\dp.rf.rf[23][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _4439_ (.A(_0103_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand3_1 _4440_ (.A(net15),
    .B(_0776_),
    .C(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__mux4_1 _4441_ (.A0(\dp.rf.rf[24][22] ),
    .A1(\dp.rf.rf[25][22] ),
    .A2(\dp.rf.rf[26][22] ),
    .A3(\dp.rf.rf[27][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(net16),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__mux4_1 _4443_ (.A0(\dp.rf.rf[16][22] ),
    .A1(\dp.rf.rf[17][22] ),
    .A2(\dp.rf.rf[18][22] ),
    .A3(\dp.rf.rf[19][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _4444_ (.A(_0103_),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__nand3_1 _4445_ (.A(_0286_),
    .B(_0781_),
    .C(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__mux4_1 _4446_ (.A0(\dp.rf.rf[12][22] ),
    .A1(\dp.rf.rf[13][22] ),
    .A2(\dp.rf.rf[14][22] ),
    .A3(\dp.rf.rf[15][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0785_));
 sky130_fd_sc_hd__mux4_1 _4447_ (.A0(\dp.rf.rf[4][22] ),
    .A1(\dp.rf.rf[5][22] ),
    .A2(\dp.rf.rf[6][22] ),
    .A3(\dp.rf.rf[7][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0786_));
 sky130_fd_sc_hd__mux2i_1 _4448_ (.A0(_0785_),
    .A1(_0786_),
    .S(_0103_),
    .Y(_0787_));
 sky130_fd_sc_hd__mux4_1 _4449_ (.A0(\dp.rf.rf[8][22] ),
    .A1(\dp.rf.rf[9][22] ),
    .A2(\dp.rf.rf[10][22] ),
    .A3(\dp.rf.rf[11][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _4450_ (.A(net16),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__mux4_1 _4451_ (.A0(\dp.rf.rf[0][22] ),
    .A1(\dp.rf.rf[1][22] ),
    .A2(\dp.rf.rf[2][22] ),
    .A3(\dp.rf.rf[3][22] ),
    .S0(net13),
    .S1(net277),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _4452_ (.A(_0103_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__and3_1 _4453_ (.A(_0286_),
    .B(_0789_),
    .C(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__a21oi_2 _4454_ (.A1(net15),
    .A2(_0787_),
    .B1(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a32oi_4 _4455_ (.A1(net17),
    .A2(_0779_),
    .A3(_0784_),
    .B1(_0793_),
    .B2(net184),
    .Y(_0794_));
 sky130_fd_sc_hd__o21ai_1 _4456_ (.A1(_0286_),
    .A2(_0119_),
    .B1(_0304_),
    .Y(_3617_));
 sky130_fd_sc_hd__nor2_1 _4457_ (.A(net179),
    .B(_3617_),
    .Y(_0795_));
 sky130_fd_sc_hd__a21oi_1 _4458_ (.A1(net179),
    .A2(_0794_),
    .B1(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__xnor2_1 _4459_ (.A(_0122_),
    .B(_0796_),
    .Y(_3356_));
 sky130_fd_sc_hd__inv_1 _4460_ (.A(_3356_),
    .Y(_3360_));
 sky130_fd_sc_hd__mux4_1 _4461_ (.A0(\dp.rf.rf[10][22] ),
    .A1(\dp.rf.rf[11][22] ),
    .A2(\dp.rf.rf[14][22] ),
    .A3(\dp.rf.rf[15][22] ),
    .S0(net209),
    .S1(net208),
    .X(_0797_));
 sky130_fd_sc_hd__nand2_1 _4462_ (.A(net8),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__mux4_1 _4463_ (.A0(\dp.rf.rf[8][22] ),
    .A1(\dp.rf.rf[9][22] ),
    .A2(\dp.rf.rf[12][22] ),
    .A3(\dp.rf.rf[13][22] ),
    .S0(net209),
    .S1(net208),
    .X(_0799_));
 sky130_fd_sc_hd__nand2_1 _4464_ (.A(net205),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand3_2 _4465_ (.A(net185),
    .B(_0798_),
    .C(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(\dp.rf.rf[6][22] ),
    .A1(\dp.rf.rf[7][22] ),
    .S(net209),
    .X(_0802_));
 sky130_fd_sc_hd__o21ai_0 _4467_ (.A1(_0148_),
    .A2(_0802_),
    .B1(_0337_),
    .Y(_0803_));
 sky130_fd_sc_hd__a221oi_1 _4468_ (.A1(\dp.rf.rf[3][22] ),
    .A2(net209),
    .B1(net201),
    .B2(\dp.rf.rf[2][22] ),
    .C1(net189),
    .Y(_0804_));
 sky130_fd_sc_hd__inv_1 _4469_ (.A(\dp.rf.rf[4][22] ),
    .Y(_0805_));
 sky130_fd_sc_hd__mux2i_1 _4470_ (.A0(\dp.rf.rf[1][22] ),
    .A1(\dp.rf.rf[5][22] ),
    .S(net208),
    .Y(_0806_));
 sky130_fd_sc_hd__a221oi_1 _4471_ (.A1(_0805_),
    .A2(net204),
    .B1(_0806_),
    .B2(net209),
    .C1(net8),
    .Y(_0807_));
 sky130_fd_sc_hd__o22ai_1 _4472_ (.A1(\dp.rf.rf[0][22] ),
    .A2(net180),
    .B1(_0807_),
    .B2(net195),
    .Y(_0808_));
 sky130_fd_sc_hd__o21ai_2 _4473_ (.A1(_0803_),
    .A2(_0804_),
    .B1(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__mux2_1 _4474_ (.A0(\dp.rf.rf[26][22] ),
    .A1(\dp.rf.rf[27][22] ),
    .S(net210),
    .X(_0810_));
 sky130_fd_sc_hd__mux2i_1 _4475_ (.A0(\dp.rf.rf[30][22] ),
    .A1(\dp.rf.rf[31][22] ),
    .S(net210),
    .Y(_0811_));
 sky130_fd_sc_hd__a21oi_1 _4476_ (.A1(net208),
    .A2(_0811_),
    .B1(net205),
    .Y(_0812_));
 sky130_fd_sc_hd__o21ai_0 _4477_ (.A1(net189),
    .A2(_0810_),
    .B1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__mux4_1 _4478_ (.A0(\dp.rf.rf[24][22] ),
    .A1(\dp.rf.rf[25][22] ),
    .A2(\dp.rf.rf[28][22] ),
    .A3(\dp.rf.rf[29][22] ),
    .S0(net210),
    .S1(net208),
    .X(_0814_));
 sky130_fd_sc_hd__a21oi_1 _4479_ (.A1(net205),
    .A2(_0814_),
    .B1(_0192_),
    .Y(_0815_));
 sky130_fd_sc_hd__a21oi_1 _4480_ (.A1(_0813_),
    .A2(_0815_),
    .B1(_0166_),
    .Y(_0816_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(\dp.rf.rf[22][22] ),
    .A1(\dp.rf.rf[23][22] ),
    .S(net210),
    .X(_0817_));
 sky130_fd_sc_hd__o21ai_0 _4482_ (.A1(_0148_),
    .A2(_0817_),
    .B1(_0337_),
    .Y(_0818_));
 sky130_fd_sc_hd__a221oi_1 _4483_ (.A1(\dp.rf.rf[19][22] ),
    .A2(net210),
    .B1(net201),
    .B2(\dp.rf.rf[18][22] ),
    .C1(net189),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_1 _4484_ (.A(\dp.rf.rf[20][22] ),
    .Y(_0820_));
 sky130_fd_sc_hd__mux2i_1 _4485_ (.A0(\dp.rf.rf[17][22] ),
    .A1(\dp.rf.rf[21][22] ),
    .S(net208),
    .Y(_0821_));
 sky130_fd_sc_hd__a221oi_1 _4486_ (.A1(_0820_),
    .A2(net204),
    .B1(_0821_),
    .B2(net210),
    .C1(net8),
    .Y(_0822_));
 sky130_fd_sc_hd__o22ai_1 _4487_ (.A1(\dp.rf.rf[16][22] ),
    .A2(net180),
    .B1(_0822_),
    .B2(net195),
    .Y(_0823_));
 sky130_fd_sc_hd__o21ai_1 _4488_ (.A1(_0818_),
    .A2(_0819_),
    .B1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__a32oi_4 _4489_ (.A1(_0209_),
    .A2(_0801_),
    .A3(_0809_),
    .B1(_0816_),
    .B2(_0824_),
    .Y(_3359_));
 sky130_fd_sc_hd__o21ai_1 _4490_ (.A1(_0057_),
    .A2(_0119_),
    .B1(_0304_),
    .Y(_3613_));
 sky130_fd_sc_hd__mux4_1 _4491_ (.A0(\dp.rf.rf[24][21] ),
    .A1(\dp.rf.rf[25][21] ),
    .A2(\dp.rf.rf[26][21] ),
    .A3(\dp.rf.rf[27][21] ),
    .S0(net213),
    .S1(net278),
    .X(_0825_));
 sky130_fd_sc_hd__mux4_1 _4492_ (.A0(\dp.rf.rf[16][21] ),
    .A1(\dp.rf.rf[17][21] ),
    .A2(\dp.rf.rf[18][21] ),
    .A3(\dp.rf.rf[19][21] ),
    .S0(net213),
    .S1(net278),
    .X(_0826_));
 sky130_fd_sc_hd__mux4_1 _4493_ (.A0(\dp.rf.rf[28][21] ),
    .A1(\dp.rf.rf[29][21] ),
    .A2(\dp.rf.rf[30][21] ),
    .A3(\dp.rf.rf[31][21] ),
    .S0(net213),
    .S1(net278),
    .X(_0827_));
 sky130_fd_sc_hd__mux4_1 _4494_ (.A0(\dp.rf.rf[20][21] ),
    .A1(\dp.rf.rf[21][21] ),
    .A2(\dp.rf.rf[22][21] ),
    .A3(\dp.rf.rf[23][21] ),
    .S0(net213),
    .S1(net278),
    .X(_0828_));
 sky130_fd_sc_hd__mux4_1 _4495_ (.A0(_0825_),
    .A1(_0826_),
    .A2(_0827_),
    .A3(_0828_),
    .S0(_0103_),
    .S1(net15),
    .X(_0829_));
 sky130_fd_sc_hd__nand2_1 _4496_ (.A(net17),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__mux4_1 _4497_ (.A0(\dp.rf.rf[8][21] ),
    .A1(\dp.rf.rf[9][21] ),
    .A2(\dp.rf.rf[10][21] ),
    .A3(\dp.rf.rf[11][21] ),
    .S0(net215),
    .S1(net14),
    .X(_0831_));
 sky130_fd_sc_hd__mux4_1 _4498_ (.A0(\dp.rf.rf[0][21] ),
    .A1(\dp.rf.rf[1][21] ),
    .A2(\dp.rf.rf[2][21] ),
    .A3(\dp.rf.rf[3][21] ),
    .S0(net215),
    .S1(net14),
    .X(_0832_));
 sky130_fd_sc_hd__mux4_1 _4499_ (.A0(\dp.rf.rf[12][21] ),
    .A1(\dp.rf.rf[13][21] ),
    .A2(\dp.rf.rf[14][21] ),
    .A3(\dp.rf.rf[15][21] ),
    .S0(net215),
    .S1(net14),
    .X(_0833_));
 sky130_fd_sc_hd__mux4_1 _4500_ (.A0(\dp.rf.rf[4][21] ),
    .A1(\dp.rf.rf[5][21] ),
    .A2(\dp.rf.rf[6][21] ),
    .A3(\dp.rf.rf[7][21] ),
    .S0(net215),
    .S1(net14),
    .X(_0834_));
 sky130_fd_sc_hd__mux4_1 _4501_ (.A0(_0831_),
    .A1(_0832_),
    .A2(_0833_),
    .A3(_0834_),
    .S0(_0103_),
    .S1(net15),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _4502_ (.A(_0086_),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_2 _4503_ (.A(_0830_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2_4 _4504_ (.A(_0311_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_1 _4505_ (.A(_0138_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__a21oi_1 _4506_ (.A1(_0138_),
    .A2(_3613_),
    .B1(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__xor2_1 _4507_ (.A(_0122_),
    .B(_0840_),
    .X(_3364_));
 sky130_fd_sc_hd__inv_1 _4508_ (.A(_3364_),
    .Y(_3368_));
 sky130_fd_sc_hd__mux4_1 _4509_ (.A0(\dp.rf.rf[26][21] ),
    .A1(\dp.rf.rf[27][21] ),
    .A2(\dp.rf.rf[30][21] ),
    .A3(\dp.rf.rf[31][21] ),
    .S0(net7),
    .S1(net206),
    .X(_0841_));
 sky130_fd_sc_hd__mux4_1 _4510_ (.A0(\dp.rf.rf[24][21] ),
    .A1(\dp.rf.rf[25][21] ),
    .A2(\dp.rf.rf[28][21] ),
    .A3(\dp.rf.rf[29][21] ),
    .S0(net7),
    .S1(net206),
    .X(_0842_));
 sky130_fd_sc_hd__a221o_1 _4511_ (.A1(_0337_),
    .A2(_0841_),
    .B1(_0842_),
    .B2(_0224_),
    .C1(net198),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(\dp.rf.rf[22][21] ),
    .A1(\dp.rf.rf[23][21] ),
    .S(net7),
    .X(_0844_));
 sky130_fd_sc_hd__o21ai_0 _4513_ (.A1(_0148_),
    .A2(_0844_),
    .B1(_0337_),
    .Y(_0845_));
 sky130_fd_sc_hd__a221oi_1 _4514_ (.A1(\dp.rf.rf[19][21] ),
    .A2(net7),
    .B1(net201),
    .B2(\dp.rf.rf[18][21] ),
    .C1(net189),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_1 _4515_ (.A(\dp.rf.rf[20][21] ),
    .Y(_0847_));
 sky130_fd_sc_hd__mux2i_1 _4516_ (.A0(\dp.rf.rf[17][21] ),
    .A1(\dp.rf.rf[21][21] ),
    .S(net206),
    .Y(_0848_));
 sky130_fd_sc_hd__a221oi_1 _4517_ (.A1(_0847_),
    .A2(net204),
    .B1(_0848_),
    .B2(net7),
    .C1(net8),
    .Y(_0849_));
 sky130_fd_sc_hd__o22ai_1 _4518_ (.A1(\dp.rf.rf[16][21] ),
    .A2(net180),
    .B1(_0849_),
    .B2(net195),
    .Y(_0850_));
 sky130_fd_sc_hd__o21ai_1 _4519_ (.A1(_0845_),
    .A2(_0846_),
    .B1(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_132 ();
 sky130_fd_sc_hd__mux4_1 _4521_ (.A0(\dp.rf.rf[10][21] ),
    .A1(\dp.rf.rf[11][21] ),
    .A2(\dp.rf.rf[14][21] ),
    .A3(\dp.rf.rf[15][21] ),
    .S0(net211),
    .S1(net207),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_1 _4522_ (.A0(\dp.rf.rf[8][21] ),
    .A1(\dp.rf.rf[9][21] ),
    .A2(\dp.rf.rf[12][21] ),
    .A3(\dp.rf.rf[13][21] ),
    .S0(net211),
    .S1(net207),
    .X(_0854_));
 sky130_fd_sc_hd__mux2i_1 _4523_ (.A0(_0853_),
    .A1(_0854_),
    .S(_0224_),
    .Y(_0855_));
 sky130_fd_sc_hd__mux4_1 _4524_ (.A0(\dp.rf.rf[2][21] ),
    .A1(\dp.rf.rf[3][21] ),
    .A2(\dp.rf.rf[6][21] ),
    .A3(\dp.rf.rf[7][21] ),
    .S0(net211),
    .S1(net207),
    .X(_0856_));
 sky130_fd_sc_hd__inv_1 _4525_ (.A(\dp.rf.rf[4][21] ),
    .Y(_0857_));
 sky130_fd_sc_hd__mux2i_1 _4526_ (.A0(\dp.rf.rf[1][21] ),
    .A1(\dp.rf.rf[5][21] ),
    .S(net207),
    .Y(_0858_));
 sky130_fd_sc_hd__a221oi_1 _4527_ (.A1(_0857_),
    .A2(net204),
    .B1(_0858_),
    .B2(net211),
    .C1(net8),
    .Y(_0859_));
 sky130_fd_sc_hd__a211oi_1 _4528_ (.A1(net8),
    .A2(_0856_),
    .B1(_0859_),
    .C1(net195),
    .Y(_0860_));
 sky130_fd_sc_hd__a21oi_2 _4529_ (.A1(net185),
    .A2(_0855_),
    .B1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__a32oi_4 _4530_ (.A1(net188),
    .A2(_0843_),
    .A3(_0851_),
    .B1(_0861_),
    .B2(_0209_),
    .Y(_3367_));
 sky130_fd_sc_hd__mux4_1 _4531_ (.A0(\dp.rf.rf[28][20] ),
    .A1(\dp.rf.rf[29][20] ),
    .A2(\dp.rf.rf[30][20] ),
    .A3(\dp.rf.rf[31][20] ),
    .S0(net212),
    .S1(net274),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_1 _4532_ (.A(net16),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__mux4_1 _4533_ (.A0(\dp.rf.rf[20][20] ),
    .A1(\dp.rf.rf[21][20] ),
    .A2(\dp.rf.rf[22][20] ),
    .A3(\dp.rf.rf[23][20] ),
    .S0(net213),
    .S1(net274),
    .X(_0864_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_0103_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__nand3_1 _4535_ (.A(net15),
    .B(_0863_),
    .C(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__mux4_1 _4536_ (.A0(\dp.rf.rf[24][20] ),
    .A1(\dp.rf.rf[25][20] ),
    .A2(\dp.rf.rf[26][20] ),
    .A3(\dp.rf.rf[27][20] ),
    .S0(net212),
    .S1(net274),
    .X(_0867_));
 sky130_fd_sc_hd__nand2_1 _4537_ (.A(net16),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__mux4_1 _4538_ (.A0(\dp.rf.rf[16][20] ),
    .A1(\dp.rf.rf[17][20] ),
    .A2(\dp.rf.rf[18][20] ),
    .A3(\dp.rf.rf[19][20] ),
    .S0(net213),
    .S1(net274),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(_0103_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand3_1 _4540_ (.A(_0286_),
    .B(_0868_),
    .C(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__mux4_1 _4541_ (.A0(\dp.rf.rf[12][20] ),
    .A1(\dp.rf.rf[13][20] ),
    .A2(\dp.rf.rf[14][20] ),
    .A3(\dp.rf.rf[15][20] ),
    .S0(net215),
    .S1(net14),
    .X(_0872_));
 sky130_fd_sc_hd__mux4_1 _4542_ (.A0(\dp.rf.rf[4][20] ),
    .A1(\dp.rf.rf[5][20] ),
    .A2(\dp.rf.rf[6][20] ),
    .A3(\dp.rf.rf[7][20] ),
    .S0(net215),
    .S1(net274),
    .X(_0873_));
 sky130_fd_sc_hd__mux2i_1 _4543_ (.A0(_0872_),
    .A1(_0873_),
    .S(_0103_),
    .Y(_0874_));
 sky130_fd_sc_hd__mux4_1 _4544_ (.A0(\dp.rf.rf[8][20] ),
    .A1(\dp.rf.rf[9][20] ),
    .A2(\dp.rf.rf[10][20] ),
    .A3(\dp.rf.rf[11][20] ),
    .S0(net215),
    .S1(net14),
    .X(_0875_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(net16),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__mux4_1 _4546_ (.A0(\dp.rf.rf[0][20] ),
    .A1(\dp.rf.rf[1][20] ),
    .A2(\dp.rf.rf[2][20] ),
    .A3(\dp.rf.rf[3][20] ),
    .S0(net215),
    .S1(net274),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _4547_ (.A(_0103_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__and3_1 _4548_ (.A(_0286_),
    .B(_0876_),
    .C(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__a21oi_2 _4549_ (.A1(net15),
    .A2(_0874_),
    .B1(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__a32oi_4 _4550_ (.A1(net17),
    .A2(_0866_),
    .A3(_0871_),
    .B1(_0880_),
    .B2(_0290_),
    .Y(_0881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_130 ();
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(net213),
    .B(_0130_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_0304_),
    .B(_0884_),
    .Y(_3609_));
 sky130_fd_sc_hd__nor2_1 _4555_ (.A(net179),
    .B(_3609_),
    .Y(_0885_));
 sky130_fd_sc_hd__a21oi_1 _4556_ (.A1(net179),
    .A2(_0881_),
    .B1(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__xnor2_1 _4557_ (.A(_0122_),
    .B(_0886_),
    .Y(_3372_));
 sky130_fd_sc_hd__inv_1 _4558_ (.A(_3372_),
    .Y(_3376_));
 sky130_fd_sc_hd__mux2_1 _4559_ (.A0(\dp.rf.rf[22][20] ),
    .A1(\dp.rf.rf[23][20] ),
    .S(net211),
    .X(_0887_));
 sky130_fd_sc_hd__o21ai_0 _4560_ (.A1(_0148_),
    .A2(_0887_),
    .B1(net182),
    .Y(_0888_));
 sky130_fd_sc_hd__a221oi_1 _4561_ (.A1(\dp.rf.rf[19][20] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[18][20] ),
    .C1(net190),
    .Y(_0889_));
 sky130_fd_sc_hd__inv_1 _4562_ (.A(\dp.rf.rf[20][20] ),
    .Y(_0890_));
 sky130_fd_sc_hd__mux2i_1 _4563_ (.A0(\dp.rf.rf[17][20] ),
    .A1(\dp.rf.rf[21][20] ),
    .S(net206),
    .Y(_0891_));
 sky130_fd_sc_hd__a221oi_1 _4564_ (.A1(_0890_),
    .A2(net204),
    .B1(_0891_),
    .B2(net211),
    .C1(net8),
    .Y(_0892_));
 sky130_fd_sc_hd__o22ai_1 _4565_ (.A1(\dp.rf.rf[16][20] ),
    .A2(net180),
    .B1(_0892_),
    .B2(net195),
    .Y(_0893_));
 sky130_fd_sc_hd__o21ai_1 _4566_ (.A1(_0888_),
    .A2(_0889_),
    .B1(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__mux4_1 _4567_ (.A0(\dp.rf.rf[26][20] ),
    .A1(\dp.rf.rf[27][20] ),
    .A2(\dp.rf.rf[30][20] ),
    .A3(\dp.rf.rf[31][20] ),
    .S0(net211),
    .S1(net206),
    .X(_0895_));
 sky130_fd_sc_hd__mux2i_1 _4568_ (.A0(\dp.rf.rf[25][20] ),
    .A1(\dp.rf.rf[29][20] ),
    .S(net206),
    .Y(_0896_));
 sky130_fd_sc_hd__mux2i_1 _4569_ (.A0(\dp.rf.rf[24][20] ),
    .A1(\dp.rf.rf[28][20] ),
    .S(net206),
    .Y(_0897_));
 sky130_fd_sc_hd__o22ai_1 _4570_ (.A1(_0415_),
    .A2(_0896_),
    .B1(_0897_),
    .B2(_0170_),
    .Y(_0898_));
 sky130_fd_sc_hd__a211o_1 _4571_ (.A1(net8),
    .A2(_0895_),
    .B1(_0898_),
    .C1(net198),
    .X(_0899_));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(\dp.rf.rf[9][20] ),
    .A1(\dp.rf.rf[11][20] ),
    .A2(\dp.rf.rf[13][20] ),
    .A3(\dp.rf.rf[15][20] ),
    .S0(net8),
    .S1(net207),
    .X(_0900_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(net211),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__mux4_1 _4574_ (.A0(\dp.rf.rf[8][20] ),
    .A1(\dp.rf.rf[10][20] ),
    .A2(\dp.rf.rf[12][20] ),
    .A3(\dp.rf.rf[14][20] ),
    .S0(net8),
    .S1(net207),
    .X(_0902_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_0245_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a31oi_4 _4576_ (.A1(net185),
    .A2(_0901_),
    .A3(_0903_),
    .B1(_0271_),
    .Y(_0904_));
 sky130_fd_sc_hd__mux2_1 _4577_ (.A0(\dp.rf.rf[6][20] ),
    .A1(\dp.rf.rf[7][20] ),
    .S(net211),
    .X(_0905_));
 sky130_fd_sc_hd__o21ai_0 _4578_ (.A1(_0148_),
    .A2(_0905_),
    .B1(net182),
    .Y(_0906_));
 sky130_fd_sc_hd__a221oi_1 _4579_ (.A1(\dp.rf.rf[3][20] ),
    .A2(net211),
    .B1(net201),
    .B2(\dp.rf.rf[2][20] ),
    .C1(net190),
    .Y(_0907_));
 sky130_fd_sc_hd__inv_1 _4580_ (.A(\dp.rf.rf[4][20] ),
    .Y(_0908_));
 sky130_fd_sc_hd__mux2i_1 _4581_ (.A0(\dp.rf.rf[1][20] ),
    .A1(\dp.rf.rf[5][20] ),
    .S(net207),
    .Y(_0909_));
 sky130_fd_sc_hd__a221oi_1 _4582_ (.A1(_0908_),
    .A2(net204),
    .B1(_0909_),
    .B2(net211),
    .C1(net8),
    .Y(_0910_));
 sky130_fd_sc_hd__o22ai_1 _4583_ (.A1(\dp.rf.rf[0][20] ),
    .A2(net180),
    .B1(_0910_),
    .B2(net195),
    .Y(_0911_));
 sky130_fd_sc_hd__o21ai_2 _4584_ (.A1(_0906_),
    .A2(_0907_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__a32oi_4 _4585_ (.A1(net188),
    .A2(_0894_),
    .A3(_0899_),
    .B1(_0904_),
    .B2(_0912_),
    .Y(_3375_));
 sky130_fd_sc_hd__nand2_4 _4586_ (.A(net26),
    .B(_0128_),
    .Y(_0913_));
 sky130_fd_sc_hd__and3_2 _4587_ (.A(net25),
    .B(_0119_),
    .C(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__a221oi_2 _4589_ (.A1(net10),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net11),
    .C1(_0914_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand2_4 _4590_ (.A(_0120_),
    .B(_0913_),
    .Y(_0917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__and2_0 _4592_ (.A(net25),
    .B(_0119_),
    .X(_0919_));
 sky130_fd_sc_hd__a211oi_1 _4593_ (.A1(net11),
    .A2(_0130_),
    .B1(_0919_),
    .C1(_0917_),
    .Y(_0920_));
 sky130_fd_sc_hd__a21oi_1 _4594_ (.A1(_0916_),
    .A2(_0917_),
    .B1(_0920_),
    .Y(_3605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_126 ();
 sky130_fd_sc_hd__mux4_1 _4597_ (.A0(\dp.rf.rf[28][19] ),
    .A1(\dp.rf.rf[29][19] ),
    .A2(\dp.rf.rf[30][19] ),
    .A3(\dp.rf.rf[31][19] ),
    .S0(net212),
    .S1(net274),
    .X(_0923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__mux4_1 _4602_ (.A0(\dp.rf.rf[20][19] ),
    .A1(\dp.rf.rf[21][19] ),
    .A2(\dp.rf.rf[22][19] ),
    .A3(\dp.rf.rf[23][19] ),
    .S0(net212),
    .S1(net274),
    .X(_0928_));
 sky130_fd_sc_hd__a22oi_2 _4603_ (.A1(_0104_),
    .A2(_0923_),
    .B1(_0928_),
    .B2(_0102_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _4604_ (.A(_0103_),
    .B(_0064_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux4_1 _4605_ (.A0(\dp.rf.rf[12][19] ),
    .A1(\dp.rf.rf[13][19] ),
    .A2(\dp.rf.rf[14][19] ),
    .A3(\dp.rf.rf[15][19] ),
    .S0(net213),
    .S1(net274),
    .X(_0931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_120 ();
 sky130_fd_sc_hd__mux4_1 _4608_ (.A0(\dp.rf.rf[4][19] ),
    .A1(\dp.rf.rf[5][19] ),
    .A2(\dp.rf.rf[6][19] ),
    .A3(\dp.rf.rf[7][19] ),
    .S0(net213),
    .S1(net274),
    .X(_0934_));
 sky130_fd_sc_hd__nor2_2 _4609_ (.A(net16),
    .B(_0064_),
    .Y(_0935_));
 sky130_fd_sc_hd__a22oi_2 _4610_ (.A1(_0930_),
    .A2(_0931_),
    .B1(_0934_),
    .B2(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__mux2i_1 _4611_ (.A0(\dp.rf.rf[26][19] ),
    .A1(\dp.rf.rf[27][19] ),
    .S(net212),
    .Y(_0937_));
 sky130_fd_sc_hd__mux2i_1 _4612_ (.A0(\dp.rf.rf[24][19] ),
    .A1(\dp.rf.rf[25][19] ),
    .S(net212),
    .Y(_0938_));
 sky130_fd_sc_hd__a22oi_1 _4613_ (.A1(_0066_),
    .A2(_0937_),
    .B1(_0938_),
    .B2(_0061_),
    .Y(_0939_));
 sky130_fd_sc_hd__mux2i_1 _4614_ (.A0(\dp.rf.rf[18][19] ),
    .A1(\dp.rf.rf[19][19] ),
    .S(net212),
    .Y(_0940_));
 sky130_fd_sc_hd__mux2i_1 _4615_ (.A0(\dp.rf.rf[16][19] ),
    .A1(\dp.rf.rf[17][19] ),
    .S(net212),
    .Y(_0941_));
 sky130_fd_sc_hd__a22oi_1 _4616_ (.A1(_0081_),
    .A2(_0940_),
    .B1(_0941_),
    .B2(_0054_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand3_1 _4617_ (.A(_0088_),
    .B(_0939_),
    .C(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor3_1 _4618_ (.A(net17),
    .B(net15),
    .C(_0103_),
    .Y(_0944_));
 sky130_fd_sc_hd__mux4_1 _4619_ (.A0(\dp.rf.rf[8][19] ),
    .A1(\dp.rf.rf[9][19] ),
    .A2(\dp.rf.rf[10][19] ),
    .A3(\dp.rf.rf[11][19] ),
    .S0(net213),
    .S1(net274),
    .X(_0945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_119 ();
 sky130_fd_sc_hd__mux4_1 _4621_ (.A0(\dp.rf.rf[0][19] ),
    .A1(\dp.rf.rf[1][19] ),
    .A2(\dp.rf.rf[2][19] ),
    .A3(\dp.rf.rf[3][19] ),
    .S0(net213),
    .S1(net274),
    .X(_0947_));
 sky130_fd_sc_hd__nor4_4 _4622_ (.A(net17),
    .B(net15),
    .C(net16),
    .D(_0289_),
    .Y(_0948_));
 sky130_fd_sc_hd__a22oi_2 _4623_ (.A1(_0944_),
    .A2(_0945_),
    .B1(_0947_),
    .B2(_0948_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand4_4 _4624_ (.A(_0929_),
    .B(_0936_),
    .C(_0943_),
    .D(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__mux2i_1 _4625_ (.A0(_3605_),
    .A1(_0950_),
    .S(net179),
    .Y(_0951_));
 sky130_fd_sc_hd__xor2_1 _4626_ (.A(_0122_),
    .B(_0951_),
    .X(_3380_));
 sky130_fd_sc_hd__inv_1 _4627_ (.A(_3380_),
    .Y(_3384_));
 sky130_fd_sc_hd__nor2_4 _4628_ (.A(_0231_),
    .B(net196),
    .Y(_0952_));
 sky130_fd_sc_hd__mux4_1 _4629_ (.A0(\dp.rf.rf[18][19] ),
    .A1(\dp.rf.rf[19][19] ),
    .A2(\dp.rf.rf[22][19] ),
    .A3(\dp.rf.rf[23][19] ),
    .S0(net209),
    .S1(net206),
    .X(_0953_));
 sky130_fd_sc_hd__nand2_1 _4630_ (.A(net8),
    .B(_0953_),
    .Y(_0954_));
 sky130_fd_sc_hd__or2_4 _4631_ (.A(net210),
    .B(net208),
    .X(_0955_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_118 ();
 sky130_fd_sc_hd__nor2_1 _4633_ (.A(\dp.rf.rf[16][19] ),
    .B(_0955_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_1 _4634_ (.A(\dp.rf.rf[16][19] ),
    .B(_0119_),
    .Y(_0958_));
 sky130_fd_sc_hd__mux2_1 _4635_ (.A0(\dp.rf.rf[17][19] ),
    .A1(\dp.rf.rf[21][19] ),
    .S(net206),
    .X(_0959_));
 sky130_fd_sc_hd__o221ai_1 _4636_ (.A1(\dp.rf.rf[20][19] ),
    .A2(_0528_),
    .B1(_0959_),
    .B2(_0245_),
    .C1(net205),
    .Y(_0960_));
 sky130_fd_sc_hd__and3_1 _4637_ (.A(_0119_),
    .B(_0954_),
    .C(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__a211oi_2 _4638_ (.A1(_0954_),
    .A2(_0957_),
    .B1(_0958_),
    .C1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__nand2_4 _4639_ (.A(net11),
    .B(_0256_),
    .Y(_0963_));
 sky130_fd_sc_hd__mux4_1 _4640_ (.A0(\dp.rf.rf[26][19] ),
    .A1(\dp.rf.rf[27][19] ),
    .A2(\dp.rf.rf[30][19] ),
    .A3(\dp.rf.rf[31][19] ),
    .S0(net209),
    .S1(net206),
    .X(_0964_));
 sky130_fd_sc_hd__nor2_1 _4641_ (.A(net205),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__mux4_1 _4642_ (.A0(\dp.rf.rf[24][19] ),
    .A1(\dp.rf.rf[25][19] ),
    .A2(\dp.rf.rf[28][19] ),
    .A3(\dp.rf.rf[29][19] ),
    .S0(net209),
    .S1(net206),
    .X(_0966_));
 sky130_fd_sc_hd__nor2_1 _4643_ (.A(net8),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__nor3_1 _4644_ (.A(_0963_),
    .B(_0965_),
    .C(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__a21oi_4 _4645_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_0347_),
    .Y(_0969_));
 sky130_fd_sc_hd__inv_1 _4646_ (.A(\dp.rf.rf[12][19] ),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2i_1 _4647_ (.A0(\dp.rf.rf[9][19] ),
    .A1(\dp.rf.rf[13][19] ),
    .S(net206),
    .Y(_0971_));
 sky130_fd_sc_hd__a221oi_1 _4648_ (.A1(_0970_),
    .A2(net203),
    .B1(_0971_),
    .B2(net209),
    .C1(net8),
    .Y(_0972_));
 sky130_fd_sc_hd__o21ai_0 _4649_ (.A1(\dp.rf.rf[8][19] ),
    .A2(_0969_),
    .B1(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__mux4_1 _4650_ (.A0(\dp.rf.rf[10][19] ),
    .A1(\dp.rf.rf[11][19] ),
    .A2(\dp.rf.rf[14][19] ),
    .A3(\dp.rf.rf[15][19] ),
    .S0(net209),
    .S1(net206),
    .X(_0974_));
 sky130_fd_sc_hd__a21oi_1 _4651_ (.A1(net8),
    .A2(_0974_),
    .B1(net199),
    .Y(_0975_));
 sky130_fd_sc_hd__mux4_1 _4652_ (.A0(\dp.rf.rf[2][19] ),
    .A1(\dp.rf.rf[3][19] ),
    .A2(\dp.rf.rf[6][19] ),
    .A3(\dp.rf.rf[7][19] ),
    .S0(net209),
    .S1(net206),
    .X(_0976_));
 sky130_fd_sc_hd__and2_0 _4653_ (.A(net8),
    .B(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__inv_1 _4654_ (.A(\dp.rf.rf[4][19] ),
    .Y(_0978_));
 sky130_fd_sc_hd__mux2i_1 _4655_ (.A0(\dp.rf.rf[1][19] ),
    .A1(\dp.rf.rf[5][19] ),
    .S(net206),
    .Y(_0979_));
 sky130_fd_sc_hd__a221oi_1 _4656_ (.A1(_0978_),
    .A2(net203),
    .B1(_0979_),
    .B2(net209),
    .C1(net8),
    .Y(_0980_));
 sky130_fd_sc_hd__o31ai_1 _4657_ (.A1(net196),
    .A2(_0977_),
    .A3(_0980_),
    .B1(net194),
    .Y(_0981_));
 sky130_fd_sc_hd__a21oi_2 _4658_ (.A1(_0973_),
    .A2(_0975_),
    .B1(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a211oi_4 _4659_ (.A1(_0952_),
    .A2(_0962_),
    .B1(_0968_),
    .C1(_0982_),
    .Y(_3383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__mux4_1 _4662_ (.A0(\dp.rf.rf[28][18] ),
    .A1(\dp.rf.rf[29][18] ),
    .A2(\dp.rf.rf[30][18] ),
    .A3(\dp.rf.rf[31][18] ),
    .S0(net212),
    .S1(net274),
    .X(_0985_));
 sky130_fd_sc_hd__mux4_1 _4663_ (.A0(\dp.rf.rf[20][18] ),
    .A1(\dp.rf.rf[21][18] ),
    .A2(\dp.rf.rf[22][18] ),
    .A3(\dp.rf.rf[23][18] ),
    .S0(net212),
    .S1(net274),
    .X(_0986_));
 sky130_fd_sc_hd__a22oi_1 _4664_ (.A1(_0104_),
    .A2(_0985_),
    .B1(_0986_),
    .B2(_0102_),
    .Y(_0987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_115 ();
 sky130_fd_sc_hd__mux4_1 _4666_ (.A0(\dp.rf.rf[12][18] ),
    .A1(\dp.rf.rf[13][18] ),
    .A2(\dp.rf.rf[14][18] ),
    .A3(\dp.rf.rf[15][18] ),
    .S0(net212),
    .S1(net274),
    .X(_0989_));
 sky130_fd_sc_hd__mux4_1 _4667_ (.A0(\dp.rf.rf[4][18] ),
    .A1(\dp.rf.rf[5][18] ),
    .A2(\dp.rf.rf[6][18] ),
    .A3(\dp.rf.rf[7][18] ),
    .S0(net212),
    .S1(net274),
    .X(_0990_));
 sky130_fd_sc_hd__a22oi_1 _4668_ (.A1(_0930_),
    .A2(_0989_),
    .B1(_0990_),
    .B2(_0935_),
    .Y(_0991_));
 sky130_fd_sc_hd__mux2i_1 _4669_ (.A0(\dp.rf.rf[26][18] ),
    .A1(\dp.rf.rf[27][18] ),
    .S(net212),
    .Y(_0992_));
 sky130_fd_sc_hd__mux2i_1 _4670_ (.A0(\dp.rf.rf[24][18] ),
    .A1(\dp.rf.rf[25][18] ),
    .S(net212),
    .Y(_0993_));
 sky130_fd_sc_hd__a22oi_1 _4671_ (.A1(_0066_),
    .A2(_0992_),
    .B1(_0993_),
    .B2(_0061_),
    .Y(_0994_));
 sky130_fd_sc_hd__mux2i_1 _4672_ (.A0(\dp.rf.rf[18][18] ),
    .A1(\dp.rf.rf[19][18] ),
    .S(net212),
    .Y(_0995_));
 sky130_fd_sc_hd__mux2i_1 _4673_ (.A0(\dp.rf.rf[16][18] ),
    .A1(\dp.rf.rf[17][18] ),
    .S(net212),
    .Y(_0996_));
 sky130_fd_sc_hd__a22oi_1 _4674_ (.A1(_0081_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0054_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand3_1 _4675_ (.A(_0088_),
    .B(_0994_),
    .C(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__mux4_1 _4676_ (.A0(\dp.rf.rf[8][18] ),
    .A1(\dp.rf.rf[9][18] ),
    .A2(\dp.rf.rf[10][18] ),
    .A3(\dp.rf.rf[11][18] ),
    .S0(net212),
    .S1(net274),
    .X(_0999_));
 sky130_fd_sc_hd__mux4_1 _4677_ (.A0(\dp.rf.rf[0][18] ),
    .A1(\dp.rf.rf[1][18] ),
    .A2(\dp.rf.rf[2][18] ),
    .A3(\dp.rf.rf[3][18] ),
    .S0(net212),
    .S1(net274),
    .X(_1000_));
 sky130_fd_sc_hd__a22oi_1 _4678_ (.A1(_0944_),
    .A2(_0999_),
    .B1(_1000_),
    .B2(_0948_),
    .Y(_1001_));
 sky130_fd_sc_hd__and4_2 _4679_ (.A(_0987_),
    .B(_0991_),
    .C(_0998_),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__a221oi_2 _4680_ (.A1(net208),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net10),
    .C1(_0914_),
    .Y(_1003_));
 sky130_fd_sc_hd__mux2i_2 _4681_ (.A0(_0916_),
    .A1(_1003_),
    .S(_0917_),
    .Y(_3601_));
 sky130_fd_sc_hd__nor2_1 _4682_ (.A(net179),
    .B(_3601_),
    .Y(_1004_));
 sky130_fd_sc_hd__a21oi_1 _4683_ (.A1(net179),
    .A2(_1002_),
    .B1(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__xnor2_1 _4684_ (.A(_0122_),
    .B(_1005_),
    .Y(_3388_));
 sky130_fd_sc_hd__inv_1 _4685_ (.A(_3388_),
    .Y(_3392_));
 sky130_fd_sc_hd__inv_1 _4686_ (.A(\dp.rf.rf[28][18] ),
    .Y(_1006_));
 sky130_fd_sc_hd__mux2i_1 _4687_ (.A0(\dp.rf.rf[25][18] ),
    .A1(\dp.rf.rf[29][18] ),
    .S(net206),
    .Y(_1007_));
 sky130_fd_sc_hd__a221oi_1 _4688_ (.A1(_1006_),
    .A2(net203),
    .B1(_1007_),
    .B2(net209),
    .C1(net8),
    .Y(_1008_));
 sky130_fd_sc_hd__o22ai_2 _4689_ (.A1(\dp.rf.rf[24][18] ),
    .A2(_0969_),
    .B1(_1008_),
    .B2(_0130_),
    .Y(_1009_));
 sky130_fd_sc_hd__mux4_1 _4690_ (.A0(\dp.rf.rf[26][18] ),
    .A1(\dp.rf.rf[27][18] ),
    .A2(\dp.rf.rf[30][18] ),
    .A3(\dp.rf.rf[31][18] ),
    .S0(net209),
    .S1(net206),
    .X(_1010_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(net182),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__inv_1 _4692_ (.A(\dp.rf.rf[20][18] ),
    .Y(_1012_));
 sky130_fd_sc_hd__mux2i_1 _4693_ (.A0(\dp.rf.rf[17][18] ),
    .A1(\dp.rf.rf[21][18] ),
    .S(net206),
    .Y(_1013_));
 sky130_fd_sc_hd__a221oi_1 _4694_ (.A1(_1012_),
    .A2(net203),
    .B1(_1013_),
    .B2(net209),
    .C1(net8),
    .Y(_1014_));
 sky130_fd_sc_hd__o22ai_2 _4695_ (.A1(\dp.rf.rf[16][18] ),
    .A2(_0955_),
    .B1(_1014_),
    .B2(_0130_),
    .Y(_1015_));
 sky130_fd_sc_hd__mux4_1 _4696_ (.A0(\dp.rf.rf[18][18] ),
    .A1(\dp.rf.rf[19][18] ),
    .A2(\dp.rf.rf[22][18] ),
    .A3(\dp.rf.rf[23][18] ),
    .S0(net209),
    .S1(net206),
    .X(_1016_));
 sky130_fd_sc_hd__a21oi_1 _4697_ (.A1(net8),
    .A2(_1016_),
    .B1(net10),
    .Y(_1017_));
 sky130_fd_sc_hd__a32oi_4 _4698_ (.A1(net10),
    .A2(_1009_),
    .A3(_1011_),
    .B1(_1015_),
    .B2(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_1 _4699_ (.A(\dp.rf.rf[12][18] ),
    .Y(_1019_));
 sky130_fd_sc_hd__mux2i_1 _4700_ (.A0(\dp.rf.rf[9][18] ),
    .A1(\dp.rf.rf[13][18] ),
    .S(net206),
    .Y(_1020_));
 sky130_fd_sc_hd__a221oi_1 _4701_ (.A1(_1019_),
    .A2(net203),
    .B1(_1020_),
    .B2(net209),
    .C1(net8),
    .Y(_1021_));
 sky130_fd_sc_hd__o21ai_1 _4702_ (.A1(\dp.rf.rf[8][18] ),
    .A2(_0969_),
    .B1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__mux4_1 _4703_ (.A0(\dp.rf.rf[10][18] ),
    .A1(\dp.rf.rf[11][18] ),
    .A2(\dp.rf.rf[14][18] ),
    .A3(\dp.rf.rf[15][18] ),
    .S0(net209),
    .S1(net206),
    .X(_1023_));
 sky130_fd_sc_hd__a21oi_1 _4704_ (.A1(net8),
    .A2(_1023_),
    .B1(net199),
    .Y(_1024_));
 sky130_fd_sc_hd__mux4_1 _4705_ (.A0(\dp.rf.rf[2][18] ),
    .A1(\dp.rf.rf[3][18] ),
    .A2(\dp.rf.rf[6][18] ),
    .A3(\dp.rf.rf[7][18] ),
    .S0(net209),
    .S1(net206),
    .X(_1025_));
 sky130_fd_sc_hd__inv_1 _4706_ (.A(\dp.rf.rf[4][18] ),
    .Y(_1026_));
 sky130_fd_sc_hd__mux2i_1 _4707_ (.A0(\dp.rf.rf[1][18] ),
    .A1(\dp.rf.rf[5][18] ),
    .S(net206),
    .Y(_1027_));
 sky130_fd_sc_hd__a221oi_1 _4708_ (.A1(_1026_),
    .A2(net203),
    .B1(_1027_),
    .B2(net209),
    .C1(net8),
    .Y(_1028_));
 sky130_fd_sc_hd__a211oi_1 _4709_ (.A1(net8),
    .A2(_1025_),
    .B1(_1028_),
    .C1(net196),
    .Y(_1029_));
 sky130_fd_sc_hd__a21oi_2 _4710_ (.A1(_1022_),
    .A2(_1024_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__a22oi_4 _4711_ (.A1(net187),
    .A2(_1018_),
    .B1(_1030_),
    .B2(net194),
    .Y(_1031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_114 ();
 sky130_fd_sc_hd__mux2i_1 _4713_ (.A0(\dp.rf.rf[26][17] ),
    .A1(\dp.rf.rf[27][17] ),
    .S(net212),
    .Y(_1032_));
 sky130_fd_sc_hd__mux2i_1 _4714_ (.A0(\dp.rf.rf[24][17] ),
    .A1(\dp.rf.rf[25][17] ),
    .S(net212),
    .Y(_1033_));
 sky130_fd_sc_hd__a22oi_1 _4715_ (.A1(_0066_),
    .A2(_1032_),
    .B1(_1033_),
    .B2(_0061_),
    .Y(_1034_));
 sky130_fd_sc_hd__mux2i_1 _4716_ (.A0(\dp.rf.rf[18][17] ),
    .A1(\dp.rf.rf[19][17] ),
    .S(net212),
    .Y(_1035_));
 sky130_fd_sc_hd__mux2i_1 _4717_ (.A0(\dp.rf.rf[16][17] ),
    .A1(\dp.rf.rf[17][17] ),
    .S(net212),
    .Y(_1036_));
 sky130_fd_sc_hd__a22oi_1 _4718_ (.A1(_0081_),
    .A2(_1035_),
    .B1(_1036_),
    .B2(_0054_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand3_1 _4719_ (.A(_0088_),
    .B(_1034_),
    .C(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__inv_1 _4720_ (.A(\dp.rf.rf[4][17] ),
    .Y(_1039_));
 sky130_fd_sc_hd__nand2_1 _4721_ (.A(net212),
    .B(\dp.rf.rf[5][17] ),
    .Y(_1040_));
 sky130_fd_sc_hd__o211ai_1 _4722_ (.A1(net212),
    .A2(_1039_),
    .B1(_0054_),
    .C1(_1040_),
    .Y(_1041_));
 sky130_fd_sc_hd__mux2i_1 _4723_ (.A0(\dp.rf.rf[6][17] ),
    .A1(\dp.rf.rf[7][17] ),
    .S(net212),
    .Y(_1042_));
 sky130_fd_sc_hd__mux2i_1 _4724_ (.A0(\dp.rf.rf[12][17] ),
    .A1(\dp.rf.rf[13][17] ),
    .S(net212),
    .Y(_1043_));
 sky130_fd_sc_hd__a22oi_1 _4725_ (.A1(_0081_),
    .A2(_1042_),
    .B1(_1043_),
    .B2(_0061_),
    .Y(_1044_));
 sky130_fd_sc_hd__mux2i_1 _4726_ (.A0(\dp.rf.rf[14][17] ),
    .A1(\dp.rf.rf[15][17] ),
    .S(net212),
    .Y(_1045_));
 sky130_fd_sc_hd__a21oi_1 _4727_ (.A1(_0066_),
    .A2(_1045_),
    .B1(_0064_),
    .Y(_1046_));
 sky130_fd_sc_hd__nand3_1 _4728_ (.A(_1041_),
    .B(_1044_),
    .C(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__mux2i_1 _4729_ (.A0(\dp.rf.rf[8][17] ),
    .A1(\dp.rf.rf[9][17] ),
    .S(net212),
    .Y(_1048_));
 sky130_fd_sc_hd__mux2i_2 _4730_ (.A0(\dp.rf.rf[10][17] ),
    .A1(\dp.rf.rf[11][17] ),
    .S(net212),
    .Y(_1049_));
 sky130_fd_sc_hd__a22oi_1 _4731_ (.A1(_0061_),
    .A2(_1048_),
    .B1(_1049_),
    .B2(_0066_),
    .Y(_1050_));
 sky130_fd_sc_hd__mux2i_1 _4732_ (.A0(\dp.rf.rf[2][17] ),
    .A1(\dp.rf.rf[3][17] ),
    .S(net212),
    .Y(_1051_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0081_),
    .B(_1051_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(net212),
    .B(\dp.rf.rf[1][17] ),
    .Y(_1053_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_0054_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand4_1 _4736_ (.A(_0046_),
    .B(_1050_),
    .C(_1052_),
    .D(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__mux4_1 _4737_ (.A0(\dp.rf.rf[28][17] ),
    .A1(\dp.rf.rf[29][17] ),
    .A2(\dp.rf.rf[30][17] ),
    .A3(\dp.rf.rf[31][17] ),
    .S0(net212),
    .S1(net274),
    .X(_1056_));
 sky130_fd_sc_hd__mux4_1 _4738_ (.A0(\dp.rf.rf[20][17] ),
    .A1(\dp.rf.rf[21][17] ),
    .A2(\dp.rf.rf[22][17] ),
    .A3(\dp.rf.rf[23][17] ),
    .S0(net212),
    .S1(net274),
    .X(_1057_));
 sky130_fd_sc_hd__a22oi_2 _4739_ (.A1(_0104_),
    .A2(_1056_),
    .B1(_1057_),
    .B2(_0102_),
    .Y(_1058_));
 sky130_fd_sc_hd__nand4_4 _4740_ (.A(_1038_),
    .B(_1047_),
    .C(_1055_),
    .D(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__clkinvlp_4 _4741_ (.A(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand3_1 _4742_ (.A(net25),
    .B(_0119_),
    .C(_0913_),
    .Y(_1061_));
 sky130_fd_sc_hd__a22oi_1 _4743_ (.A1(net8),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net208),
    .Y(_1062_));
 sky130_fd_sc_hd__and3_1 _4744_ (.A(_1061_),
    .B(_0917_),
    .C(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__a31oi_2 _4745_ (.A1(_0120_),
    .A2(_0913_),
    .A3(_1003_),
    .B1(_1063_),
    .Y(_3597_));
 sky130_fd_sc_hd__nor2_1 _4746_ (.A(net179),
    .B(_3597_),
    .Y(_1064_));
 sky130_fd_sc_hd__a21oi_1 _4747_ (.A1(net179),
    .A2(_1060_),
    .B1(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__xnor2_1 _4748_ (.A(_0122_),
    .B(_1065_),
    .Y(_3396_));
 sky130_fd_sc_hd__inv_1 _4749_ (.A(_3396_),
    .Y(_3400_));
 sky130_fd_sc_hd__mux2i_1 _4750_ (.A0(\dp.rf.rf[18][17] ),
    .A1(\dp.rf.rf[22][17] ),
    .S(net206),
    .Y(_1066_));
 sky130_fd_sc_hd__o211ai_1 _4751_ (.A1(net205),
    .A2(_1066_),
    .B1(_0148_),
    .C1(_0245_),
    .Y(_1067_));
 sky130_fd_sc_hd__a21oi_1 _4752_ (.A1(_0119_),
    .A2(_1067_),
    .B1(\dp.rf.rf[16][17] ),
    .Y(_1068_));
 sky130_fd_sc_hd__mux2i_1 _4753_ (.A0(\dp.rf.rf[19][17] ),
    .A1(\dp.rf.rf[23][17] ),
    .S(net206),
    .Y(_1069_));
 sky130_fd_sc_hd__nand2_2 _4754_ (.A(net209),
    .B(net8),
    .Y(_1070_));
 sky130_fd_sc_hd__o22ai_1 _4755_ (.A1(_0247_),
    .A2(_1066_),
    .B1(_1069_),
    .B2(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__inv_1 _4756_ (.A(\dp.rf.rf[20][17] ),
    .Y(_1072_));
 sky130_fd_sc_hd__mux2i_1 _4757_ (.A0(\dp.rf.rf[17][17] ),
    .A1(\dp.rf.rf[21][17] ),
    .S(net206),
    .Y(_1073_));
 sky130_fd_sc_hd__a221oi_1 _4758_ (.A1(_1072_),
    .A2(net203),
    .B1(_1073_),
    .B2(net209),
    .C1(net8),
    .Y(_1074_));
 sky130_fd_sc_hd__nor3_1 _4759_ (.A(_0130_),
    .B(_1071_),
    .C(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__nor4_1 _4760_ (.A(_0231_),
    .B(net196),
    .C(_1068_),
    .D(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__mux4_1 _4761_ (.A0(\dp.rf.rf[26][17] ),
    .A1(\dp.rf.rf[27][17] ),
    .A2(\dp.rf.rf[30][17] ),
    .A3(\dp.rf.rf[31][17] ),
    .S0(net209),
    .S1(net206),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(net8),
    .B(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__inv_1 _4763_ (.A(\dp.rf.rf[28][17] ),
    .Y(_1079_));
 sky130_fd_sc_hd__mux2i_1 _4764_ (.A0(\dp.rf.rf[25][17] ),
    .A1(\dp.rf.rf[29][17] ),
    .S(net206),
    .Y(_1080_));
 sky130_fd_sc_hd__a221oi_1 _4765_ (.A1(_1079_),
    .A2(net203),
    .B1(_1080_),
    .B2(net209),
    .C1(net8),
    .Y(_1081_));
 sky130_fd_sc_hd__o22ai_1 _4766_ (.A1(\dp.rf.rf[24][17] ),
    .A2(_0955_),
    .B1(_1081_),
    .B2(_0130_),
    .Y(_1082_));
 sky130_fd_sc_hd__a21oi_1 _4767_ (.A1(_1078_),
    .A2(_1082_),
    .B1(_0963_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux2i_1 _4768_ (.A0(\dp.rf.rf[9][17] ),
    .A1(\dp.rf.rf[13][17] ),
    .S(net206),
    .Y(_1084_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(net209),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__o22a_1 _4770_ (.A1(\dp.rf.rf[12][17] ),
    .A2(_0528_),
    .B1(_0955_),
    .B2(\dp.rf.rf[8][17] ),
    .X(_1086_));
 sky130_fd_sc_hd__mux2i_1 _4771_ (.A0(\dp.rf.rf[11][17] ),
    .A1(\dp.rf.rf[15][17] ),
    .S(net206),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2i_1 _4772_ (.A0(\dp.rf.rf[10][17] ),
    .A1(\dp.rf.rf[14][17] ),
    .S(net206),
    .Y(_1088_));
 sky130_fd_sc_hd__o22ai_1 _4773_ (.A1(_1070_),
    .A2(_1087_),
    .B1(_1088_),
    .B2(_0247_),
    .Y(_1089_));
 sky130_fd_sc_hd__a31oi_1 _4774_ (.A1(net205),
    .A2(_1085_),
    .A3(_1086_),
    .B1(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__mux4_1 _4775_ (.A0(\dp.rf.rf[2][17] ),
    .A1(\dp.rf.rf[3][17] ),
    .A2(\dp.rf.rf[6][17] ),
    .A3(\dp.rf.rf[7][17] ),
    .S0(net209),
    .S1(net206),
    .X(_1091_));
 sky130_fd_sc_hd__and2_0 _4776_ (.A(net8),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2i_1 _4777_ (.A0(\dp.rf.rf[1][17] ),
    .A1(\dp.rf.rf[5][17] ),
    .S(net206),
    .Y(_1093_));
 sky130_fd_sc_hd__a221oi_1 _4778_ (.A1(_1039_),
    .A2(net203),
    .B1(_1093_),
    .B2(net209),
    .C1(net8),
    .Y(_1094_));
 sky130_fd_sc_hd__nor3_1 _4779_ (.A(net210),
    .B(net8),
    .C(net208),
    .Y(_1095_));
 sky130_fd_sc_hd__a2111oi_4 _4780_ (.A1(_0115_),
    .A2(_0117_),
    .B1(_1095_),
    .C1(net11),
    .D1(net10),
    .Y(_1096_));
 sky130_fd_sc_hd__o21ai_0 _4781_ (.A1(_1092_),
    .A2(_1094_),
    .B1(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__o31ai_1 _4782_ (.A1(net11),
    .A2(net199),
    .A3(_1090_),
    .B1(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__or3_4 _4783_ (.A(_1076_),
    .B(_1083_),
    .C(_1098_),
    .X(_3395_));
 sky130_fd_sc_hd__clkinv_4 _4784_ (.A(_3395_),
    .Y(_3399_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_113 ();
 sky130_fd_sc_hd__mux2i_2 _4786_ (.A0(\dp.rf.rf[26][16] ),
    .A1(\dp.rf.rf[27][16] ),
    .S(net212),
    .Y(_1100_));
 sky130_fd_sc_hd__mux2i_1 _4787_ (.A0(\dp.rf.rf[24][16] ),
    .A1(\dp.rf.rf[25][16] ),
    .S(net212),
    .Y(_1101_));
 sky130_fd_sc_hd__a22oi_1 _4788_ (.A1(_0066_),
    .A2(_1100_),
    .B1(_1101_),
    .B2(_0061_),
    .Y(_1102_));
 sky130_fd_sc_hd__mux2i_1 _4789_ (.A0(\dp.rf.rf[18][16] ),
    .A1(\dp.rf.rf[19][16] ),
    .S(net212),
    .Y(_1103_));
 sky130_fd_sc_hd__mux2i_1 _4790_ (.A0(\dp.rf.rf[16][16] ),
    .A1(\dp.rf.rf[17][16] ),
    .S(net212),
    .Y(_1104_));
 sky130_fd_sc_hd__a22oi_1 _4791_ (.A1(_0081_),
    .A2(_1103_),
    .B1(_1104_),
    .B2(_0054_),
    .Y(_1105_));
 sky130_fd_sc_hd__nand3_1 _4792_ (.A(_0088_),
    .B(_1102_),
    .C(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__inv_1 _4793_ (.A(\dp.rf.rf[4][16] ),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(net212),
    .B(\dp.rf.rf[5][16] ),
    .Y(_1108_));
 sky130_fd_sc_hd__o211ai_1 _4795_ (.A1(net212),
    .A2(_1107_),
    .B1(_0054_),
    .C1(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__mux2i_1 _4796_ (.A0(\dp.rf.rf[6][16] ),
    .A1(\dp.rf.rf[7][16] ),
    .S(net212),
    .Y(_1110_));
 sky130_fd_sc_hd__mux2i_1 _4797_ (.A0(\dp.rf.rf[12][16] ),
    .A1(\dp.rf.rf[13][16] ),
    .S(net212),
    .Y(_1111_));
 sky130_fd_sc_hd__a22oi_1 _4798_ (.A1(_0081_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(_0061_),
    .Y(_1112_));
 sky130_fd_sc_hd__mux2i_1 _4799_ (.A0(\dp.rf.rf[14][16] ),
    .A1(\dp.rf.rf[15][16] ),
    .S(net212),
    .Y(_1113_));
 sky130_fd_sc_hd__a21oi_1 _4800_ (.A1(_0066_),
    .A2(_1113_),
    .B1(_0064_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand3_1 _4801_ (.A(_1109_),
    .B(_1112_),
    .C(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__mux2i_1 _4802_ (.A0(\dp.rf.rf[8][16] ),
    .A1(\dp.rf.rf[9][16] ),
    .S(net212),
    .Y(_1116_));
 sky130_fd_sc_hd__mux2i_1 _4803_ (.A0(\dp.rf.rf[10][16] ),
    .A1(\dp.rf.rf[11][16] ),
    .S(net212),
    .Y(_1117_));
 sky130_fd_sc_hd__a22oi_1 _4804_ (.A1(_0061_),
    .A2(_1116_),
    .B1(_1117_),
    .B2(_0066_),
    .Y(_1118_));
 sky130_fd_sc_hd__mux2i_1 _4805_ (.A0(\dp.rf.rf[2][16] ),
    .A1(\dp.rf.rf[3][16] ),
    .S(net212),
    .Y(_1119_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_0081_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(net212),
    .B(\dp.rf.rf[1][16] ),
    .Y(_1121_));
 sky130_fd_sc_hd__nand2_1 _4808_ (.A(_0054_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand4_1 _4809_ (.A(_0046_),
    .B(_1118_),
    .C(_1120_),
    .D(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__mux4_1 _4810_ (.A0(\dp.rf.rf[28][16] ),
    .A1(\dp.rf.rf[29][16] ),
    .A2(\dp.rf.rf[30][16] ),
    .A3(\dp.rf.rf[31][16] ),
    .S0(net212),
    .S1(net274),
    .X(_1124_));
 sky130_fd_sc_hd__mux4_1 _4811_ (.A0(\dp.rf.rf[20][16] ),
    .A1(\dp.rf.rf[21][16] ),
    .A2(\dp.rf.rf[22][16] ),
    .A3(\dp.rf.rf[23][16] ),
    .S0(net212),
    .S1(net274),
    .X(_1125_));
 sky130_fd_sc_hd__a22oi_1 _4812_ (.A1(_0104_),
    .A2(_1124_),
    .B1(_1125_),
    .B2(_0102_),
    .Y(_1126_));
 sky130_fd_sc_hd__and4_2 _4813_ (.A(_1106_),
    .B(_1115_),
    .C(_1123_),
    .D(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__a221oi_4 _4814_ (.A1(net210),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net8),
    .C1(_0914_),
    .Y(_1128_));
 sky130_fd_sc_hd__nor3b_1 _4815_ (.A(_0914_),
    .B(_0917_),
    .C_N(_1062_),
    .Y(_1129_));
 sky130_fd_sc_hd__a21oi_1 _4816_ (.A1(_0917_),
    .A2(_1128_),
    .B1(_1129_),
    .Y(_3593_));
 sky130_fd_sc_hd__nor2_1 _4817_ (.A(net178),
    .B(_3593_),
    .Y(_1130_));
 sky130_fd_sc_hd__a21oi_1 _4818_ (.A1(net178),
    .A2(_1127_),
    .B1(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__xnor2_1 _4819_ (.A(_0122_),
    .B(_1131_),
    .Y(_3404_));
 sky130_fd_sc_hd__inv_1 _4820_ (.A(_3404_),
    .Y(_3408_));
 sky130_fd_sc_hd__mux2i_1 _4821_ (.A0(\dp.rf.rf[9][16] ),
    .A1(\dp.rf.rf[13][16] ),
    .S(net206),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(net209),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__o22a_1 _4823_ (.A1(\dp.rf.rf[12][16] ),
    .A2(_0528_),
    .B1(_0955_),
    .B2(\dp.rf.rf[8][16] ),
    .X(_1134_));
 sky130_fd_sc_hd__mux2i_1 _4824_ (.A0(\dp.rf.rf[11][16] ),
    .A1(\dp.rf.rf[15][16] ),
    .S(net206),
    .Y(_1135_));
 sky130_fd_sc_hd__mux2i_1 _4825_ (.A0(\dp.rf.rf[10][16] ),
    .A1(\dp.rf.rf[14][16] ),
    .S(net206),
    .Y(_1136_));
 sky130_fd_sc_hd__o22ai_1 _4826_ (.A1(_1070_),
    .A2(_1135_),
    .B1(_1136_),
    .B2(_0247_),
    .Y(_1137_));
 sky130_fd_sc_hd__a31oi_2 _4827_ (.A1(net205),
    .A2(_1133_),
    .A3(_1134_),
    .B1(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__mux4_1 _4828_ (.A0(\dp.rf.rf[2][16] ),
    .A1(\dp.rf.rf[3][16] ),
    .A2(\dp.rf.rf[6][16] ),
    .A3(\dp.rf.rf[7][16] ),
    .S0(net209),
    .S1(net206),
    .X(_1139_));
 sky130_fd_sc_hd__and2_0 _4829_ (.A(net8),
    .B(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__mux2i_1 _4830_ (.A0(\dp.rf.rf[1][16] ),
    .A1(\dp.rf.rf[5][16] ),
    .S(net206),
    .Y(_1141_));
 sky130_fd_sc_hd__a221oi_1 _4831_ (.A1(_1107_),
    .A2(net203),
    .B1(_1141_),
    .B2(net209),
    .C1(net8),
    .Y(_1142_));
 sky130_fd_sc_hd__o21ai_1 _4832_ (.A1(_1140_),
    .A2(_1142_),
    .B1(_1096_),
    .Y(_1143_));
 sky130_fd_sc_hd__o31ai_4 _4833_ (.A1(net11),
    .A2(net199),
    .A3(_1138_),
    .B1(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__inv_1 _4834_ (.A(\dp.rf.rf[28][16] ),
    .Y(_1145_));
 sky130_fd_sc_hd__mux2i_1 _4835_ (.A0(\dp.rf.rf[25][16] ),
    .A1(\dp.rf.rf[29][16] ),
    .S(net206),
    .Y(_1146_));
 sky130_fd_sc_hd__a221oi_2 _4836_ (.A1(_1145_),
    .A2(net203),
    .B1(_1146_),
    .B2(net209),
    .C1(net8),
    .Y(_1147_));
 sky130_fd_sc_hd__o22ai_2 _4837_ (.A1(\dp.rf.rf[24][16] ),
    .A2(_0969_),
    .B1(_1147_),
    .B2(_0130_),
    .Y(_1148_));
 sky130_fd_sc_hd__mux4_1 _4838_ (.A0(\dp.rf.rf[26][16] ),
    .A1(\dp.rf.rf[27][16] ),
    .A2(\dp.rf.rf[30][16] ),
    .A3(\dp.rf.rf[31][16] ),
    .S0(net209),
    .S1(net206),
    .X(_1149_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(net182),
    .B(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__mux2i_1 _4840_ (.A0(\dp.rf.rf[18][16] ),
    .A1(\dp.rf.rf[22][16] ),
    .S(net206),
    .Y(_1151_));
 sky130_fd_sc_hd__mux2i_1 _4841_ (.A0(\dp.rf.rf[19][16] ),
    .A1(\dp.rf.rf[23][16] ),
    .S(net206),
    .Y(_1152_));
 sky130_fd_sc_hd__o221ai_1 _4842_ (.A1(_0247_),
    .A2(_1151_),
    .B1(_1152_),
    .B2(_1070_),
    .C1(_0145_),
    .Y(_1153_));
 sky130_fd_sc_hd__mux2i_1 _4843_ (.A0(\dp.rf.rf[17][16] ),
    .A1(\dp.rf.rf[21][16] ),
    .S(net206),
    .Y(_1154_));
 sky130_fd_sc_hd__nor3b_1 _4844_ (.A(\dp.rf.rf[20][16] ),
    .B(net209),
    .C_N(net206),
    .Y(_1155_));
 sky130_fd_sc_hd__nor3_1 _4845_ (.A(\dp.rf.rf[16][16] ),
    .B(net209),
    .C(net206),
    .Y(_1156_));
 sky130_fd_sc_hd__a2111oi_1 _4846_ (.A1(net209),
    .A2(_1154_),
    .B1(_1155_),
    .C1(_1156_),
    .D1(net8),
    .Y(_1157_));
 sky130_fd_sc_hd__o21ai_1 _4847_ (.A1(_1153_),
    .A2(_1157_),
    .B1(net187),
    .Y(_1158_));
 sky130_fd_sc_hd__a31oi_4 _4848_ (.A1(net10),
    .A2(_1148_),
    .A3(_1150_),
    .B1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__or2_4 _4849_ (.A(_1144_),
    .B(_1159_),
    .X(_3403_));
 sky130_fd_sc_hd__clkinv_2 _4850_ (.A(_3403_),
    .Y(_3407_));
 sky130_fd_sc_hd__mux4_1 _4851_ (.A0(\dp.rf.rf[24][15] ),
    .A1(\dp.rf.rf[25][15] ),
    .A2(\dp.rf.rf[26][15] ),
    .A3(\dp.rf.rf[27][15] ),
    .S0(net213),
    .S1(net278),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _4852_ (.A0(\dp.rf.rf[16][15] ),
    .A1(\dp.rf.rf[17][15] ),
    .A2(\dp.rf.rf[18][15] ),
    .A3(\dp.rf.rf[19][15] ),
    .S0(net213),
    .S1(net278),
    .X(_1161_));
 sky130_fd_sc_hd__mux4_1 _4853_ (.A0(\dp.rf.rf[28][15] ),
    .A1(\dp.rf.rf[29][15] ),
    .A2(\dp.rf.rf[30][15] ),
    .A3(\dp.rf.rf[31][15] ),
    .S0(net213),
    .S1(net278),
    .X(_1162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_112 ();
 sky130_fd_sc_hd__mux4_1 _4855_ (.A0(\dp.rf.rf[20][15] ),
    .A1(\dp.rf.rf[21][15] ),
    .A2(\dp.rf.rf[22][15] ),
    .A3(\dp.rf.rf[23][15] ),
    .S0(net213),
    .S1(net278),
    .X(_1164_));
 sky130_fd_sc_hd__mux4_1 _4856_ (.A0(_1160_),
    .A1(_1161_),
    .A2(_1162_),
    .A3(_1164_),
    .S0(_0103_),
    .S1(net15),
    .X(_1165_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(net17),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__mux4_1 _4858_ (.A0(\dp.rf.rf[8][15] ),
    .A1(\dp.rf.rf[9][15] ),
    .A2(\dp.rf.rf[10][15] ),
    .A3(\dp.rf.rf[11][15] ),
    .S0(net215),
    .S1(net14),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_1 _4859_ (.A0(\dp.rf.rf[0][15] ),
    .A1(\dp.rf.rf[1][15] ),
    .A2(\dp.rf.rf[2][15] ),
    .A3(\dp.rf.rf[3][15] ),
    .S0(net215),
    .S1(net14),
    .X(_1168_));
 sky130_fd_sc_hd__mux4_1 _4860_ (.A0(\dp.rf.rf[12][15] ),
    .A1(\dp.rf.rf[13][15] ),
    .A2(\dp.rf.rf[14][15] ),
    .A3(\dp.rf.rf[15][15] ),
    .S0(net215),
    .S1(net14),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\dp.rf.rf[4][15] ),
    .A1(\dp.rf.rf[5][15] ),
    .A2(\dp.rf.rf[6][15] ),
    .A3(\dp.rf.rf[7][15] ),
    .S0(net215),
    .S1(net14),
    .X(_1170_));
 sky130_fd_sc_hd__mux4_1 _4862_ (.A0(_1167_),
    .A1(_1168_),
    .A2(_1169_),
    .A3(_1170_),
    .S0(_0103_),
    .S1(net15),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_0086_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_1166_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2_4 _4865_ (.A(_0311_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__a221oi_4 _4867_ (.A1(net6),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net210),
    .C1(_0914_),
    .Y(_1176_));
 sky130_fd_sc_hd__mux2i_4 _4868_ (.A0(_1128_),
    .A1(_1176_),
    .S(_0917_),
    .Y(_3589_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_0138_),
    .B(_3589_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21ai_0 _4870_ (.A1(_0138_),
    .A2(_1174_),
    .B1(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__xnor2_1 _4871_ (.A(_0122_),
    .B(_1178_),
    .Y(_3412_));
 sky130_fd_sc_hd__inv_1 _4872_ (.A(_3412_),
    .Y(_3416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__mux4_1 _4874_ (.A0(\dp.rf.rf[26][15] ),
    .A1(\dp.rf.rf[27][15] ),
    .A2(\dp.rf.rf[30][15] ),
    .A3(\dp.rf.rf[31][15] ),
    .S0(net7),
    .S1(net206),
    .X(_1180_));
 sky130_fd_sc_hd__mux4_1 _4875_ (.A0(\dp.rf.rf[24][15] ),
    .A1(\dp.rf.rf[25][15] ),
    .A2(\dp.rf.rf[28][15] ),
    .A3(\dp.rf.rf[29][15] ),
    .S0(net7),
    .S1(net206),
    .X(_1181_));
 sky130_fd_sc_hd__a221oi_1 _4876_ (.A1(_0337_),
    .A2(_1180_),
    .B1(_1181_),
    .B2(_0224_),
    .C1(net198),
    .Y(_1182_));
 sky130_fd_sc_hd__nor2_1 _4877_ (.A(_0166_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(\dp.rf.rf[22][15] ),
    .A1(\dp.rf.rf[23][15] ),
    .S(net7),
    .X(_1184_));
 sky130_fd_sc_hd__o21ai_0 _4879_ (.A1(_0148_),
    .A2(_1184_),
    .B1(_0337_),
    .Y(_1185_));
 sky130_fd_sc_hd__a221oi_1 _4880_ (.A1(\dp.rf.rf[19][15] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[18][15] ),
    .C1(net189),
    .Y(_1186_));
 sky130_fd_sc_hd__inv_1 _4881_ (.A(\dp.rf.rf[20][15] ),
    .Y(_1187_));
 sky130_fd_sc_hd__mux2i_1 _4882_ (.A0(\dp.rf.rf[17][15] ),
    .A1(\dp.rf.rf[21][15] ),
    .S(net206),
    .Y(_1188_));
 sky130_fd_sc_hd__a221oi_1 _4883_ (.A1(_1187_),
    .A2(net204),
    .B1(_1188_),
    .B2(net7),
    .C1(net8),
    .Y(_1189_));
 sky130_fd_sc_hd__o22ai_1 _4884_ (.A1(\dp.rf.rf[16][15] ),
    .A2(net180),
    .B1(_1189_),
    .B2(_0202_),
    .Y(_1190_));
 sky130_fd_sc_hd__o21ai_1 _4885_ (.A1(_1185_),
    .A2(_1186_),
    .B1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__mux4_1 _4886_ (.A0(\dp.rf.rf[2][15] ),
    .A1(\dp.rf.rf[3][15] ),
    .A2(\dp.rf.rf[6][15] ),
    .A3(\dp.rf.rf[7][15] ),
    .S0(net211),
    .S1(net207),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(net8),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__mux2_1 _4888_ (.A0(\dp.rf.rf[1][15] ),
    .A1(\dp.rf.rf[5][15] ),
    .S(net207),
    .X(_1194_));
 sky130_fd_sc_hd__o221ai_1 _4889_ (.A1(\dp.rf.rf[4][15] ),
    .A2(_0528_),
    .B1(_1194_),
    .B2(_0245_),
    .C1(_0224_),
    .Y(_1195_));
 sky130_fd_sc_hd__a31o_1 _4890_ (.A1(_0493_),
    .A2(_1193_),
    .A3(_1195_),
    .B1(_0271_),
    .X(_1196_));
 sky130_fd_sc_hd__mux2i_1 _4891_ (.A0(\dp.rf.rf[14][15] ),
    .A1(\dp.rf.rf[15][15] ),
    .S(net211),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_1 _4892_ (.A(net207),
    .B(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__a221o_1 _4893_ (.A1(\dp.rf.rf[11][15] ),
    .A2(net211),
    .B1(net200),
    .B2(\dp.rf.rf[10][15] ),
    .C1(net189),
    .X(_1199_));
 sky130_fd_sc_hd__mux4_1 _4894_ (.A0(\dp.rf.rf[8][15] ),
    .A1(\dp.rf.rf[9][15] ),
    .A2(\dp.rf.rf[12][15] ),
    .A3(\dp.rf.rf[13][15] ),
    .S0(net211),
    .S1(net207),
    .X(_1200_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(_0224_),
    .B(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _4896_ (.A(net185),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a31oi_4 _4897_ (.A1(_0337_),
    .A2(_1198_),
    .A3(_1199_),
    .B1(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__o2bb2ai_4 _4898_ (.A1_N(_1183_),
    .A2_N(_1191_),
    .B1(_1196_),
    .B2(_1203_),
    .Y(_3411_));
 sky130_fd_sc_hd__clkinv_2 _4899_ (.A(_3411_),
    .Y(_3415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_109 ();
 sky130_fd_sc_hd__a22oi_1 _4901_ (.A1(net5),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net6),
    .Y(_1205_));
 sky130_fd_sc_hd__and3_1 _4902_ (.A(_1061_),
    .B(_0917_),
    .C(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a31oi_4 _4903_ (.A1(_0120_),
    .A2(_0913_),
    .A3(_1176_),
    .B1(_1206_),
    .Y(_3585_));
 sky130_fd_sc_hd__nor2_1 _4904_ (.A(_0132_),
    .B(_3585_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux4_1 _4905_ (.A0(\dp.rf.rf[24][14] ),
    .A1(\dp.rf.rf[25][14] ),
    .A2(\dp.rf.rf[26][14] ),
    .A3(\dp.rf.rf[27][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1208_));
 sky130_fd_sc_hd__mux4_1 _4906_ (.A0(\dp.rf.rf[16][14] ),
    .A1(\dp.rf.rf[17][14] ),
    .A2(\dp.rf.rf[18][14] ),
    .A3(\dp.rf.rf[19][14] ),
    .S0(net214),
    .S1(net277),
    .X(_1209_));
 sky130_fd_sc_hd__mux4_1 _4907_ (.A0(\dp.rf.rf[28][14] ),
    .A1(\dp.rf.rf[29][14] ),
    .A2(\dp.rf.rf[30][14] ),
    .A3(\dp.rf.rf[31][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1210_));
 sky130_fd_sc_hd__mux4_1 _4908_ (.A0(\dp.rf.rf[20][14] ),
    .A1(\dp.rf.rf[21][14] ),
    .A2(\dp.rf.rf[22][14] ),
    .A3(\dp.rf.rf[23][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1211_));
 sky130_fd_sc_hd__mux4_1 _4909_ (.A0(_1208_),
    .A1(_1209_),
    .A2(_1210_),
    .A3(_1211_),
    .S0(_0103_),
    .S1(net15),
    .X(_1212_));
 sky130_fd_sc_hd__mux4_1 _4910_ (.A0(\dp.rf.rf[8][14] ),
    .A1(\dp.rf.rf[9][14] ),
    .A2(\dp.rf.rf[10][14] ),
    .A3(\dp.rf.rf[11][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1213_));
 sky130_fd_sc_hd__mux4_1 _4911_ (.A0(\dp.rf.rf[0][14] ),
    .A1(\dp.rf.rf[1][14] ),
    .A2(\dp.rf.rf[2][14] ),
    .A3(\dp.rf.rf[3][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1214_));
 sky130_fd_sc_hd__mux4_1 _4912_ (.A0(\dp.rf.rf[12][14] ),
    .A1(\dp.rf.rf[13][14] ),
    .A2(\dp.rf.rf[14][14] ),
    .A3(\dp.rf.rf[15][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1215_));
 sky130_fd_sc_hd__mux4_1 _4913_ (.A0(\dp.rf.rf[4][14] ),
    .A1(\dp.rf.rf[5][14] ),
    .A2(\dp.rf.rf[6][14] ),
    .A3(\dp.rf.rf[7][14] ),
    .S0(net214),
    .S1(net278),
    .X(_1216_));
 sky130_fd_sc_hd__mux4_1 _4914_ (.A0(_1213_),
    .A1(_1214_),
    .A2(_1215_),
    .A3(_1216_),
    .S0(_0103_),
    .S1(net15),
    .X(_1217_));
 sky130_fd_sc_hd__a22o_2 _4915_ (.A1(net17),
    .A2(_1212_),
    .B1(_1217_),
    .B2(net184),
    .X(_1218_));
 sky130_fd_sc_hd__nor2_1 _4916_ (.A(_0138_),
    .B(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__nor2_1 _4917_ (.A(_1207_),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__xnor2_1 _4918_ (.A(_0122_),
    .B(_1220_),
    .Y(_3420_));
 sky130_fd_sc_hd__inv_1 _4919_ (.A(_3420_),
    .Y(_3424_));
 sky130_fd_sc_hd__mux4_1 _4920_ (.A0(\dp.rf.rf[10][14] ),
    .A1(\dp.rf.rf[11][14] ),
    .A2(\dp.rf.rf[14][14] ),
    .A3(\dp.rf.rf[15][14] ),
    .S0(net7),
    .S1(net9),
    .X(_1221_));
 sky130_fd_sc_hd__nand2_1 _4921_ (.A(net8),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__mux4_1 _4922_ (.A0(\dp.rf.rf[8][14] ),
    .A1(\dp.rf.rf[9][14] ),
    .A2(\dp.rf.rf[12][14] ),
    .A3(\dp.rf.rf[13][14] ),
    .S0(net7),
    .S1(net9),
    .X(_1223_));
 sky130_fd_sc_hd__nand2_1 _4923_ (.A(net205),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand3_1 _4924_ (.A(net186),
    .B(_1222_),
    .C(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__mux2_1 _4925_ (.A0(\dp.rf.rf[6][14] ),
    .A1(\dp.rf.rf[7][14] ),
    .S(net7),
    .X(_1226_));
 sky130_fd_sc_hd__o21ai_0 _4926_ (.A1(_0148_),
    .A2(_1226_),
    .B1(net183),
    .Y(_1227_));
 sky130_fd_sc_hd__a221oi_1 _4927_ (.A1(\dp.rf.rf[3][14] ),
    .A2(net7),
    .B1(_0176_),
    .B2(\dp.rf.rf[2][14] ),
    .C1(net191),
    .Y(_1228_));
 sky130_fd_sc_hd__inv_1 _4928_ (.A(\dp.rf.rf[4][14] ),
    .Y(_1229_));
 sky130_fd_sc_hd__mux2i_1 _4929_ (.A0(\dp.rf.rf[1][14] ),
    .A1(\dp.rf.rf[5][14] ),
    .S(net9),
    .Y(_1230_));
 sky130_fd_sc_hd__a221oi_1 _4930_ (.A1(_1229_),
    .A2(_0263_),
    .B1(_1230_),
    .B2(net7),
    .C1(net8),
    .Y(_1231_));
 sky130_fd_sc_hd__o22ai_1 _4931_ (.A1(\dp.rf.rf[0][14] ),
    .A2(_0348_),
    .B1(_1231_),
    .B2(net197),
    .Y(_1232_));
 sky130_fd_sc_hd__o21ai_0 _4932_ (.A1(_1227_),
    .A2(_1228_),
    .B1(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__mux4_1 _4933_ (.A0(\dp.rf.rf[26][14] ),
    .A1(\dp.rf.rf[27][14] ),
    .A2(\dp.rf.rf[30][14] ),
    .A3(\dp.rf.rf[31][14] ),
    .S0(net7),
    .S1(net9),
    .X(_1234_));
 sky130_fd_sc_hd__nand2_1 _4934_ (.A(net8),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__mux4_1 _4935_ (.A0(\dp.rf.rf[24][14] ),
    .A1(\dp.rf.rf[25][14] ),
    .A2(\dp.rf.rf[28][14] ),
    .A3(\dp.rf.rf[29][14] ),
    .S0(net7),
    .S1(net9),
    .X(_1236_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(net205),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__a31oi_1 _4937_ (.A1(net10),
    .A2(_1235_),
    .A3(_1237_),
    .B1(_0166_),
    .Y(_1238_));
 sky130_fd_sc_hd__mux2_1 _4938_ (.A0(\dp.rf.rf[22][14] ),
    .A1(\dp.rf.rf[23][14] ),
    .S(net7),
    .X(_1239_));
 sky130_fd_sc_hd__o21ai_0 _4939_ (.A1(_0148_),
    .A2(_1239_),
    .B1(net183),
    .Y(_1240_));
 sky130_fd_sc_hd__a221oi_1 _4940_ (.A1(\dp.rf.rf[19][14] ),
    .A2(net7),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][14] ),
    .C1(net191),
    .Y(_1241_));
 sky130_fd_sc_hd__inv_1 _4941_ (.A(\dp.rf.rf[20][14] ),
    .Y(_1242_));
 sky130_fd_sc_hd__mux2i_1 _4942_ (.A0(\dp.rf.rf[17][14] ),
    .A1(\dp.rf.rf[21][14] ),
    .S(net9),
    .Y(_1243_));
 sky130_fd_sc_hd__a221oi_1 _4943_ (.A1(_1242_),
    .A2(_0263_),
    .B1(_1243_),
    .B2(net7),
    .C1(net8),
    .Y(_1244_));
 sky130_fd_sc_hd__o22ai_1 _4944_ (.A1(\dp.rf.rf[16][14] ),
    .A2(_0348_),
    .B1(_1244_),
    .B2(net197),
    .Y(_1245_));
 sky130_fd_sc_hd__o21ai_0 _4945_ (.A1(_1240_),
    .A2(_1241_),
    .B1(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__a32o_4 _4946_ (.A1(net193),
    .A2(_1225_),
    .A3(_1233_),
    .B1(_1238_),
    .B2(_1246_),
    .X(_3419_));
 sky130_fd_sc_hd__inv_2 _4947_ (.A(_3419_),
    .Y(_3423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_107 ();
 sky130_fd_sc_hd__a221oi_1 _4950_ (.A1(net4),
    .A2(_0130_),
    .B1(_0133_),
    .B2(net5),
    .C1(_0914_),
    .Y(_1249_));
 sky130_fd_sc_hd__nor3b_1 _4951_ (.A(_0914_),
    .B(_0917_),
    .C_N(_1205_),
    .Y(_1250_));
 sky130_fd_sc_hd__a21oi_2 _4952_ (.A1(_0917_),
    .A2(_1249_),
    .B1(_1250_),
    .Y(_3581_));
 sky130_fd_sc_hd__nor2_1 _4953_ (.A(_0132_),
    .B(_3581_),
    .Y(_1251_));
 sky130_fd_sc_hd__mux4_1 _4954_ (.A0(\dp.rf.rf[24][13] ),
    .A1(\dp.rf.rf[25][13] ),
    .A2(\dp.rf.rf[26][13] ),
    .A3(\dp.rf.rf[27][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1252_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\dp.rf.rf[16][13] ),
    .A1(\dp.rf.rf[17][13] ),
    .A2(\dp.rf.rf[18][13] ),
    .A3(\dp.rf.rf[19][13] ),
    .S0(net214),
    .S1(net277),
    .X(_1253_));
 sky130_fd_sc_hd__mux4_1 _4956_ (.A0(\dp.rf.rf[28][13] ),
    .A1(\dp.rf.rf[29][13] ),
    .A2(\dp.rf.rf[30][13] ),
    .A3(\dp.rf.rf[31][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1254_));
 sky130_fd_sc_hd__mux4_1 _4957_ (.A0(\dp.rf.rf[20][13] ),
    .A1(\dp.rf.rf[21][13] ),
    .A2(\dp.rf.rf[22][13] ),
    .A3(\dp.rf.rf[23][13] ),
    .S0(net214),
    .S1(net277),
    .X(_1255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_106 ();
 sky130_fd_sc_hd__mux4_1 _4959_ (.A0(_1252_),
    .A1(_1253_),
    .A2(_1254_),
    .A3(_1255_),
    .S0(_0103_),
    .S1(net15),
    .X(_1257_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_105 ();
 sky130_fd_sc_hd__mux4_1 _4961_ (.A0(\dp.rf.rf[8][13] ),
    .A1(\dp.rf.rf[9][13] ),
    .A2(\dp.rf.rf[10][13] ),
    .A3(\dp.rf.rf[11][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1259_));
 sky130_fd_sc_hd__mux4_1 _4962_ (.A0(\dp.rf.rf[0][13] ),
    .A1(\dp.rf.rf[1][13] ),
    .A2(\dp.rf.rf[2][13] ),
    .A3(\dp.rf.rf[3][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1260_));
 sky130_fd_sc_hd__mux4_1 _4963_ (.A0(\dp.rf.rf[12][13] ),
    .A1(\dp.rf.rf[13][13] ),
    .A2(\dp.rf.rf[14][13] ),
    .A3(\dp.rf.rf[15][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1261_));
 sky130_fd_sc_hd__mux4_1 _4964_ (.A0(\dp.rf.rf[4][13] ),
    .A1(\dp.rf.rf[5][13] ),
    .A2(\dp.rf.rf[6][13] ),
    .A3(\dp.rf.rf[7][13] ),
    .S0(net214),
    .S1(net278),
    .X(_1262_));
 sky130_fd_sc_hd__mux4_1 _4965_ (.A0(_1259_),
    .A1(_1260_),
    .A2(_1261_),
    .A3(_1262_),
    .S0(_0103_),
    .S1(net15),
    .X(_1263_));
 sky130_fd_sc_hd__a22o_2 _4966_ (.A1(net17),
    .A2(_1257_),
    .B1(_1263_),
    .B2(net184),
    .X(_1264_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_0138_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__nor2_1 _4968_ (.A(_1251_),
    .B(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__xnor2_1 _4969_ (.A(_0122_),
    .B(_1266_),
    .Y(_3428_));
 sky130_fd_sc_hd__inv_1 _4970_ (.A(_3428_),
    .Y(_3432_));
 sky130_fd_sc_hd__mux4_1 _4971_ (.A0(\dp.rf.rf[26][13] ),
    .A1(\dp.rf.rf[27][13] ),
    .A2(\dp.rf.rf[30][13] ),
    .A3(\dp.rf.rf[31][13] ),
    .S0(net7),
    .S1(net9),
    .X(_1267_));
 sky130_fd_sc_hd__mux4_1 _4972_ (.A0(\dp.rf.rf[24][13] ),
    .A1(\dp.rf.rf[25][13] ),
    .A2(\dp.rf.rf[28][13] ),
    .A3(\dp.rf.rf[29][13] ),
    .S0(net7),
    .S1(net9),
    .X(_1268_));
 sky130_fd_sc_hd__a221oi_1 _4973_ (.A1(net183),
    .A2(_1267_),
    .B1(_1268_),
    .B2(net205),
    .C1(net199),
    .Y(_1269_));
 sky130_fd_sc_hd__nor2_1 _4974_ (.A(_0166_),
    .B(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(\dp.rf.rf[22][13] ),
    .A1(\dp.rf.rf[23][13] ),
    .S(net7),
    .X(_1271_));
 sky130_fd_sc_hd__o21ai_0 _4976_ (.A1(_0148_),
    .A2(_1271_),
    .B1(net183),
    .Y(_1272_));
 sky130_fd_sc_hd__a221oi_1 _4977_ (.A1(\dp.rf.rf[19][13] ),
    .A2(net7),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][13] ),
    .C1(net191),
    .Y(_1273_));
 sky130_fd_sc_hd__inv_1 _4978_ (.A(\dp.rf.rf[20][13] ),
    .Y(_1274_));
 sky130_fd_sc_hd__mux2i_1 _4979_ (.A0(\dp.rf.rf[17][13] ),
    .A1(\dp.rf.rf[21][13] ),
    .S(net9),
    .Y(_1275_));
 sky130_fd_sc_hd__a221oi_1 _4980_ (.A1(_1274_),
    .A2(_0263_),
    .B1(_1275_),
    .B2(net7),
    .C1(net8),
    .Y(_1276_));
 sky130_fd_sc_hd__o22ai_1 _4981_ (.A1(\dp.rf.rf[16][13] ),
    .A2(_0348_),
    .B1(_1276_),
    .B2(net197),
    .Y(_1277_));
 sky130_fd_sc_hd__o21ai_0 _4982_ (.A1(_1272_),
    .A2(_1273_),
    .B1(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__mux4_1 _4983_ (.A0(\dp.rf.rf[10][13] ),
    .A1(\dp.rf.rf[11][13] ),
    .A2(\dp.rf.rf[14][13] ),
    .A3(\dp.rf.rf[15][13] ),
    .S0(net7),
    .S1(net9),
    .X(_1279_));
 sky130_fd_sc_hd__mux4_1 _4984_ (.A0(\dp.rf.rf[8][13] ),
    .A1(\dp.rf.rf[9][13] ),
    .A2(\dp.rf.rf[12][13] ),
    .A3(\dp.rf.rf[13][13] ),
    .S0(net7),
    .S1(net9),
    .X(_1280_));
 sky130_fd_sc_hd__mux2i_2 _4985_ (.A0(_1279_),
    .A1(_1280_),
    .S(net205),
    .Y(_1281_));
 sky130_fd_sc_hd__mux4_1 _4986_ (.A0(\dp.rf.rf[2][13] ),
    .A1(\dp.rf.rf[3][13] ),
    .A2(\dp.rf.rf[6][13] ),
    .A3(\dp.rf.rf[7][13] ),
    .S0(net7),
    .S1(net9),
    .X(_1282_));
 sky130_fd_sc_hd__inv_1 _4987_ (.A(\dp.rf.rf[4][13] ),
    .Y(_1283_));
 sky130_fd_sc_hd__mux2i_1 _4988_ (.A0(\dp.rf.rf[1][13] ),
    .A1(\dp.rf.rf[5][13] ),
    .S(net9),
    .Y(_1284_));
 sky130_fd_sc_hd__a221oi_1 _4989_ (.A1(_1283_),
    .A2(_0263_),
    .B1(_1284_),
    .B2(net7),
    .C1(net8),
    .Y(_1285_));
 sky130_fd_sc_hd__a211oi_1 _4990_ (.A1(net8),
    .A2(_1282_),
    .B1(_1285_),
    .C1(net197),
    .Y(_1286_));
 sky130_fd_sc_hd__a211oi_2 _4991_ (.A1(net186),
    .A2(_1281_),
    .B1(_1286_),
    .C1(_0271_),
    .Y(_1287_));
 sky130_fd_sc_hd__a21o_4 _4992_ (.A1(_1270_),
    .A2(_1278_),
    .B1(_1287_),
    .X(_3427_));
 sky130_fd_sc_hd__inv_2 _4993_ (.A(_3427_),
    .Y(_3431_));
 sky130_fd_sc_hd__o21ai_0 _4994_ (.A1(_0130_),
    .A2(_0133_),
    .B1(net4),
    .Y(_1288_));
 sky130_fd_sc_hd__nand2_2 _4995_ (.A(_1061_),
    .B(_1288_),
    .Y(_3577_));
 sky130_fd_sc_hd__mux4_1 _4996_ (.A0(\dp.rf.rf[24][12] ),
    .A1(\dp.rf.rf[25][12] ),
    .A2(\dp.rf.rf[26][12] ),
    .A3(\dp.rf.rf[27][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_1 _4997_ (.A0(\dp.rf.rf[16][12] ),
    .A1(\dp.rf.rf[17][12] ),
    .A2(\dp.rf.rf[18][12] ),
    .A3(\dp.rf.rf[19][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1290_));
 sky130_fd_sc_hd__mux4_1 _4998_ (.A0(\dp.rf.rf[28][12] ),
    .A1(\dp.rf.rf[29][12] ),
    .A2(\dp.rf.rf[30][12] ),
    .A3(\dp.rf.rf[31][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_1 _4999_ (.A0(\dp.rf.rf[20][12] ),
    .A1(\dp.rf.rf[21][12] ),
    .A2(\dp.rf.rf[22][12] ),
    .A3(\dp.rf.rf[23][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1292_));
 sky130_fd_sc_hd__mux4_1 _5000_ (.A0(_1289_),
    .A1(_1290_),
    .A2(_1291_),
    .A3(_1292_),
    .S0(_0103_),
    .S1(net15),
    .X(_1293_));
 sky130_fd_sc_hd__mux4_1 _5001_ (.A0(\dp.rf.rf[8][12] ),
    .A1(\dp.rf.rf[9][12] ),
    .A2(\dp.rf.rf[10][12] ),
    .A3(\dp.rf.rf[11][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1294_));
 sky130_fd_sc_hd__mux4_1 _5002_ (.A0(\dp.rf.rf[0][12] ),
    .A1(\dp.rf.rf[1][12] ),
    .A2(\dp.rf.rf[2][12] ),
    .A3(\dp.rf.rf[3][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1295_));
 sky130_fd_sc_hd__mux4_1 _5003_ (.A0(\dp.rf.rf[12][12] ),
    .A1(\dp.rf.rf[13][12] ),
    .A2(\dp.rf.rf[14][12] ),
    .A3(\dp.rf.rf[15][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1296_));
 sky130_fd_sc_hd__mux4_1 _5004_ (.A0(\dp.rf.rf[4][12] ),
    .A1(\dp.rf.rf[5][12] ),
    .A2(\dp.rf.rf[6][12] ),
    .A3(\dp.rf.rf[7][12] ),
    .S0(net214),
    .S1(net277),
    .X(_1297_));
 sky130_fd_sc_hd__mux4_2 _5005_ (.A0(_1294_),
    .A1(_1295_),
    .A2(_1296_),
    .A3(_1297_),
    .S0(_0103_),
    .S1(net15),
    .X(_1298_));
 sky130_fd_sc_hd__a22oi_4 _5006_ (.A1(net17),
    .A2(_1293_),
    .B1(_1298_),
    .B2(net184),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(_0132_),
    .B(_1299_),
    .Y(_1300_));
 sky130_fd_sc_hd__o21ai_0 _5008_ (.A1(_0132_),
    .A2(_3577_),
    .B1(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__xor2_1 _5009_ (.A(_0122_),
    .B(_1301_),
    .X(_3436_));
 sky130_fd_sc_hd__inv_1 _5010_ (.A(_3436_),
    .Y(_3440_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(\dp.rf.rf[22][12] ),
    .A1(\dp.rf.rf[23][12] ),
    .S(net210),
    .X(_1302_));
 sky130_fd_sc_hd__o21ai_0 _5012_ (.A1(_0148_),
    .A2(_1302_),
    .B1(net183),
    .Y(_1303_));
 sky130_fd_sc_hd__a221oi_1 _5013_ (.A1(\dp.rf.rf[19][12] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][12] ),
    .C1(net191),
    .Y(_1304_));
 sky130_fd_sc_hd__inv_1 _5014_ (.A(\dp.rf.rf[20][12] ),
    .Y(_1305_));
 sky130_fd_sc_hd__mux2i_1 _5015_ (.A0(\dp.rf.rf[17][12] ),
    .A1(\dp.rf.rf[21][12] ),
    .S(net208),
    .Y(_1306_));
 sky130_fd_sc_hd__a221oi_1 _5016_ (.A1(_1305_),
    .A2(_0263_),
    .B1(_1306_),
    .B2(net210),
    .C1(net8),
    .Y(_1307_));
 sky130_fd_sc_hd__o22ai_1 _5017_ (.A1(\dp.rf.rf[16][12] ),
    .A2(_0348_),
    .B1(_1307_),
    .B2(net197),
    .Y(_1308_));
 sky130_fd_sc_hd__o21ai_1 _5018_ (.A1(_1303_),
    .A2(_1304_),
    .B1(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__mux2_1 _5019_ (.A0(\dp.rf.rf[30][12] ),
    .A1(\dp.rf.rf[31][12] ),
    .S(net210),
    .X(_1310_));
 sky130_fd_sc_hd__o21ai_0 _5020_ (.A1(_0148_),
    .A2(_1310_),
    .B1(net183),
    .Y(_1311_));
 sky130_fd_sc_hd__a221oi_1 _5021_ (.A1(\dp.rf.rf[27][12] ),
    .A2(net210),
    .B1(net200),
    .B2(\dp.rf.rf[26][12] ),
    .C1(net191),
    .Y(_1312_));
 sky130_fd_sc_hd__mux2i_1 _5022_ (.A0(\dp.rf.rf[25][12] ),
    .A1(\dp.rf.rf[29][12] ),
    .S(net208),
    .Y(_1313_));
 sky130_fd_sc_hd__nand2_1 _5023_ (.A(net210),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__o221ai_1 _5024_ (.A1(\dp.rf.rf[28][12] ),
    .A2(_0528_),
    .B1(_0955_),
    .B2(\dp.rf.rf[24][12] ),
    .C1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__o221ai_1 _5025_ (.A1(_1311_),
    .A2(_1312_),
    .B1(_1315_),
    .B2(net8),
    .C1(net186),
    .Y(_1316_));
 sky130_fd_sc_hd__mux4_1 _5026_ (.A0(\dp.rf.rf[8][12] ),
    .A1(\dp.rf.rf[9][12] ),
    .A2(\dp.rf.rf[12][12] ),
    .A3(\dp.rf.rf[13][12] ),
    .S0(net210),
    .S1(net208),
    .X(_1317_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(net205),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__mux4_1 _5028_ (.A0(\dp.rf.rf[10][12] ),
    .A1(\dp.rf.rf[11][12] ),
    .A2(\dp.rf.rf[14][12] ),
    .A3(\dp.rf.rf[15][12] ),
    .S0(net210),
    .S1(net208),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(net8),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__a31oi_2 _5030_ (.A1(net186),
    .A2(_1318_),
    .A3(_1320_),
    .B1(_0271_),
    .Y(_1321_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(\dp.rf.rf[6][12] ),
    .A1(\dp.rf.rf[7][12] ),
    .S(net210),
    .X(_1322_));
 sky130_fd_sc_hd__o21ai_0 _5032_ (.A1(_0148_),
    .A2(_1322_),
    .B1(net183),
    .Y(_1323_));
 sky130_fd_sc_hd__a221oi_1 _5033_ (.A1(\dp.rf.rf[3][12] ),
    .A2(net210),
    .B1(net200),
    .B2(\dp.rf.rf[2][12] ),
    .C1(net189),
    .Y(_1324_));
 sky130_fd_sc_hd__inv_1 _5034_ (.A(\dp.rf.rf[4][12] ),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2i_1 _5035_ (.A0(\dp.rf.rf[1][12] ),
    .A1(\dp.rf.rf[5][12] ),
    .S(net208),
    .Y(_1326_));
 sky130_fd_sc_hd__a221oi_1 _5036_ (.A1(_1325_),
    .A2(net204),
    .B1(_1326_),
    .B2(net210),
    .C1(net8),
    .Y(_1327_));
 sky130_fd_sc_hd__o22ai_1 _5037_ (.A1(\dp.rf.rf[0][12] ),
    .A2(net180),
    .B1(_1327_),
    .B2(_0202_),
    .Y(_1328_));
 sky130_fd_sc_hd__o21ai_1 _5038_ (.A1(_1323_),
    .A2(_1324_),
    .B1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__a32o_4 _5039_ (.A1(_0232_),
    .A2(_1309_),
    .A3(_1316_),
    .B1(_1321_),
    .B2(_1329_),
    .X(_3435_));
 sky130_fd_sc_hd__clkinv_2 _5040_ (.A(_3435_),
    .Y(_3439_));
 sky130_fd_sc_hd__mux4_1 _5041_ (.A0(\dp.rf.rf[24][11] ),
    .A1(\dp.rf.rf[25][11] ),
    .A2(\dp.rf.rf[26][11] ),
    .A3(\dp.rf.rf[27][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_1 _5042_ (.A0(\dp.rf.rf[16][11] ),
    .A1(\dp.rf.rf[17][11] ),
    .A2(\dp.rf.rf[18][11] ),
    .A3(\dp.rf.rf[19][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_1 _5043_ (.A0(\dp.rf.rf[28][11] ),
    .A1(\dp.rf.rf[29][11] ),
    .A2(\dp.rf.rf[30][11] ),
    .A3(\dp.rf.rf[31][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1332_));
 sky130_fd_sc_hd__mux4_1 _5044_ (.A0(\dp.rf.rf[20][11] ),
    .A1(\dp.rf.rf[21][11] ),
    .A2(\dp.rf.rf[22][11] ),
    .A3(\dp.rf.rf[23][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1333_));
 sky130_fd_sc_hd__mux4_1 _5045_ (.A0(_1330_),
    .A1(_1331_),
    .A2(_1332_),
    .A3(_1333_),
    .S0(_0103_),
    .S1(net15),
    .X(_1334_));
 sky130_fd_sc_hd__mux4_1 _5046_ (.A0(\dp.rf.rf[8][11] ),
    .A1(\dp.rf.rf[9][11] ),
    .A2(\dp.rf.rf[10][11] ),
    .A3(\dp.rf.rf[11][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1335_));
 sky130_fd_sc_hd__mux4_1 _5047_ (.A0(\dp.rf.rf[0][11] ),
    .A1(\dp.rf.rf[1][11] ),
    .A2(\dp.rf.rf[2][11] ),
    .A3(\dp.rf.rf[3][11] ),
    .S0(net13),
    .S1(net277),
    .X(_1336_));
 sky130_fd_sc_hd__mux4_1 _5048_ (.A0(\dp.rf.rf[12][11] ),
    .A1(\dp.rf.rf[13][11] ),
    .A2(\dp.rf.rf[14][11] ),
    .A3(\dp.rf.rf[15][11] ),
    .S0(net214),
    .S1(net278),
    .X(_1337_));
 sky130_fd_sc_hd__mux4_1 _5049_ (.A0(\dp.rf.rf[4][11] ),
    .A1(\dp.rf.rf[5][11] ),
    .A2(\dp.rf.rf[6][11] ),
    .A3(\dp.rf.rf[7][11] ),
    .S0(net13),
    .S1(net278),
    .X(_1338_));
 sky130_fd_sc_hd__mux4_2 _5050_ (.A0(_1335_),
    .A1(_1336_),
    .A2(_1337_),
    .A3(_1338_),
    .S0(_0103_),
    .S1(net15),
    .X(_1339_));
 sky130_fd_sc_hd__mux2i_4 _5051_ (.A0(_1334_),
    .A1(_1339_),
    .S(_0086_),
    .Y(_1340_));
 sky130_fd_sc_hd__and2_0 _5052_ (.A(net29),
    .B(_0042_),
    .X(_1341_));
 sky130_fd_sc_hd__a22oi_2 _5053_ (.A1(net30),
    .A2(_1341_),
    .B1(_0133_),
    .B2(net13),
    .Y(_1342_));
 sky130_fd_sc_hd__o21ai_4 _5054_ (.A1(_0304_),
    .A2(_0917_),
    .B1(_1342_),
    .Y(_3573_));
 sky130_fd_sc_hd__nand2_1 _5055_ (.A(_0138_),
    .B(_3573_),
    .Y(_1343_));
 sky130_fd_sc_hd__o31ai_1 _5056_ (.A1(_0138_),
    .A2(_0401_),
    .A3(_1340_),
    .B1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__xnor2_1 _5057_ (.A(_0122_),
    .B(_1344_),
    .Y(_3444_));
 sky130_fd_sc_hd__inv_1 _5058_ (.A(_3444_),
    .Y(_3448_));
 sky130_fd_sc_hd__mux4_1 _5059_ (.A0(\dp.rf.rf[2][11] ),
    .A1(\dp.rf.rf[3][11] ),
    .A2(\dp.rf.rf[6][11] ),
    .A3(\dp.rf.rf[7][11] ),
    .S0(net210),
    .S1(net9),
    .X(_1345_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(net8),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__mux2_1 _5061_ (.A0(\dp.rf.rf[1][11] ),
    .A1(\dp.rf.rf[5][11] ),
    .S(net9),
    .X(_1347_));
 sky130_fd_sc_hd__o221ai_1 _5062_ (.A1(\dp.rf.rf[4][11] ),
    .A2(_0528_),
    .B1(_1347_),
    .B2(_0245_),
    .C1(net205),
    .Y(_1348_));
 sky130_fd_sc_hd__nand3_1 _5063_ (.A(_0493_),
    .B(_1346_),
    .C(_1348_),
    .Y(_1349_));
 sky130_fd_sc_hd__mux4_1 _5064_ (.A0(\dp.rf.rf[10][11] ),
    .A1(\dp.rf.rf[11][11] ),
    .A2(\dp.rf.rf[14][11] ),
    .A3(\dp.rf.rf[15][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1350_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(net8),
    .B(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__mux4_1 _5066_ (.A0(\dp.rf.rf[8][11] ),
    .A1(\dp.rf.rf[9][11] ),
    .A2(\dp.rf.rf[12][11] ),
    .A3(\dp.rf.rf[13][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1352_));
 sky130_fd_sc_hd__nand2_1 _5067_ (.A(net205),
    .B(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand3_1 _5068_ (.A(net186),
    .B(_1351_),
    .C(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__mux4_1 _5069_ (.A0(\dp.rf.rf[26][11] ),
    .A1(\dp.rf.rf[27][11] ),
    .A2(\dp.rf.rf[30][11] ),
    .A3(\dp.rf.rf[31][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1355_));
 sky130_fd_sc_hd__nand2_1 _5070_ (.A(net8),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__mux4_1 _5071_ (.A0(\dp.rf.rf[24][11] ),
    .A1(\dp.rf.rf[25][11] ),
    .A2(\dp.rf.rf[28][11] ),
    .A3(\dp.rf.rf[29][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1357_));
 sky130_fd_sc_hd__nand2_1 _5072_ (.A(net205),
    .B(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__a31oi_1 _5073_ (.A1(net10),
    .A2(_1356_),
    .A3(_1358_),
    .B1(_0166_),
    .Y(_1359_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(\dp.rf.rf[22][11] ),
    .A1(\dp.rf.rf[23][11] ),
    .S(net7),
    .X(_1360_));
 sky130_fd_sc_hd__o21ai_0 _5075_ (.A1(_0148_),
    .A2(_1360_),
    .B1(net183),
    .Y(_1361_));
 sky130_fd_sc_hd__a221oi_1 _5076_ (.A1(\dp.rf.rf[19][11] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[18][11] ),
    .C1(net191),
    .Y(_1362_));
 sky130_fd_sc_hd__inv_1 _5077_ (.A(\dp.rf.rf[20][11] ),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2i_1 _5078_ (.A0(\dp.rf.rf[17][11] ),
    .A1(\dp.rf.rf[21][11] ),
    .S(net9),
    .Y(_1364_));
 sky130_fd_sc_hd__a221oi_1 _5079_ (.A1(_1363_),
    .A2(_0263_),
    .B1(_1364_),
    .B2(net7),
    .C1(net8),
    .Y(_1365_));
 sky130_fd_sc_hd__o22ai_1 _5080_ (.A1(\dp.rf.rf[16][11] ),
    .A2(net180),
    .B1(_1365_),
    .B2(_0202_),
    .Y(_1366_));
 sky130_fd_sc_hd__o21ai_0 _5081_ (.A1(_1361_),
    .A2(_1362_),
    .B1(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__a32o_4 _5082_ (.A1(net193),
    .A2(_1349_),
    .A3(_1354_),
    .B1(_1359_),
    .B2(_1367_),
    .X(_3443_));
 sky130_fd_sc_hd__clkinv_2 _5083_ (.A(_3443_),
    .Y(_3447_));
 sky130_fd_sc_hd__and2_1 _5084_ (.A(net24),
    .B(_0119_),
    .X(_3569_));
 sky130_fd_sc_hd__mux4_1 _5085_ (.A0(\dp.rf.rf[24][10] ),
    .A1(\dp.rf.rf[25][10] ),
    .A2(\dp.rf.rf[26][10] ),
    .A3(\dp.rf.rf[27][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1368_));
 sky130_fd_sc_hd__mux4_1 _5086_ (.A0(\dp.rf.rf[16][10] ),
    .A1(\dp.rf.rf[17][10] ),
    .A2(\dp.rf.rf[18][10] ),
    .A3(\dp.rf.rf[19][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1369_));
 sky130_fd_sc_hd__mux4_1 _5087_ (.A0(\dp.rf.rf[28][10] ),
    .A1(\dp.rf.rf[29][10] ),
    .A2(\dp.rf.rf[30][10] ),
    .A3(\dp.rf.rf[31][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1370_));
 sky130_fd_sc_hd__mux4_1 _5088_ (.A0(\dp.rf.rf[20][10] ),
    .A1(\dp.rf.rf[21][10] ),
    .A2(\dp.rf.rf[22][10] ),
    .A3(\dp.rf.rf[23][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1371_));
 sky130_fd_sc_hd__mux4_1 _5089_ (.A0(_1368_),
    .A1(_1369_),
    .A2(_1370_),
    .A3(_1371_),
    .S0(_0103_),
    .S1(net15),
    .X(_1372_));
 sky130_fd_sc_hd__mux4_1 _5090_ (.A0(\dp.rf.rf[8][10] ),
    .A1(\dp.rf.rf[9][10] ),
    .A2(\dp.rf.rf[10][10] ),
    .A3(\dp.rf.rf[11][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1373_));
 sky130_fd_sc_hd__mux4_1 _5091_ (.A0(\dp.rf.rf[0][10] ),
    .A1(\dp.rf.rf[1][10] ),
    .A2(\dp.rf.rf[2][10] ),
    .A3(\dp.rf.rf[3][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1374_));
 sky130_fd_sc_hd__mux4_1 _5092_ (.A0(\dp.rf.rf[12][10] ),
    .A1(\dp.rf.rf[13][10] ),
    .A2(\dp.rf.rf[14][10] ),
    .A3(\dp.rf.rf[15][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1375_));
 sky130_fd_sc_hd__mux4_1 _5093_ (.A0(\dp.rf.rf[4][10] ),
    .A1(\dp.rf.rf[5][10] ),
    .A2(\dp.rf.rf[6][10] ),
    .A3(\dp.rf.rf[7][10] ),
    .S0(net214),
    .S1(net278),
    .X(_1376_));
 sky130_fd_sc_hd__mux4_1 _5094_ (.A0(_1373_),
    .A1(_1374_),
    .A2(_1375_),
    .A3(_1376_),
    .S0(_0103_),
    .S1(net15),
    .X(_1377_));
 sky130_fd_sc_hd__a22o_2 _5095_ (.A1(net17),
    .A2(_1372_),
    .B1(_1377_),
    .B2(net184),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(_3569_),
    .A1(_1378_),
    .S(_0132_),
    .X(_1379_));
 sky130_fd_sc_hd__xnor2_1 _5097_ (.A(_0122_),
    .B(_1379_),
    .Y(_3452_));
 sky130_fd_sc_hd__inv_1 _5098_ (.A(_3452_),
    .Y(_3456_));
 sky130_fd_sc_hd__mux4_1 _5099_ (.A0(\dp.rf.rf[10][10] ),
    .A1(\dp.rf.rf[11][10] ),
    .A2(\dp.rf.rf[14][10] ),
    .A3(\dp.rf.rf[15][10] ),
    .S0(net7),
    .S1(net9),
    .X(_1380_));
 sky130_fd_sc_hd__nand2_1 _5100_ (.A(net8),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__mux4_1 _5101_ (.A0(\dp.rf.rf[8][10] ),
    .A1(\dp.rf.rf[9][10] ),
    .A2(\dp.rf.rf[12][10] ),
    .A3(\dp.rf.rf[13][10] ),
    .S0(net7),
    .S1(net9),
    .X(_1382_));
 sky130_fd_sc_hd__nand2_1 _5102_ (.A(net205),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand3_1 _5103_ (.A(net186),
    .B(_1381_),
    .C(_1383_),
    .Y(_1384_));
 sky130_fd_sc_hd__mux2_1 _5104_ (.A0(\dp.rf.rf[6][10] ),
    .A1(\dp.rf.rf[7][10] ),
    .S(net7),
    .X(_1385_));
 sky130_fd_sc_hd__o21ai_0 _5105_ (.A1(_0148_),
    .A2(_1385_),
    .B1(net183),
    .Y(_1386_));
 sky130_fd_sc_hd__a221oi_1 _5106_ (.A1(\dp.rf.rf[3][10] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[2][10] ),
    .C1(net191),
    .Y(_1387_));
 sky130_fd_sc_hd__inv_1 _5107_ (.A(\dp.rf.rf[4][10] ),
    .Y(_1388_));
 sky130_fd_sc_hd__mux2i_1 _5108_ (.A0(\dp.rf.rf[1][10] ),
    .A1(\dp.rf.rf[5][10] ),
    .S(net9),
    .Y(_1389_));
 sky130_fd_sc_hd__a221oi_1 _5109_ (.A1(_1388_),
    .A2(_0263_),
    .B1(_1389_),
    .B2(net7),
    .C1(net8),
    .Y(_1390_));
 sky130_fd_sc_hd__o22ai_1 _5110_ (.A1(\dp.rf.rf[0][10] ),
    .A2(_0348_),
    .B1(_1390_),
    .B2(net197),
    .Y(_1391_));
 sky130_fd_sc_hd__o21ai_1 _5111_ (.A1(_1386_),
    .A2(_1387_),
    .B1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux4_1 _5112_ (.A0(\dp.rf.rf[26][10] ),
    .A1(\dp.rf.rf[27][10] ),
    .A2(\dp.rf.rf[30][10] ),
    .A3(\dp.rf.rf[31][10] ),
    .S0(net7),
    .S1(net9),
    .X(_1393_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(net8),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__mux4_1 _5114_ (.A0(\dp.rf.rf[24][10] ),
    .A1(\dp.rf.rf[25][10] ),
    .A2(\dp.rf.rf[28][10] ),
    .A3(\dp.rf.rf[29][10] ),
    .S0(net7),
    .S1(net9),
    .X(_1395_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(net205),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__a31oi_1 _5116_ (.A1(net10),
    .A2(_1394_),
    .A3(_1396_),
    .B1(_0166_),
    .Y(_1397_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(\dp.rf.rf[22][10] ),
    .A1(\dp.rf.rf[23][10] ),
    .S(net7),
    .X(_1398_));
 sky130_fd_sc_hd__o21ai_0 _5118_ (.A1(_0148_),
    .A2(_1398_),
    .B1(net183),
    .Y(_1399_));
 sky130_fd_sc_hd__a221oi_1 _5119_ (.A1(\dp.rf.rf[19][10] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[18][10] ),
    .C1(net191),
    .Y(_1400_));
 sky130_fd_sc_hd__inv_1 _5120_ (.A(\dp.rf.rf[20][10] ),
    .Y(_1401_));
 sky130_fd_sc_hd__mux2i_1 _5121_ (.A0(\dp.rf.rf[17][10] ),
    .A1(\dp.rf.rf[21][10] ),
    .S(net9),
    .Y(_1402_));
 sky130_fd_sc_hd__a221oi_1 _5122_ (.A1(_1401_),
    .A2(_0263_),
    .B1(_1402_),
    .B2(net7),
    .C1(net8),
    .Y(_1403_));
 sky130_fd_sc_hd__o22ai_1 _5123_ (.A1(\dp.rf.rf[16][10] ),
    .A2(_0348_),
    .B1(_1403_),
    .B2(net197),
    .Y(_1404_));
 sky130_fd_sc_hd__o21ai_0 _5124_ (.A1(_1399_),
    .A2(_1400_),
    .B1(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__a32o_4 _5125_ (.A1(net193),
    .A2(_1384_),
    .A3(_1392_),
    .B1(_1397_),
    .B2(_1405_),
    .X(_3451_));
 sky130_fd_sc_hd__clkinv_4 _5126_ (.A(_3451_),
    .Y(_3455_));
 sky130_fd_sc_hd__and2_1 _5127_ (.A(net22),
    .B(_0119_),
    .X(_3565_));
 sky130_fd_sc_hd__mux4_1 _5128_ (.A0(\dp.rf.rf[24][9] ),
    .A1(\dp.rf.rf[25][9] ),
    .A2(\dp.rf.rf[26][9] ),
    .A3(\dp.rf.rf[27][9] ),
    .S0(net13),
    .S1(net278),
    .X(_1406_));
 sky130_fd_sc_hd__mux4_1 _5129_ (.A0(\dp.rf.rf[16][9] ),
    .A1(\dp.rf.rf[17][9] ),
    .A2(\dp.rf.rf[18][9] ),
    .A3(\dp.rf.rf[19][9] ),
    .S0(net13),
    .S1(net278),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_1 _5130_ (.A0(\dp.rf.rf[28][9] ),
    .A1(\dp.rf.rf[29][9] ),
    .A2(\dp.rf.rf[30][9] ),
    .A3(\dp.rf.rf[31][9] ),
    .S0(net13),
    .S1(net278),
    .X(_1408_));
 sky130_fd_sc_hd__mux4_1 _5131_ (.A0(\dp.rf.rf[20][9] ),
    .A1(\dp.rf.rf[21][9] ),
    .A2(\dp.rf.rf[22][9] ),
    .A3(\dp.rf.rf[23][9] ),
    .S0(net13),
    .S1(net278),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_1 _5132_ (.A0(_1406_),
    .A1(_1407_),
    .A2(_1408_),
    .A3(_1409_),
    .S0(_0103_),
    .S1(net15),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_1 _5133_ (.A(net17),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux4_1 _5134_ (.A0(\dp.rf.rf[8][9] ),
    .A1(\dp.rf.rf[9][9] ),
    .A2(\dp.rf.rf[10][9] ),
    .A3(\dp.rf.rf[11][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1412_));
 sky130_fd_sc_hd__mux4_1 _5135_ (.A0(\dp.rf.rf[0][9] ),
    .A1(\dp.rf.rf[1][9] ),
    .A2(\dp.rf.rf[2][9] ),
    .A3(\dp.rf.rf[3][9] ),
    .S0(net215),
    .S1(net14),
    .X(_1413_));
 sky130_fd_sc_hd__mux4_1 _5136_ (.A0(\dp.rf.rf[12][9] ),
    .A1(\dp.rf.rf[13][9] ),
    .A2(\dp.rf.rf[14][9] ),
    .A3(\dp.rf.rf[15][9] ),
    .S0(net215),
    .S1(net14),
    .X(_1414_));
 sky130_fd_sc_hd__mux4_1 _5137_ (.A0(\dp.rf.rf[4][9] ),
    .A1(\dp.rf.rf[5][9] ),
    .A2(\dp.rf.rf[6][9] ),
    .A3(\dp.rf.rf[7][9] ),
    .S0(net215),
    .S1(net14),
    .X(_1415_));
 sky130_fd_sc_hd__mux4_2 _5138_ (.A0(_1412_),
    .A1(_1413_),
    .A2(_1414_),
    .A3(_1415_),
    .S0(_0103_),
    .S1(net15),
    .X(_1416_));
 sky130_fd_sc_hd__nand2_1 _5139_ (.A(_0086_),
    .B(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_1411_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_4 _5141_ (.A(_0311_),
    .B(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__nor2_1 _5142_ (.A(_0138_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__a21oi_1 _5143_ (.A1(_0138_),
    .A2(_3565_),
    .B1(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__xor2_1 _5144_ (.A(_0122_),
    .B(_1421_),
    .X(_3460_));
 sky130_fd_sc_hd__inv_1 _5145_ (.A(_3460_),
    .Y(_3464_));
 sky130_fd_sc_hd__mux2_1 _5146_ (.A0(\dp.rf.rf[1][9] ),
    .A1(\dp.rf.rf[5][9] ),
    .S(net208),
    .X(_1422_));
 sky130_fd_sc_hd__o22ai_1 _5147_ (.A1(\dp.rf.rf[4][9] ),
    .A2(_0528_),
    .B1(_1422_),
    .B2(_0245_),
    .Y(_1423_));
 sky130_fd_sc_hd__mux4_1 _5148_ (.A0(\dp.rf.rf[2][9] ),
    .A1(\dp.rf.rf[3][9] ),
    .A2(\dp.rf.rf[6][9] ),
    .A3(\dp.rf.rf[7][9] ),
    .S0(net211),
    .S1(net207),
    .X(_1424_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(net8),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__o211ai_2 _5150_ (.A1(net8),
    .A2(_1423_),
    .B1(_1425_),
    .C1(_0493_),
    .Y(_1426_));
 sky130_fd_sc_hd__mux4_1 _5151_ (.A0(\dp.rf.rf[10][9] ),
    .A1(\dp.rf.rf[11][9] ),
    .A2(\dp.rf.rf[14][9] ),
    .A3(\dp.rf.rf[15][9] ),
    .S0(net7),
    .S1(net9),
    .X(_1427_));
 sky130_fd_sc_hd__nand2_1 _5152_ (.A(net8),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__mux4_1 _5153_ (.A0(\dp.rf.rf[8][9] ),
    .A1(\dp.rf.rf[9][9] ),
    .A2(\dp.rf.rf[12][9] ),
    .A3(\dp.rf.rf[13][9] ),
    .S0(net7),
    .S1(net9),
    .X(_1429_));
 sky130_fd_sc_hd__nand2_1 _5154_ (.A(_0224_),
    .B(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand3_2 _5155_ (.A(net186),
    .B(_1428_),
    .C(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__mux4_1 _5156_ (.A0(\dp.rf.rf[26][9] ),
    .A1(\dp.rf.rf[27][9] ),
    .A2(\dp.rf.rf[30][9] ),
    .A3(\dp.rf.rf[31][9] ),
    .S0(net7),
    .S1(net9),
    .X(_1432_));
 sky130_fd_sc_hd__nand2_1 _5157_ (.A(net8),
    .B(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__mux4_1 _5158_ (.A0(\dp.rf.rf[24][9] ),
    .A1(\dp.rf.rf[25][9] ),
    .A2(\dp.rf.rf[28][9] ),
    .A3(\dp.rf.rf[29][9] ),
    .S0(net7),
    .S1(net9),
    .X(_1434_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(net205),
    .B(_1434_),
    .Y(_1435_));
 sky130_fd_sc_hd__a31oi_2 _5160_ (.A1(net10),
    .A2(_1433_),
    .A3(_1435_),
    .B1(_0166_),
    .Y(_1436_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(\dp.rf.rf[22][9] ),
    .A1(\dp.rf.rf[23][9] ),
    .S(net7),
    .X(_1437_));
 sky130_fd_sc_hd__o21ai_0 _5162_ (.A1(_0148_),
    .A2(_1437_),
    .B1(net183),
    .Y(_1438_));
 sky130_fd_sc_hd__a221oi_1 _5163_ (.A1(\dp.rf.rf[19][9] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[18][9] ),
    .C1(net189),
    .Y(_1439_));
 sky130_fd_sc_hd__inv_1 _5164_ (.A(\dp.rf.rf[20][9] ),
    .Y(_1440_));
 sky130_fd_sc_hd__mux2i_1 _5165_ (.A0(\dp.rf.rf[17][9] ),
    .A1(\dp.rf.rf[21][9] ),
    .S(net9),
    .Y(_1441_));
 sky130_fd_sc_hd__a221oi_1 _5166_ (.A1(_1440_),
    .A2(_0263_),
    .B1(_1441_),
    .B2(net7),
    .C1(net8),
    .Y(_1442_));
 sky130_fd_sc_hd__o22ai_1 _5167_ (.A1(\dp.rf.rf[16][9] ),
    .A2(net180),
    .B1(_1442_),
    .B2(_0202_),
    .Y(_1443_));
 sky130_fd_sc_hd__o21ai_1 _5168_ (.A1(_1438_),
    .A2(_1439_),
    .B1(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__a32oi_4 _5169_ (.A1(net193),
    .A2(_1431_),
    .A3(_1426_),
    .B1(_1436_),
    .B2(_1444_),
    .Y(_3463_));
 sky130_fd_sc_hd__mux4_1 _5170_ (.A0(\dp.rf.rf[24][8] ),
    .A1(\dp.rf.rf[25][8] ),
    .A2(\dp.rf.rf[26][8] ),
    .A3(\dp.rf.rf[27][8] ),
    .S0(net214),
    .S1(net277),
    .X(_1445_));
 sky130_fd_sc_hd__mux4_1 _5171_ (.A0(\dp.rf.rf[16][8] ),
    .A1(\dp.rf.rf[17][8] ),
    .A2(\dp.rf.rf[18][8] ),
    .A3(\dp.rf.rf[19][8] ),
    .S0(net214),
    .S1(net277),
    .X(_1446_));
 sky130_fd_sc_hd__mux4_1 _5172_ (.A0(\dp.rf.rf[28][8] ),
    .A1(\dp.rf.rf[29][8] ),
    .A2(\dp.rf.rf[30][8] ),
    .A3(\dp.rf.rf[31][8] ),
    .S0(net214),
    .S1(net277),
    .X(_1447_));
 sky130_fd_sc_hd__mux4_1 _5173_ (.A0(\dp.rf.rf[20][8] ),
    .A1(\dp.rf.rf[21][8] ),
    .A2(\dp.rf.rf[22][8] ),
    .A3(\dp.rf.rf[23][8] ),
    .S0(net214),
    .S1(net278),
    .X(_1448_));
 sky130_fd_sc_hd__mux4_1 _5174_ (.A0(_1445_),
    .A1(_1446_),
    .A2(_1447_),
    .A3(_1448_),
    .S0(_0103_),
    .S1(net15),
    .X(_1449_));
 sky130_fd_sc_hd__mux4_1 _5175_ (.A0(\dp.rf.rf[8][8] ),
    .A1(\dp.rf.rf[9][8] ),
    .A2(\dp.rf.rf[10][8] ),
    .A3(\dp.rf.rf[11][8] ),
    .S0(net214),
    .S1(net278),
    .X(_1450_));
 sky130_fd_sc_hd__mux4_1 _5176_ (.A0(\dp.rf.rf[0][8] ),
    .A1(\dp.rf.rf[1][8] ),
    .A2(\dp.rf.rf[2][8] ),
    .A3(\dp.rf.rf[3][8] ),
    .S0(net214),
    .S1(net278),
    .X(_1451_));
 sky130_fd_sc_hd__mux4_1 _5177_ (.A0(\dp.rf.rf[12][8] ),
    .A1(\dp.rf.rf[13][8] ),
    .A2(\dp.rf.rf[14][8] ),
    .A3(\dp.rf.rf[15][8] ),
    .S0(net214),
    .S1(net278),
    .X(_1452_));
 sky130_fd_sc_hd__mux4_1 _5178_ (.A0(\dp.rf.rf[4][8] ),
    .A1(\dp.rf.rf[5][8] ),
    .A2(\dp.rf.rf[6][8] ),
    .A3(\dp.rf.rf[7][8] ),
    .S0(net214),
    .S1(net278),
    .X(_1453_));
 sky130_fd_sc_hd__mux4_2 _5179_ (.A0(_1450_),
    .A1(_1451_),
    .A2(_1452_),
    .A3(_1453_),
    .S0(_0103_),
    .S1(net15),
    .X(_1454_));
 sky130_fd_sc_hd__a22oi_4 _5180_ (.A1(net17),
    .A2(_1449_),
    .B1(_1454_),
    .B2(net184),
    .Y(_1455_));
 sky130_fd_sc_hd__and2_1 _5181_ (.A(net21),
    .B(_0119_),
    .X(_3561_));
 sky130_fd_sc_hd__nor2_1 _5182_ (.A(_0132_),
    .B(_3561_),
    .Y(_1456_));
 sky130_fd_sc_hd__a21oi_1 _5183_ (.A1(_0132_),
    .A2(_1455_),
    .B1(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__xnor2_1 _5184_ (.A(_0122_),
    .B(_1457_),
    .Y(_3468_));
 sky130_fd_sc_hd__inv_1 _5185_ (.A(_3468_),
    .Y(_3472_));
 sky130_fd_sc_hd__mux4_1 _5186_ (.A0(\dp.rf.rf[24][8] ),
    .A1(\dp.rf.rf[25][8] ),
    .A2(\dp.rf.rf[28][8] ),
    .A3(\dp.rf.rf[29][8] ),
    .S0(net210),
    .S1(net208),
    .X(_1458_));
 sky130_fd_sc_hd__a21oi_1 _5187_ (.A1(net205),
    .A2(_1458_),
    .B1(net199),
    .Y(_1459_));
 sky130_fd_sc_hd__mux4_1 _5188_ (.A0(\dp.rf.rf[26][8] ),
    .A1(\dp.rf.rf[27][8] ),
    .A2(\dp.rf.rf[30][8] ),
    .A3(\dp.rf.rf[31][8] ),
    .S0(net210),
    .S1(net208),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(_0406_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__o21ai_2 _5190_ (.A1(_0166_),
    .A2(_1459_),
    .B1(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__mux4_1 _5191_ (.A0(\dp.rf.rf[18][8] ),
    .A1(\dp.rf.rf[19][8] ),
    .A2(\dp.rf.rf[22][8] ),
    .A3(\dp.rf.rf[23][8] ),
    .S0(net210),
    .S1(net208),
    .X(_1463_));
 sky130_fd_sc_hd__nand2_1 _5192_ (.A(net183),
    .B(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__inv_1 _5193_ (.A(\dp.rf.rf[20][8] ),
    .Y(_1465_));
 sky130_fd_sc_hd__mux2i_1 _5194_ (.A0(\dp.rf.rf[17][8] ),
    .A1(\dp.rf.rf[21][8] ),
    .S(net208),
    .Y(_1466_));
 sky130_fd_sc_hd__a221oi_1 _5195_ (.A1(_1465_),
    .A2(_0263_),
    .B1(_1466_),
    .B2(net210),
    .C1(net8),
    .Y(_1467_));
 sky130_fd_sc_hd__o22ai_1 _5196_ (.A1(\dp.rf.rf[16][8] ),
    .A2(_0348_),
    .B1(_1467_),
    .B2(net197),
    .Y(_1468_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(_1464_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__mux4_1 _5198_ (.A0(\dp.rf.rf[9][8] ),
    .A1(\dp.rf.rf[11][8] ),
    .A2(\dp.rf.rf[13][8] ),
    .A3(\dp.rf.rf[15][8] ),
    .S0(net8),
    .S1(net9),
    .X(_1470_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(net7),
    .B(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__mux4_1 _5200_ (.A0(\dp.rf.rf[8][8] ),
    .A1(\dp.rf.rf[10][8] ),
    .A2(\dp.rf.rf[12][8] ),
    .A3(\dp.rf.rf[14][8] ),
    .S0(net8),
    .S1(net9),
    .X(_1472_));
 sky130_fd_sc_hd__nand2_1 _5201_ (.A(_0245_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__a31oi_4 _5202_ (.A1(net186),
    .A2(_1471_),
    .A3(_1473_),
    .B1(_0271_),
    .Y(_1474_));
 sky130_fd_sc_hd__mux2_1 _5203_ (.A0(\dp.rf.rf[6][8] ),
    .A1(\dp.rf.rf[7][8] ),
    .S(net7),
    .X(_1475_));
 sky130_fd_sc_hd__o21ai_0 _5204_ (.A1(_0148_),
    .A2(_1475_),
    .B1(net183),
    .Y(_1476_));
 sky130_fd_sc_hd__a221oi_1 _5205_ (.A1(\dp.rf.rf[3][8] ),
    .A2(net7),
    .B1(_0176_),
    .B2(\dp.rf.rf[2][8] ),
    .C1(net191),
    .Y(_1477_));
 sky130_fd_sc_hd__inv_1 _5206_ (.A(\dp.rf.rf[4][8] ),
    .Y(_1478_));
 sky130_fd_sc_hd__mux2i_1 _5207_ (.A0(\dp.rf.rf[1][8] ),
    .A1(\dp.rf.rf[5][8] ),
    .S(net9),
    .Y(_1479_));
 sky130_fd_sc_hd__a221oi_1 _5208_ (.A1(_1478_),
    .A2(_0263_),
    .B1(_1479_),
    .B2(net7),
    .C1(net8),
    .Y(_1480_));
 sky130_fd_sc_hd__o22ai_1 _5209_ (.A1(\dp.rf.rf[0][8] ),
    .A2(_0348_),
    .B1(_1480_),
    .B2(net197),
    .Y(_1481_));
 sky130_fd_sc_hd__o21ai_2 _5210_ (.A1(_1476_),
    .A2(_1477_),
    .B1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hd__a22oi_4 _5211_ (.A1(_1462_),
    .A2(_1469_),
    .B1(_1474_),
    .B2(_1482_),
    .Y(_3471_));
 sky130_fd_sc_hd__mux4_1 _5212_ (.A0(\dp.rf.rf[12][7] ),
    .A1(\dp.rf.rf[13][7] ),
    .A2(\dp.rf.rf[14][7] ),
    .A3(\dp.rf.rf[15][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_1 _5213_ (.A(net16),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__mux4_1 _5214_ (.A0(\dp.rf.rf[4][7] ),
    .A1(\dp.rf.rf[5][7] ),
    .A2(\dp.rf.rf[6][7] ),
    .A3(\dp.rf.rf[7][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1485_));
 sky130_fd_sc_hd__nand2_1 _5215_ (.A(_0103_),
    .B(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand3_1 _5216_ (.A(net15),
    .B(_1484_),
    .C(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__mux4_1 _5217_ (.A0(\dp.rf.rf[8][7] ),
    .A1(\dp.rf.rf[9][7] ),
    .A2(\dp.rf.rf[10][7] ),
    .A3(\dp.rf.rf[11][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1488_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(net16),
    .B(_1488_),
    .Y(_1489_));
 sky130_fd_sc_hd__mux4_1 _5219_ (.A0(\dp.rf.rf[0][7] ),
    .A1(\dp.rf.rf[1][7] ),
    .A2(\dp.rf.rf[2][7] ),
    .A3(\dp.rf.rf[3][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _5220_ (.A(_0103_),
    .B(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__nand3_1 _5221_ (.A(_0286_),
    .B(_1489_),
    .C(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__mux4_1 _5222_ (.A0(\dp.rf.rf[28][7] ),
    .A1(\dp.rf.rf[29][7] ),
    .A2(\dp.rf.rf[30][7] ),
    .A3(\dp.rf.rf[31][7] ),
    .S0(net214),
    .S1(net277),
    .X(_1493_));
 sky130_fd_sc_hd__mux4_1 _5223_ (.A0(\dp.rf.rf[20][7] ),
    .A1(\dp.rf.rf[21][7] ),
    .A2(\dp.rf.rf[22][7] ),
    .A3(\dp.rf.rf[23][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1494_));
 sky130_fd_sc_hd__mux2i_1 _5224_ (.A0(_1493_),
    .A1(_1494_),
    .S(_0103_),
    .Y(_1495_));
 sky130_fd_sc_hd__mux4_1 _5225_ (.A0(\dp.rf.rf[24][7] ),
    .A1(\dp.rf.rf[25][7] ),
    .A2(\dp.rf.rf[26][7] ),
    .A3(\dp.rf.rf[27][7] ),
    .S0(net214),
    .S1(net277),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _5226_ (.A(net16),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux4_1 _5227_ (.A0(\dp.rf.rf[16][7] ),
    .A1(\dp.rf.rf[17][7] ),
    .A2(\dp.rf.rf[18][7] ),
    .A3(\dp.rf.rf[19][7] ),
    .S0(net13),
    .S1(net277),
    .X(_1498_));
 sky130_fd_sc_hd__nand2_1 _5228_ (.A(_0103_),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__and3_1 _5229_ (.A(_0286_),
    .B(_1497_),
    .C(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__a21oi_1 _5230_ (.A1(net15),
    .A2(_1495_),
    .B1(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__a32oi_4 _5231_ (.A1(net184),
    .A2(_1487_),
    .A3(_1492_),
    .B1(_1501_),
    .B2(net17),
    .Y(_1502_));
 sky130_fd_sc_hd__inv_1 _5232_ (.A(_1502_),
    .Y(net162));
 sky130_fd_sc_hd__and2_1 _5233_ (.A(net20),
    .B(_0119_),
    .X(_3557_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_0138_),
    .B(_3557_),
    .Y(_1503_));
 sky130_fd_sc_hd__o21ai_0 _5235_ (.A1(_0138_),
    .A2(_1502_),
    .B1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__xnor2_1 _5236_ (.A(_0122_),
    .B(_1504_),
    .Y(_3476_));
 sky130_fd_sc_hd__inv_1 _5237_ (.A(_3476_),
    .Y(_3480_));
 sky130_fd_sc_hd__mux4_1 _5238_ (.A0(\dp.rf.rf[8][7] ),
    .A1(\dp.rf.rf[9][7] ),
    .A2(\dp.rf.rf[12][7] ),
    .A3(\dp.rf.rf[13][7] ),
    .S0(net210),
    .S1(net208),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(net205),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__mux4_1 _5240_ (.A0(\dp.rf.rf[10][7] ),
    .A1(\dp.rf.rf[11][7] ),
    .A2(\dp.rf.rf[14][7] ),
    .A3(\dp.rf.rf[15][7] ),
    .S0(net210),
    .S1(net208),
    .X(_1507_));
 sky130_fd_sc_hd__a21oi_1 _5241_ (.A1(net183),
    .A2(_1507_),
    .B1(_0192_),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_1506_),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(\dp.rf.rf[6][7] ),
    .A1(\dp.rf.rf[7][7] ),
    .S(net210),
    .X(_1510_));
 sky130_fd_sc_hd__o21ai_0 _5244_ (.A1(_0148_),
    .A2(_1510_),
    .B1(net183),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _5245_ (.A1(\dp.rf.rf[3][7] ),
    .A2(net209),
    .B1(net200),
    .B2(\dp.rf.rf[2][7] ),
    .C1(net189),
    .Y(_1512_));
 sky130_fd_sc_hd__inv_1 _5246_ (.A(\dp.rf.rf[4][7] ),
    .Y(_1513_));
 sky130_fd_sc_hd__mux2i_1 _5247_ (.A0(\dp.rf.rf[1][7] ),
    .A1(\dp.rf.rf[5][7] ),
    .S(net208),
    .Y(_1514_));
 sky130_fd_sc_hd__a221oi_1 _5248_ (.A1(_1513_),
    .A2(net204),
    .B1(_1514_),
    .B2(net210),
    .C1(net8),
    .Y(_1515_));
 sky130_fd_sc_hd__o22ai_1 _5249_ (.A1(\dp.rf.rf[0][7] ),
    .A2(net180),
    .B1(_1515_),
    .B2(_0202_),
    .Y(_1516_));
 sky130_fd_sc_hd__o21ai_2 _5250_ (.A1(_1511_),
    .A2(_1512_),
    .B1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__mux4_1 _5251_ (.A0(\dp.rf.rf[24][7] ),
    .A1(\dp.rf.rf[25][7] ),
    .A2(\dp.rf.rf[28][7] ),
    .A3(\dp.rf.rf[29][7] ),
    .S0(net210),
    .S1(net208),
    .X(_1518_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(net205),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__mux4_1 _5253_ (.A0(\dp.rf.rf[26][7] ),
    .A1(\dp.rf.rf[27][7] ),
    .A2(\dp.rf.rf[30][7] ),
    .A3(\dp.rf.rf[31][7] ),
    .S0(net210),
    .S1(net208),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _5254_ (.A(net8),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__a31oi_2 _5255_ (.A1(net10),
    .A2(_1519_),
    .A3(_1521_),
    .B1(_0166_),
    .Y(_1522_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(\dp.rf.rf[22][7] ),
    .A1(\dp.rf.rf[23][7] ),
    .S(net210),
    .X(_1523_));
 sky130_fd_sc_hd__o21ai_0 _5257_ (.A1(_0148_),
    .A2(_1523_),
    .B1(net183),
    .Y(_1524_));
 sky130_fd_sc_hd__a221oi_1 _5258_ (.A1(\dp.rf.rf[19][7] ),
    .A2(net210),
    .B1(net200),
    .B2(\dp.rf.rf[18][7] ),
    .C1(net189),
    .Y(_1525_));
 sky130_fd_sc_hd__inv_1 _5259_ (.A(\dp.rf.rf[20][7] ),
    .Y(_1526_));
 sky130_fd_sc_hd__mux2i_1 _5260_ (.A0(\dp.rf.rf[17][7] ),
    .A1(\dp.rf.rf[21][7] ),
    .S(net208),
    .Y(_1527_));
 sky130_fd_sc_hd__a221oi_1 _5261_ (.A1(_1526_),
    .A2(net204),
    .B1(_1527_),
    .B2(net210),
    .C1(net8),
    .Y(_1528_));
 sky130_fd_sc_hd__o22ai_1 _5262_ (.A1(\dp.rf.rf[16][7] ),
    .A2(net180),
    .B1(_1528_),
    .B2(_0202_),
    .Y(_1529_));
 sky130_fd_sc_hd__o21ai_1 _5263_ (.A1(_1524_),
    .A2(_1525_),
    .B1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hd__a32oi_4 _5264_ (.A1(_1509_),
    .A2(net193),
    .A3(_1517_),
    .B1(_1522_),
    .B2(_1530_),
    .Y(_3479_));
 sky130_fd_sc_hd__mux4_1 _5265_ (.A0(\dp.rf.rf[24][6] ),
    .A1(\dp.rf.rf[25][6] ),
    .A2(\dp.rf.rf[26][6] ),
    .A3(\dp.rf.rf[27][6] ),
    .S0(net213),
    .S1(net278),
    .X(_1531_));
 sky130_fd_sc_hd__mux4_1 _5266_ (.A0(\dp.rf.rf[16][6] ),
    .A1(\dp.rf.rf[17][6] ),
    .A2(\dp.rf.rf[18][6] ),
    .A3(\dp.rf.rf[19][6] ),
    .S0(net213),
    .S1(net278),
    .X(_1532_));
 sky130_fd_sc_hd__mux4_1 _5267_ (.A0(\dp.rf.rf[28][6] ),
    .A1(\dp.rf.rf[29][6] ),
    .A2(\dp.rf.rf[30][6] ),
    .A3(\dp.rf.rf[31][6] ),
    .S0(net213),
    .S1(net278),
    .X(_1533_));
 sky130_fd_sc_hd__mux4_1 _5268_ (.A0(\dp.rf.rf[20][6] ),
    .A1(\dp.rf.rf[21][6] ),
    .A2(\dp.rf.rf[22][6] ),
    .A3(\dp.rf.rf[23][6] ),
    .S0(net213),
    .S1(net278),
    .X(_1534_));
 sky130_fd_sc_hd__mux4_1 _5269_ (.A0(_1531_),
    .A1(_1532_),
    .A2(_1533_),
    .A3(_1534_),
    .S0(_0103_),
    .S1(net15),
    .X(_1535_));
 sky130_fd_sc_hd__mux4_1 _5270_ (.A0(\dp.rf.rf[8][6] ),
    .A1(\dp.rf.rf[9][6] ),
    .A2(\dp.rf.rf[10][6] ),
    .A3(\dp.rf.rf[11][6] ),
    .S0(net215),
    .S1(net14),
    .X(_1536_));
 sky130_fd_sc_hd__mux4_1 _5271_ (.A0(\dp.rf.rf[0][6] ),
    .A1(\dp.rf.rf[1][6] ),
    .A2(\dp.rf.rf[2][6] ),
    .A3(\dp.rf.rf[3][6] ),
    .S0(net215),
    .S1(net14),
    .X(_1537_));
 sky130_fd_sc_hd__mux4_1 _5272_ (.A0(\dp.rf.rf[12][6] ),
    .A1(\dp.rf.rf[13][6] ),
    .A2(\dp.rf.rf[14][6] ),
    .A3(\dp.rf.rf[15][6] ),
    .S0(net215),
    .S1(net14),
    .X(_1538_));
 sky130_fd_sc_hd__mux4_1 _5273_ (.A0(\dp.rf.rf[4][6] ),
    .A1(\dp.rf.rf[5][6] ),
    .A2(\dp.rf.rf[6][6] ),
    .A3(\dp.rf.rf[7][6] ),
    .S0(net215),
    .S1(net14),
    .X(_1539_));
 sky130_fd_sc_hd__mux4_1 _5274_ (.A0(_1536_),
    .A1(_1537_),
    .A2(_1538_),
    .A3(_1539_),
    .S0(_0103_),
    .S1(net15),
    .X(_1540_));
 sky130_fd_sc_hd__a22o_4 _5275_ (.A1(net17),
    .A2(_1535_),
    .B1(_1540_),
    .B2(net184),
    .X(net161));
 sky130_fd_sc_hd__and2_1 _5276_ (.A(net19),
    .B(_0119_),
    .X(_3553_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(net161),
    .A1(_3553_),
    .S(_0138_),
    .X(_1541_));
 sky130_fd_sc_hd__xnor2_1 _5278_ (.A(_0122_),
    .B(_1541_),
    .Y(_3484_));
 sky130_fd_sc_hd__inv_1 _5279_ (.A(_3484_),
    .Y(_3488_));
 sky130_fd_sc_hd__mux4_1 _5280_ (.A0(\dp.rf.rf[10][6] ),
    .A1(\dp.rf.rf[11][6] ),
    .A2(\dp.rf.rf[14][6] ),
    .A3(\dp.rf.rf[15][6] ),
    .S0(net211),
    .S1(net207),
    .X(_1542_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(net8),
    .B(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__mux4_1 _5282_ (.A0(\dp.rf.rf[8][6] ),
    .A1(\dp.rf.rf[9][6] ),
    .A2(\dp.rf.rf[12][6] ),
    .A3(\dp.rf.rf[13][6] ),
    .S0(net211),
    .S1(net207),
    .X(_1544_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_0224_),
    .B(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand3_2 _5284_ (.A(net185),
    .B(_1543_),
    .C(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(\dp.rf.rf[6][6] ),
    .A1(\dp.rf.rf[7][6] ),
    .S(net211),
    .X(_1547_));
 sky130_fd_sc_hd__o21ai_0 _5286_ (.A1(_0148_),
    .A2(_1547_),
    .B1(_0337_),
    .Y(_1548_));
 sky130_fd_sc_hd__a221oi_1 _5287_ (.A1(\dp.rf.rf[3][6] ),
    .A2(net211),
    .B1(net200),
    .B2(\dp.rf.rf[2][6] ),
    .C1(net189),
    .Y(_1549_));
 sky130_fd_sc_hd__inv_1 _5288_ (.A(\dp.rf.rf[4][6] ),
    .Y(_1550_));
 sky130_fd_sc_hd__mux2i_1 _5289_ (.A0(\dp.rf.rf[1][6] ),
    .A1(\dp.rf.rf[5][6] ),
    .S(net207),
    .Y(_1551_));
 sky130_fd_sc_hd__a221oi_1 _5290_ (.A1(_1550_),
    .A2(net204),
    .B1(_1551_),
    .B2(net211),
    .C1(net8),
    .Y(_1552_));
 sky130_fd_sc_hd__o22ai_1 _5291_ (.A1(\dp.rf.rf[0][6] ),
    .A2(net180),
    .B1(_1552_),
    .B2(_0202_),
    .Y(_1553_));
 sky130_fd_sc_hd__o21ai_2 _5292_ (.A1(_1548_),
    .A2(_1549_),
    .B1(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__mux4_1 _5293_ (.A0(\dp.rf.rf[26][6] ),
    .A1(\dp.rf.rf[27][6] ),
    .A2(\dp.rf.rf[30][6] ),
    .A3(\dp.rf.rf[31][6] ),
    .S0(net7),
    .S1(net208),
    .X(_1555_));
 sky130_fd_sc_hd__nand2_1 _5294_ (.A(net8),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__mux4_1 _5295_ (.A0(\dp.rf.rf[24][6] ),
    .A1(\dp.rf.rf[25][6] ),
    .A2(\dp.rf.rf[28][6] ),
    .A3(\dp.rf.rf[29][6] ),
    .S0(net7),
    .S1(net208),
    .X(_1557_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_0224_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__a31oi_2 _5297_ (.A1(net10),
    .A2(_1556_),
    .A3(_1558_),
    .B1(_0166_),
    .Y(_1559_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(\dp.rf.rf[22][6] ),
    .A1(\dp.rf.rf[23][6] ),
    .S(net7),
    .X(_1560_));
 sky130_fd_sc_hd__o21ai_0 _5299_ (.A1(_0148_),
    .A2(_1560_),
    .B1(_0337_),
    .Y(_1561_));
 sky130_fd_sc_hd__a221oi_1 _5300_ (.A1(\dp.rf.rf[19][6] ),
    .A2(net7),
    .B1(net200),
    .B2(\dp.rf.rf[18][6] ),
    .C1(net189),
    .Y(_1562_));
 sky130_fd_sc_hd__inv_1 _5301_ (.A(\dp.rf.rf[20][6] ),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2i_1 _5302_ (.A0(\dp.rf.rf[17][6] ),
    .A1(\dp.rf.rf[21][6] ),
    .S(net206),
    .Y(_1564_));
 sky130_fd_sc_hd__a221oi_1 _5303_ (.A1(_1563_),
    .A2(net204),
    .B1(_1564_),
    .B2(net7),
    .C1(net8),
    .Y(_1565_));
 sky130_fd_sc_hd__o22ai_1 _5304_ (.A1(\dp.rf.rf[16][6] ),
    .A2(net180),
    .B1(_1565_),
    .B2(_0202_),
    .Y(_1566_));
 sky130_fd_sc_hd__o21ai_1 _5305_ (.A1(_1561_),
    .A2(_1562_),
    .B1(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__a32oi_4 _5306_ (.A1(_1546_),
    .A2(net193),
    .A3(_1554_),
    .B1(_1567_),
    .B2(_1559_),
    .Y(_3487_));
 sky130_fd_sc_hd__mux4_1 _5307_ (.A0(\dp.rf.rf[24][5] ),
    .A1(\dp.rf.rf[25][5] ),
    .A2(\dp.rf.rf[26][5] ),
    .A3(\dp.rf.rf[27][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_1 _5308_ (.A0(\dp.rf.rf[16][5] ),
    .A1(\dp.rf.rf[17][5] ),
    .A2(\dp.rf.rf[18][5] ),
    .A3(\dp.rf.rf[19][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_1 _5309_ (.A0(\dp.rf.rf[28][5] ),
    .A1(\dp.rf.rf[29][5] ),
    .A2(\dp.rf.rf[30][5] ),
    .A3(\dp.rf.rf[31][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1570_));
 sky130_fd_sc_hd__mux4_1 _5310_ (.A0(\dp.rf.rf[20][5] ),
    .A1(\dp.rf.rf[21][5] ),
    .A2(\dp.rf.rf[22][5] ),
    .A3(\dp.rf.rf[23][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1571_));
 sky130_fd_sc_hd__mux4_2 _5311_ (.A0(_1568_),
    .A1(_1569_),
    .A2(_1570_),
    .A3(_1571_),
    .S0(_0103_),
    .S1(net15),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_1 _5312_ (.A0(\dp.rf.rf[8][5] ),
    .A1(\dp.rf.rf[9][5] ),
    .A2(\dp.rf.rf[10][5] ),
    .A3(\dp.rf.rf[11][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1573_));
 sky130_fd_sc_hd__mux4_1 _5313_ (.A0(\dp.rf.rf[0][5] ),
    .A1(\dp.rf.rf[1][5] ),
    .A2(\dp.rf.rf[2][5] ),
    .A3(\dp.rf.rf[3][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1574_));
 sky130_fd_sc_hd__mux4_1 _5314_ (.A0(\dp.rf.rf[12][5] ),
    .A1(\dp.rf.rf[13][5] ),
    .A2(\dp.rf.rf[14][5] ),
    .A3(\dp.rf.rf[15][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1575_));
 sky130_fd_sc_hd__mux4_1 _5315_ (.A0(\dp.rf.rf[4][5] ),
    .A1(\dp.rf.rf[5][5] ),
    .A2(\dp.rf.rf[6][5] ),
    .A3(\dp.rf.rf[7][5] ),
    .S0(net214),
    .S1(net277),
    .X(_1576_));
 sky130_fd_sc_hd__mux4_1 _5316_ (.A0(_1573_),
    .A1(_1574_),
    .A2(_1575_),
    .A3(_1576_),
    .S0(_0103_),
    .S1(net15),
    .X(_1577_));
 sky130_fd_sc_hd__mux2i_4 _5317_ (.A0(_1572_),
    .A1(_1577_),
    .S(_0086_),
    .Y(_1578_));
 sky130_fd_sc_hd__nor2_2 _5318_ (.A(_0401_),
    .B(_1578_),
    .Y(net160));
 sky130_fd_sc_hd__and2_1 _5319_ (.A(net18),
    .B(_0119_),
    .X(_3549_));
 sky130_fd_sc_hd__nor3_1 _5320_ (.A(_0138_),
    .B(_0401_),
    .C(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__a21oi_1 _5321_ (.A1(_0138_),
    .A2(_3549_),
    .B1(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__xor2_1 _5322_ (.A(_0122_),
    .B(_1580_),
    .X(_3492_));
 sky130_fd_sc_hd__inv_1 _5323_ (.A(_3492_),
    .Y(_3496_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(\dp.rf.rf[26][5] ),
    .A1(\dp.rf.rf[27][5] ),
    .S(net7),
    .X(_1581_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(\dp.rf.rf[30][5] ),
    .A1(\dp.rf.rf[31][5] ),
    .S(net7),
    .X(_1582_));
 sky130_fd_sc_hd__o221ai_1 _5326_ (.A1(net191),
    .A2(_1581_),
    .B1(_1582_),
    .B2(_0148_),
    .C1(net8),
    .Y(_1583_));
 sky130_fd_sc_hd__mux4_1 _5327_ (.A0(\dp.rf.rf[24][5] ),
    .A1(\dp.rf.rf[25][5] ),
    .A2(\dp.rf.rf[28][5] ),
    .A3(\dp.rf.rf[29][5] ),
    .S0(net7),
    .S1(net9),
    .X(_1584_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(net205),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__nand3_1 _5329_ (.A(net186),
    .B(_1583_),
    .C(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__nor2b_1 _5330_ (.A(net7),
    .B_N(\dp.rf.rf[22][5] ),
    .Y(_1587_));
 sky130_fd_sc_hd__a211oi_1 _5331_ (.A1(\dp.rf.rf[23][5] ),
    .A2(net7),
    .B1(_0148_),
    .C1(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__a221oi_1 _5332_ (.A1(\dp.rf.rf[19][5] ),
    .A2(net7),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][5] ),
    .C1(net191),
    .Y(_1589_));
 sky130_fd_sc_hd__inv_1 _5333_ (.A(\dp.rf.rf[20][5] ),
    .Y(_1590_));
 sky130_fd_sc_hd__mux2i_1 _5334_ (.A0(\dp.rf.rf[17][5] ),
    .A1(\dp.rf.rf[21][5] ),
    .S(net208),
    .Y(_1591_));
 sky130_fd_sc_hd__a221oi_1 _5335_ (.A1(_1590_),
    .A2(_0263_),
    .B1(_1591_),
    .B2(net7),
    .C1(net8),
    .Y(_1592_));
 sky130_fd_sc_hd__o22ai_1 _5336_ (.A1(\dp.rf.rf[16][5] ),
    .A2(_0348_),
    .B1(_1592_),
    .B2(net197),
    .Y(_1593_));
 sky130_fd_sc_hd__o31ai_2 _5337_ (.A1(net192),
    .A2(_1588_),
    .A3(_1589_),
    .B1(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__mux4_1 _5338_ (.A0(\dp.rf.rf[10][5] ),
    .A1(\dp.rf.rf[11][5] ),
    .A2(\dp.rf.rf[14][5] ),
    .A3(\dp.rf.rf[15][5] ),
    .S0(net210),
    .S1(net208),
    .X(_1595_));
 sky130_fd_sc_hd__mux4_1 _5339_ (.A0(\dp.rf.rf[8][5] ),
    .A1(\dp.rf.rf[9][5] ),
    .A2(\dp.rf.rf[12][5] ),
    .A3(\dp.rf.rf[13][5] ),
    .S0(net210),
    .S1(net208),
    .X(_1596_));
 sky130_fd_sc_hd__mux2i_1 _5340_ (.A0(_1595_),
    .A1(_1596_),
    .S(net205),
    .Y(_1597_));
 sky130_fd_sc_hd__mux4_1 _5341_ (.A0(\dp.rf.rf[2][5] ),
    .A1(\dp.rf.rf[3][5] ),
    .A2(\dp.rf.rf[6][5] ),
    .A3(\dp.rf.rf[7][5] ),
    .S0(net210),
    .S1(net208),
    .X(_1598_));
 sky130_fd_sc_hd__inv_1 _5342_ (.A(\dp.rf.rf[4][5] ),
    .Y(_1599_));
 sky130_fd_sc_hd__mux2i_1 _5343_ (.A0(\dp.rf.rf[1][5] ),
    .A1(\dp.rf.rf[5][5] ),
    .S(net208),
    .Y(_1600_));
 sky130_fd_sc_hd__a221oi_1 _5344_ (.A1(_1599_),
    .A2(_0263_),
    .B1(_1600_),
    .B2(net210),
    .C1(net8),
    .Y(_1601_));
 sky130_fd_sc_hd__a211oi_1 _5345_ (.A1(net8),
    .A2(_1598_),
    .B1(_1601_),
    .C1(net197),
    .Y(_1602_));
 sky130_fd_sc_hd__a211oi_2 _5346_ (.A1(net186),
    .A2(_1597_),
    .B1(_1602_),
    .C1(_0271_),
    .Y(_1603_));
 sky130_fd_sc_hd__a31oi_4 _5347_ (.A1(_0232_),
    .A2(_1586_),
    .A3(_1594_),
    .B1(_1603_),
    .Y(_3495_));
 sky130_fd_sc_hd__nor2_2 _5348_ (.A(_0042_),
    .B(_0130_),
    .Y(_1604_));
 sky130_fd_sc_hd__a22oi_4 _5349_ (.A1(net3),
    .A2(_0042_),
    .B1(_1604_),
    .B2(net17),
    .Y(_1605_));
 sky130_fd_sc_hd__inv_1 _5350_ (.A(_1605_),
    .Y(_3545_));
 sky130_fd_sc_hd__mux4_1 _5351_ (.A0(\dp.rf.rf[4][4] ),
    .A1(\dp.rf.rf[5][4] ),
    .A2(\dp.rf.rf[6][4] ),
    .A3(\dp.rf.rf[7][4] ),
    .S0(net215),
    .S1(net14),
    .X(_1606_));
 sky130_fd_sc_hd__mux4_1 _5352_ (.A0(\dp.rf.rf[0][4] ),
    .A1(\dp.rf.rf[1][4] ),
    .A2(\dp.rf.rf[2][4] ),
    .A3(\dp.rf.rf[3][4] ),
    .S0(net215),
    .S1(net14),
    .X(_1607_));
 sky130_fd_sc_hd__mux2i_2 _5353_ (.A0(_1606_),
    .A1(_1607_),
    .S(_0286_),
    .Y(_1608_));
 sky130_fd_sc_hd__mux4_1 _5354_ (.A0(\dp.rf.rf[28][4] ),
    .A1(\dp.rf.rf[29][4] ),
    .A2(\dp.rf.rf[30][4] ),
    .A3(\dp.rf.rf[31][4] ),
    .S0(net213),
    .S1(net278),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_1 _5355_ (.A0(\dp.rf.rf[20][4] ),
    .A1(\dp.rf.rf[21][4] ),
    .A2(\dp.rf.rf[22][4] ),
    .A3(\dp.rf.rf[23][4] ),
    .S0(net213),
    .S1(net278),
    .X(_1610_));
 sky130_fd_sc_hd__mux4_1 _5356_ (.A0(\dp.rf.rf[24][4] ),
    .A1(\dp.rf.rf[25][4] ),
    .A2(\dp.rf.rf[26][4] ),
    .A3(\dp.rf.rf[27][4] ),
    .S0(net213),
    .S1(net278),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_1 _5357_ (.A0(\dp.rf.rf[16][4] ),
    .A1(\dp.rf.rf[17][4] ),
    .A2(\dp.rf.rf[18][4] ),
    .A3(\dp.rf.rf[19][4] ),
    .S0(net213),
    .S1(net278),
    .X(_1612_));
 sky130_fd_sc_hd__mux4_1 _5358_ (.A0(_1609_),
    .A1(_1610_),
    .A2(_1611_),
    .A3(_1612_),
    .S0(_0103_),
    .S1(_0286_),
    .X(_1613_));
 sky130_fd_sc_hd__nor2_1 _5359_ (.A(_0086_),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__mux4_1 _5360_ (.A0(\dp.rf.rf[12][4] ),
    .A1(\dp.rf.rf[13][4] ),
    .A2(\dp.rf.rf[14][4] ),
    .A3(\dp.rf.rf[15][4] ),
    .S0(net215),
    .S1(net14),
    .X(_1615_));
 sky130_fd_sc_hd__mux4_1 _5361_ (.A0(\dp.rf.rf[8][4] ),
    .A1(\dp.rf.rf[9][4] ),
    .A2(\dp.rf.rf[10][4] ),
    .A3(\dp.rf.rf[11][4] ),
    .S0(net215),
    .S1(net14),
    .X(_1616_));
 sky130_fd_sc_hd__o22ai_1 _5362_ (.A1(_0449_),
    .A2(_1615_),
    .B1(_1616_),
    .B2(_0448_),
    .Y(_1617_));
 sky130_fd_sc_hd__a2111o_4 _5363_ (.A1(_0394_),
    .A2(_1608_),
    .B1(_1617_),
    .C1(_0401_),
    .D1(_1614_),
    .X(_1618_));
 sky130_fd_sc_hd__inv_1 _5364_ (.A(net428),
    .Y(net159));
 sky130_fd_sc_hd__mux2i_4 _5365_ (.A0(_1605_),
    .A1(_1618_),
    .S(net178),
    .Y(_1619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__xnor2_1 _5368_ (.A(_0122_),
    .B(_1619_),
    .Y(_3500_));
 sky130_fd_sc_hd__inv_1 _5369_ (.A(_3500_),
    .Y(_3504_));
 sky130_fd_sc_hd__mux4_1 _5370_ (.A0(\dp.rf.rf[9][4] ),
    .A1(\dp.rf.rf[11][4] ),
    .A2(\dp.rf.rf[13][4] ),
    .A3(\dp.rf.rf[15][4] ),
    .S0(net8),
    .S1(net207),
    .X(_1622_));
 sky130_fd_sc_hd__nand2_1 _5371_ (.A(net211),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__mux4_1 _5372_ (.A0(\dp.rf.rf[8][4] ),
    .A1(\dp.rf.rf[10][4] ),
    .A2(\dp.rf.rf[12][4] ),
    .A3(\dp.rf.rf[14][4] ),
    .S0(net8),
    .S1(net207),
    .X(_1624_));
 sky130_fd_sc_hd__nand2_1 _5373_ (.A(_0245_),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand3_1 _5374_ (.A(net185),
    .B(_1623_),
    .C(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(\dp.rf.rf[1][4] ),
    .A1(\dp.rf.rf[5][4] ),
    .S(net207),
    .X(_1627_));
 sky130_fd_sc_hd__o22ai_1 _5376_ (.A1(\dp.rf.rf[4][4] ),
    .A2(_0528_),
    .B1(_1627_),
    .B2(_0245_),
    .Y(_1628_));
 sky130_fd_sc_hd__mux4_1 _5377_ (.A0(\dp.rf.rf[2][4] ),
    .A1(\dp.rf.rf[3][4] ),
    .A2(\dp.rf.rf[6][4] ),
    .A3(\dp.rf.rf[7][4] ),
    .S0(net211),
    .S1(net207),
    .X(_1629_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(net8),
    .B(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__o211ai_2 _5379_ (.A1(net8),
    .A2(_1628_),
    .B1(_1630_),
    .C1(_0493_),
    .Y(_1631_));
 sky130_fd_sc_hd__mux4_1 _5380_ (.A0(\dp.rf.rf[24][4] ),
    .A1(\dp.rf.rf[25][4] ),
    .A2(\dp.rf.rf[28][4] ),
    .A3(\dp.rf.rf[29][4] ),
    .S0(net7),
    .S1(net206),
    .X(_1632_));
 sky130_fd_sc_hd__nand2_1 _5381_ (.A(net205),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__mux4_1 _5382_ (.A0(\dp.rf.rf[26][4] ),
    .A1(\dp.rf.rf[27][4] ),
    .A2(\dp.rf.rf[30][4] ),
    .A3(\dp.rf.rf[31][4] ),
    .S0(net7),
    .S1(net206),
    .X(_1634_));
 sky130_fd_sc_hd__nand2_1 _5383_ (.A(net8),
    .B(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__nand3_1 _5384_ (.A(net185),
    .B(_1633_),
    .C(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__mux2i_1 _5385_ (.A0(\dp.rf.rf[16][4] ),
    .A1(\dp.rf.rf[20][4] ),
    .S(net206),
    .Y(_1637_));
 sky130_fd_sc_hd__mux2i_1 _5386_ (.A0(\dp.rf.rf[17][4] ),
    .A1(\dp.rf.rf[21][4] ),
    .S(net206),
    .Y(_1638_));
 sky130_fd_sc_hd__o221ai_1 _5387_ (.A1(_0170_),
    .A2(_1637_),
    .B1(_1638_),
    .B2(_0415_),
    .C1(_0145_),
    .Y(_1639_));
 sky130_fd_sc_hd__mux4_1 _5388_ (.A0(\dp.rf.rf[18][4] ),
    .A1(\dp.rf.rf[19][4] ),
    .A2(\dp.rf.rf[22][4] ),
    .A3(\dp.rf.rf[23][4] ),
    .S0(net7),
    .S1(net206),
    .X(_1640_));
 sky130_fd_sc_hd__a22o_1 _5389_ (.A1(net188),
    .A2(_1639_),
    .B1(_1640_),
    .B2(_0406_),
    .X(_1641_));
 sky130_fd_sc_hd__a32o_4 _5390_ (.A1(_0209_),
    .A2(_1626_),
    .A3(_1631_),
    .B1(_1636_),
    .B2(_1641_),
    .X(_3499_));
 sky130_fd_sc_hd__clkinv_2 _5391_ (.A(_3499_),
    .Y(_3503_));
 sky130_fd_sc_hd__a22o_2 _5392_ (.A1(net2),
    .A2(_0042_),
    .B1(_1604_),
    .B2(net16),
    .X(_3539_));
 sky130_fd_sc_hd__mux4_1 _5393_ (.A0(\dp.rf.rf[24][3] ),
    .A1(\dp.rf.rf[25][3] ),
    .A2(\dp.rf.rf[26][3] ),
    .A3(\dp.rf.rf[27][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1642_));
 sky130_fd_sc_hd__mux4_1 _5394_ (.A0(\dp.rf.rf[16][3] ),
    .A1(\dp.rf.rf[17][3] ),
    .A2(\dp.rf.rf[18][3] ),
    .A3(\dp.rf.rf[19][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1643_));
 sky130_fd_sc_hd__mux4_1 _5395_ (.A0(\dp.rf.rf[28][3] ),
    .A1(\dp.rf.rf[29][3] ),
    .A2(\dp.rf.rf[30][3] ),
    .A3(\dp.rf.rf[31][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1644_));
 sky130_fd_sc_hd__mux4_1 _5396_ (.A0(\dp.rf.rf[20][3] ),
    .A1(\dp.rf.rf[21][3] ),
    .A2(\dp.rf.rf[22][3] ),
    .A3(\dp.rf.rf[23][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1645_));
 sky130_fd_sc_hd__mux4_1 _5397_ (.A0(_1642_),
    .A1(_1643_),
    .A2(_1644_),
    .A3(_1645_),
    .S0(_0103_),
    .S1(net15),
    .X(_1646_));
 sky130_fd_sc_hd__mux4_1 _5398_ (.A0(\dp.rf.rf[8][3] ),
    .A1(\dp.rf.rf[9][3] ),
    .A2(\dp.rf.rf[10][3] ),
    .A3(\dp.rf.rf[11][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1647_));
 sky130_fd_sc_hd__mux4_1 _5399_ (.A0(\dp.rf.rf[0][3] ),
    .A1(\dp.rf.rf[1][3] ),
    .A2(\dp.rf.rf[2][3] ),
    .A3(\dp.rf.rf[3][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1648_));
 sky130_fd_sc_hd__mux4_1 _5400_ (.A0(\dp.rf.rf[12][3] ),
    .A1(\dp.rf.rf[13][3] ),
    .A2(\dp.rf.rf[14][3] ),
    .A3(\dp.rf.rf[15][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1649_));
 sky130_fd_sc_hd__mux4_1 _5401_ (.A0(\dp.rf.rf[4][3] ),
    .A1(\dp.rf.rf[5][3] ),
    .A2(\dp.rf.rf[6][3] ),
    .A3(\dp.rf.rf[7][3] ),
    .S0(net13),
    .S1(net277),
    .X(_1650_));
 sky130_fd_sc_hd__mux4_1 _5402_ (.A0(_1647_),
    .A1(_1648_),
    .A2(_1649_),
    .A3(_1650_),
    .S0(_0103_),
    .S1(net15),
    .X(_1651_));
 sky130_fd_sc_hd__a22o_4 _5403_ (.A1(net17),
    .A2(_1646_),
    .B1(_1651_),
    .B2(net184),
    .X(net158));
 sky130_fd_sc_hd__mux2_8 _5404_ (.A0(_3539_),
    .A1(net158),
    .S(net178),
    .X(_1652_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_100 ();
 sky130_fd_sc_hd__xnor2_1 _5408_ (.A(_0122_),
    .B(_1652_),
    .Y(_3508_));
 sky130_fd_sc_hd__inv_1 _5409_ (.A(_3508_),
    .Y(_3512_));
 sky130_fd_sc_hd__a221o_1 _5410_ (.A1(\dp.rf.rf[19][3] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][3] ),
    .C1(net191),
    .X(_1656_));
 sky130_fd_sc_hd__mux2i_1 _5411_ (.A0(\dp.rf.rf[22][3] ),
    .A1(\dp.rf.rf[23][3] ),
    .S(net210),
    .Y(_1657_));
 sky130_fd_sc_hd__a211oi_1 _5412_ (.A1(net208),
    .A2(_1657_),
    .B1(_0130_),
    .C1(net205),
    .Y(_1658_));
 sky130_fd_sc_hd__mux4_1 _5413_ (.A0(\dp.rf.rf[16][3] ),
    .A1(\dp.rf.rf[17][3] ),
    .A2(\dp.rf.rf[20][3] ),
    .A3(\dp.rf.rf[21][3] ),
    .S0(net210),
    .S1(net208),
    .X(_1659_));
 sky130_fd_sc_hd__nand2_1 _5414_ (.A(net205),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(_0232_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a21oi_1 _5416_ (.A1(_1656_),
    .A2(_1658_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__a21o_1 _5417_ (.A1(_0231_),
    .A2(_1095_),
    .B1(net197),
    .X(_1663_));
 sky130_fd_sc_hd__inv_1 _5418_ (.A(\dp.rf.rf[4][3] ),
    .Y(_1664_));
 sky130_fd_sc_hd__mux2i_1 _5419_ (.A0(\dp.rf.rf[1][3] ),
    .A1(\dp.rf.rf[5][3] ),
    .S(net208),
    .Y(_1665_));
 sky130_fd_sc_hd__a221oi_1 _5420_ (.A1(_1664_),
    .A2(net204),
    .B1(_1665_),
    .B2(net210),
    .C1(net8),
    .Y(_1666_));
 sky130_fd_sc_hd__nor3_1 _5421_ (.A(net11),
    .B(_0130_),
    .C(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand2_1 _5422_ (.A(_0231_),
    .B(_0347_),
    .Y(_1668_));
 sky130_fd_sc_hd__a21oi_1 _5423_ (.A1(_0119_),
    .A2(_1668_),
    .B1(\dp.rf.rf[0][3] ),
    .Y(_1669_));
 sky130_fd_sc_hd__mux2i_1 _5424_ (.A0(\dp.rf.rf[6][3] ),
    .A1(\dp.rf.rf[7][3] ),
    .S(net210),
    .Y(_1670_));
 sky130_fd_sc_hd__a21oi_1 _5425_ (.A1(net208),
    .A2(_1670_),
    .B1(net192),
    .Y(_1671_));
 sky130_fd_sc_hd__a221o_1 _5426_ (.A1(\dp.rf.rf[3][3] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[2][3] ),
    .C1(_0221_),
    .X(_1672_));
 sky130_fd_sc_hd__a2bb2oi_1 _5427_ (.A1_N(_1667_),
    .A2_N(_1669_),
    .B1(_1671_),
    .B2(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(\dp.rf.rf[26][3] ),
    .A1(\dp.rf.rf[30][3] ),
    .S(net208),
    .X(_1674_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(net210),
    .B(net208),
    .Y(_1675_));
 sky130_fd_sc_hd__o221ai_1 _5430_ (.A1(net210),
    .A2(_1674_),
    .B1(_1675_),
    .B2(\dp.rf.rf[31][3] ),
    .C1(net8),
    .Y(_1676_));
 sky130_fd_sc_hd__a2111oi_0 _5431_ (.A1(_0115_),
    .A2(_0117_),
    .B1(\dp.rf.rf[27][3] ),
    .C1(_0245_),
    .D1(net208),
    .Y(_1677_));
 sky130_fd_sc_hd__mux4_1 _5432_ (.A0(\dp.rf.rf[24][3] ),
    .A1(\dp.rf.rf[25][3] ),
    .A2(\dp.rf.rf[28][3] ),
    .A3(\dp.rf.rf[29][3] ),
    .S0(net210),
    .S1(net208),
    .X(_1678_));
 sky130_fd_sc_hd__nand2_1 _5433_ (.A(net205),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__o2111ai_1 _5434_ (.A1(_1676_),
    .A2(_1677_),
    .B1(_1679_),
    .C1(_0119_),
    .D1(net11),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(net186),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__a221o_1 _5436_ (.A1(\dp.rf.rf[11][3] ),
    .A2(net210),
    .B1(net200),
    .B2(\dp.rf.rf[10][3] ),
    .C1(net189),
    .X(_1682_));
 sky130_fd_sc_hd__mux2i_1 _5437_ (.A0(\dp.rf.rf[14][3] ),
    .A1(\dp.rf.rf[15][3] ),
    .S(net210),
    .Y(_1683_));
 sky130_fd_sc_hd__a21oi_1 _5438_ (.A1(net208),
    .A2(_1683_),
    .B1(net192),
    .Y(_1684_));
 sky130_fd_sc_hd__mux4_1 _5439_ (.A0(\dp.rf.rf[8][3] ),
    .A1(\dp.rf.rf[9][3] ),
    .A2(\dp.rf.rf[12][3] ),
    .A3(\dp.rf.rf[13][3] ),
    .S0(net210),
    .S1(net208),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _5440_ (.A(net205),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_0231_),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a21oi_1 _5442_ (.A1(_1682_),
    .A2(_1684_),
    .B1(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__o32a_4 _5443_ (.A1(_1662_),
    .A2(_1663_),
    .A3(_1673_),
    .B1(_1681_),
    .B2(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_99 ();
 sky130_fd_sc_hd__a22o_2 _5445_ (.A1(net32),
    .A2(_0042_),
    .B1(_1604_),
    .B2(net15),
    .X(_3535_));
 sky130_fd_sc_hd__mux4_1 _5446_ (.A0(\dp.rf.rf[24][2] ),
    .A1(\dp.rf.rf[25][2] ),
    .A2(\dp.rf.rf[26][2] ),
    .A3(\dp.rf.rf[27][2] ),
    .S0(net213),
    .S1(net277),
    .X(_1690_));
 sky130_fd_sc_hd__mux4_1 _5447_ (.A0(\dp.rf.rf[16][2] ),
    .A1(\dp.rf.rf[17][2] ),
    .A2(\dp.rf.rf[18][2] ),
    .A3(\dp.rf.rf[19][2] ),
    .S0(net213),
    .S1(net277),
    .X(_1691_));
 sky130_fd_sc_hd__mux4_2 _5448_ (.A0(\dp.rf.rf[28][2] ),
    .A1(\dp.rf.rf[29][2] ),
    .A2(\dp.rf.rf[30][2] ),
    .A3(\dp.rf.rf[31][2] ),
    .S0(net213),
    .S1(net277),
    .X(_1692_));
 sky130_fd_sc_hd__mux4_1 _5449_ (.A0(\dp.rf.rf[20][2] ),
    .A1(\dp.rf.rf[21][2] ),
    .A2(\dp.rf.rf[22][2] ),
    .A3(\dp.rf.rf[23][2] ),
    .S0(net213),
    .S1(net277),
    .X(_1693_));
 sky130_fd_sc_hd__mux4_2 _5450_ (.A0(_1690_),
    .A1(_1691_),
    .A2(_1692_),
    .A3(_1693_),
    .S0(_0103_),
    .S1(net15),
    .X(_1694_));
 sky130_fd_sc_hd__mux4_1 _5451_ (.A0(\dp.rf.rf[8][2] ),
    .A1(\dp.rf.rf[9][2] ),
    .A2(\dp.rf.rf[10][2] ),
    .A3(\dp.rf.rf[11][2] ),
    .S0(net13),
    .S1(net277),
    .X(_1695_));
 sky130_fd_sc_hd__mux4_1 _5452_ (.A0(\dp.rf.rf[0][2] ),
    .A1(\dp.rf.rf[1][2] ),
    .A2(\dp.rf.rf[2][2] ),
    .A3(\dp.rf.rf[3][2] ),
    .S0(net13),
    .S1(net277),
    .X(_1696_));
 sky130_fd_sc_hd__mux4_1 _5453_ (.A0(\dp.rf.rf[12][2] ),
    .A1(\dp.rf.rf[13][2] ),
    .A2(\dp.rf.rf[14][2] ),
    .A3(\dp.rf.rf[15][2] ),
    .S0(net13),
    .S1(net277),
    .X(_1697_));
 sky130_fd_sc_hd__mux4_1 _5454_ (.A0(\dp.rf.rf[4][2] ),
    .A1(\dp.rf.rf[5][2] ),
    .A2(\dp.rf.rf[6][2] ),
    .A3(\dp.rf.rf[7][2] ),
    .S0(net13),
    .S1(net277),
    .X(_1698_));
 sky130_fd_sc_hd__mux4_2 _5455_ (.A0(_1695_),
    .A1(_1696_),
    .A2(_1697_),
    .A3(_1698_),
    .S0(_0103_),
    .S1(net15),
    .X(_1699_));
 sky130_fd_sc_hd__a22oi_4 _5456_ (.A1(_1694_),
    .A2(net17),
    .B1(_1699_),
    .B2(net184),
    .Y(_1700_));
 sky130_fd_sc_hd__inv_1 _5457_ (.A(_1700_),
    .Y(net155));
 sky130_fd_sc_hd__nand2_4 _5458_ (.A(_1700_),
    .B(net178),
    .Y(_1701_));
 sky130_fd_sc_hd__o21a_4 _5459_ (.A1(net178),
    .A2(_3535_),
    .B1(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_97 ();
 sky130_fd_sc_hd__xnor2_1 _5462_ (.A(_0122_),
    .B(_1702_),
    .Y(_3516_));
 sky130_fd_sc_hd__inv_1 _5463_ (.A(_3516_),
    .Y(_3520_));
 sky130_fd_sc_hd__nor2b_1 _5464_ (.A(net208),
    .B_N(\dp.rf.rf[17][2] ),
    .Y(_1705_));
 sky130_fd_sc_hd__a211oi_2 _5465_ (.A1(net434),
    .A2(net208),
    .B1(_1705_),
    .C1(_0245_),
    .Y(_1706_));
 sky130_fd_sc_hd__o221ai_2 _5466_ (.A1(net436),
    .A2(_0528_),
    .B1(_0955_),
    .B2(\dp.rf.rf[16][2] ),
    .C1(net205),
    .Y(_1707_));
 sky130_fd_sc_hd__a221oi_2 _5467_ (.A1(\dp.rf.rf[19][2] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[18][2] ),
    .C1(_0221_),
    .Y(_1708_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(\dp.rf.rf[22][2] ),
    .A1(\dp.rf.rf[23][2] ),
    .S(net210),
    .X(_1709_));
 sky130_fd_sc_hd__o21ai_1 _5469_ (.A1(_0148_),
    .A2(_1709_),
    .B1(net8),
    .Y(_1710_));
 sky130_fd_sc_hd__o22ai_4 _5470_ (.A1(_1706_),
    .A2(_1707_),
    .B1(_1708_),
    .B2(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__nor2b_1 _5471_ (.A(net210),
    .B_N(\dp.rf.rf[30][2] ),
    .Y(_1712_));
 sky130_fd_sc_hd__a211oi_1 _5472_ (.A1(\dp.rf.rf[31][2] ),
    .A2(net210),
    .B1(_0148_),
    .C1(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__a221oi_1 _5473_ (.A1(\dp.rf.rf[27][2] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[26][2] ),
    .C1(_0221_),
    .Y(_1714_));
 sky130_fd_sc_hd__nor4_1 _5474_ (.A(_0212_),
    .B(_0963_),
    .C(_1713_),
    .D(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__nor2b_1 _5475_ (.A(net208),
    .B_N(\dp.rf.rf[25][2] ),
    .Y(_1716_));
 sky130_fd_sc_hd__a211oi_1 _5476_ (.A1(\dp.rf.rf[29][2] ),
    .A2(net208),
    .B1(_1716_),
    .C1(_0245_),
    .Y(_1717_));
 sky130_fd_sc_hd__o22ai_1 _5477_ (.A1(\dp.rf.rf[28][2] ),
    .A2(_0528_),
    .B1(_0955_),
    .B2(\dp.rf.rf[24][2] ),
    .Y(_1718_));
 sky130_fd_sc_hd__nor4_1 _5478_ (.A(net8),
    .B(_0963_),
    .C(_1717_),
    .D(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__a211oi_4 _5479_ (.A1(_0952_),
    .A2(_1711_),
    .B1(_1715_),
    .C1(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__mux4_1 _5480_ (.A0(\dp.rf.rf[10][2] ),
    .A1(\dp.rf.rf[11][2] ),
    .A2(\dp.rf.rf[14][2] ),
    .A3(\dp.rf.rf[15][2] ),
    .S0(net210),
    .S1(net208),
    .X(_1721_));
 sky130_fd_sc_hd__mux4_1 _5481_ (.A0(\dp.rf.rf[8][2] ),
    .A1(\dp.rf.rf[9][2] ),
    .A2(\dp.rf.rf[12][2] ),
    .A3(\dp.rf.rf[13][2] ),
    .S0(net210),
    .S1(net208),
    .X(_1722_));
 sky130_fd_sc_hd__mux2i_2 _5482_ (.A0(_1721_),
    .A1(_1722_),
    .S(net205),
    .Y(_1723_));
 sky130_fd_sc_hd__mux2i_1 _5483_ (.A0(\dp.rf.rf[6][2] ),
    .A1(\dp.rf.rf[7][2] ),
    .S(net210),
    .Y(_1724_));
 sky130_fd_sc_hd__a221oi_1 _5484_ (.A1(\dp.rf.rf[3][2] ),
    .A2(net210),
    .B1(_0176_),
    .B2(\dp.rf.rf[2][2] ),
    .C1(net191),
    .Y(_1725_));
 sky130_fd_sc_hd__a211o_1 _5485_ (.A1(net208),
    .A2(_1724_),
    .B1(_1725_),
    .C1(net192),
    .X(_1726_));
 sky130_fd_sc_hd__mux2i_1 _5486_ (.A0(\dp.rf.rf[1][2] ),
    .A1(\dp.rf.rf[5][2] ),
    .S(net208),
    .Y(_1727_));
 sky130_fd_sc_hd__nor2_1 _5487_ (.A(\dp.rf.rf[4][2] ),
    .B(_0528_),
    .Y(_1728_));
 sky130_fd_sc_hd__a211oi_1 _5488_ (.A1(net210),
    .A2(_1727_),
    .B1(_1728_),
    .C1(net8),
    .Y(_1729_));
 sky130_fd_sc_hd__o22ai_1 _5489_ (.A1(\dp.rf.rf[0][2] ),
    .A2(_0348_),
    .B1(_1729_),
    .B2(net197),
    .Y(_1730_));
 sky130_fd_sc_hd__a221o_4 _5490_ (.A1(net186),
    .A2(_1723_),
    .B1(_1726_),
    .B2(_1730_),
    .C1(_0271_),
    .X(_1731_));
 sky130_fd_sc_hd__nand2_4 _5491_ (.A(_1720_),
    .B(_1731_),
    .Y(_3515_));
 sky130_fd_sc_hd__inv_1 _5492_ (.A(_3515_),
    .Y(_3519_));
 sky130_fd_sc_hd__a22o_1 _5493_ (.A1(net31),
    .A2(_0042_),
    .B1(_1604_),
    .B2(net277),
    .X(_3272_));
 sky130_fd_sc_hd__a221oi_1 _5494_ (.A1(net16),
    .A2(\dp.rf.rf[8][1] ),
    .B1(_0081_),
    .B2(\dp.rf.rf[0][1] ),
    .C1(net15),
    .Y(_1732_));
 sky130_fd_sc_hd__inv_1 _5495_ (.A(\dp.rf.rf[4][1] ),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5496_ (.A(net16),
    .B(\dp.rf.rf[12][1] ),
    .Y(_1734_));
 sky130_fd_sc_hd__o211a_1 _5497_ (.A1(net16),
    .A2(_1733_),
    .B1(_1734_),
    .C1(net15),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_1 _5498_ (.A0(\dp.rf.rf[1][1] ),
    .A1(\dp.rf.rf[5][1] ),
    .A2(\dp.rf.rf[9][1] ),
    .A3(\dp.rf.rf[13][1] ),
    .S0(net15),
    .S1(net16),
    .X(_1736_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(net212),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__o31a_1 _5500_ (.A1(net212),
    .A2(_1732_),
    .A3(_1735_),
    .B1(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__mux2i_1 _5501_ (.A0(\dp.rf.rf[18][1] ),
    .A1(\dp.rf.rf[19][1] ),
    .S(net212),
    .Y(_1739_));
 sky130_fd_sc_hd__mux2i_1 _5502_ (.A0(\dp.rf.rf[24][1] ),
    .A1(\dp.rf.rf[25][1] ),
    .S(net212),
    .Y(_1740_));
 sky130_fd_sc_hd__a22oi_1 _5503_ (.A1(_0081_),
    .A2(_1739_),
    .B1(_1740_),
    .B2(_0061_),
    .Y(_1741_));
 sky130_fd_sc_hd__mux2i_1 _5504_ (.A0(\dp.rf.rf[26][1] ),
    .A1(\dp.rf.rf[27][1] ),
    .S(net212),
    .Y(_1742_));
 sky130_fd_sc_hd__mux2i_1 _5505_ (.A0(\dp.rf.rf[16][1] ),
    .A1(\dp.rf.rf[17][1] ),
    .S(net212),
    .Y(_1743_));
 sky130_fd_sc_hd__a22oi_1 _5506_ (.A1(_0066_),
    .A2(_1742_),
    .B1(_1743_),
    .B2(_0054_),
    .Y(_1744_));
 sky130_fd_sc_hd__nand3_1 _5507_ (.A(_0088_),
    .B(_1741_),
    .C(_1744_),
    .Y(_1745_));
 sky130_fd_sc_hd__mux4_1 _5508_ (.A0(\dp.rf.rf[6][1] ),
    .A1(\dp.rf.rf[7][1] ),
    .A2(\dp.rf.rf[14][1] ),
    .A3(\dp.rf.rf[15][1] ),
    .S0(net212),
    .S1(net16),
    .X(_1746_));
 sky130_fd_sc_hd__mux4_1 _5509_ (.A0(\dp.rf.rf[2][1] ),
    .A1(\dp.rf.rf[3][1] ),
    .A2(\dp.rf.rf[10][1] ),
    .A3(\dp.rf.rf[11][1] ),
    .S0(net212),
    .S1(net16),
    .X(_1747_));
 sky130_fd_sc_hd__mux2i_1 _5510_ (.A0(_1746_),
    .A1(_1747_),
    .S(_0286_),
    .Y(_1748_));
 sky130_fd_sc_hd__mux4_1 _5511_ (.A0(\dp.rf.rf[28][1] ),
    .A1(\dp.rf.rf[29][1] ),
    .A2(\dp.rf.rf[30][1] ),
    .A3(\dp.rf.rf[31][1] ),
    .S0(net212),
    .S1(net274),
    .X(_1749_));
 sky130_fd_sc_hd__mux4_1 _5512_ (.A0(\dp.rf.rf[20][1] ),
    .A1(\dp.rf.rf[21][1] ),
    .A2(\dp.rf.rf[22][1] ),
    .A3(\dp.rf.rf[23][1] ),
    .S0(net212),
    .S1(net274),
    .X(_1750_));
 sky130_fd_sc_hd__mux2i_1 _5513_ (.A0(_1749_),
    .A1(_1750_),
    .S(_0103_),
    .Y(_1751_));
 sky130_fd_sc_hd__o32a_1 _5514_ (.A1(net17),
    .A2(_0057_),
    .A3(_1748_),
    .B1(_1751_),
    .B2(_0101_),
    .X(_1752_));
 sky130_fd_sc_hd__o311ai_4 _5515_ (.A1(_1738_),
    .A2(net274),
    .A3(net17),
    .B1(_1745_),
    .C1(_1752_),
    .Y(net144));
 sky130_fd_sc_hd__a221o_2 _5516_ (.A1(net31),
    .A2(_0042_),
    .B1(_1604_),
    .B2(net277),
    .C1(net178),
    .X(_1753_));
 sky130_fd_sc_hd__o21a_4 _5517_ (.A1(net409),
    .A2(_0138_),
    .B1(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_93 ();
 sky130_fd_sc_hd__xnor2_2 _5522_ (.A(_0122_),
    .B(_1754_),
    .Y(_3267_));
 sky130_fd_sc_hd__inv_1 _5523_ (.A(_3267_),
    .Y(_3526_));
 sky130_fd_sc_hd__mux2i_1 _5524_ (.A0(\dp.rf.rf[24][1] ),
    .A1(\dp.rf.rf[28][1] ),
    .S(net206),
    .Y(_1759_));
 sky130_fd_sc_hd__mux2i_1 _5525_ (.A0(\dp.rf.rf[25][1] ),
    .A1(\dp.rf.rf[29][1] ),
    .S(net206),
    .Y(_1760_));
 sky130_fd_sc_hd__o22ai_1 _5526_ (.A1(_0170_),
    .A2(_1759_),
    .B1(_1760_),
    .B2(_0415_),
    .Y(_1761_));
 sky130_fd_sc_hd__o21ai_2 _5527_ (.A1(net198),
    .A2(_1761_),
    .B1(net187),
    .Y(_1762_));
 sky130_fd_sc_hd__nand4_1 _5528_ (.A(\dp.rf.rf[26][1] ),
    .B(net1),
    .C(net12),
    .D(net23),
    .Y(_1763_));
 sky130_fd_sc_hd__o2bb2ai_1 _5529_ (.A1_N(\dp.rf.rf[26][1] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__and2_0 _5530_ (.A(\dp.rf.rf[27][1] ),
    .B(net209),
    .X(_1765_));
 sky130_fd_sc_hd__mux2i_1 _5531_ (.A0(\dp.rf.rf[30][1] ),
    .A1(\dp.rf.rf[31][1] ),
    .S(net209),
    .Y(_1766_));
 sky130_fd_sc_hd__a21oi_1 _5532_ (.A1(net206),
    .A2(_1766_),
    .B1(_0231_),
    .Y(_1767_));
 sky130_fd_sc_hd__o311ai_4 _5533_ (.A1(_0221_),
    .A2(_1764_),
    .A3(_1765_),
    .B1(_1767_),
    .C1(net182),
    .Y(_1768_));
 sky130_fd_sc_hd__nand4_1 _5534_ (.A(\dp.rf.rf[18][1] ),
    .B(net1),
    .C(net12),
    .D(net23),
    .Y(_1769_));
 sky130_fd_sc_hd__o2bb2ai_1 _5535_ (.A1_N(\dp.rf.rf[18][1] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__and2_0 _5536_ (.A(\dp.rf.rf[19][1] ),
    .B(net209),
    .X(_1771_));
 sky130_fd_sc_hd__mux2i_1 _5537_ (.A0(\dp.rf.rf[22][1] ),
    .A1(\dp.rf.rf[23][1] ),
    .S(net209),
    .Y(_1772_));
 sky130_fd_sc_hd__nand2_1 _5538_ (.A(net206),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__o311ai_2 _5539_ (.A1(_0221_),
    .A2(_1770_),
    .A3(_1771_),
    .B1(_1773_),
    .C1(net182),
    .Y(_1774_));
 sky130_fd_sc_hd__inv_1 _5540_ (.A(\dp.rf.rf[20][1] ),
    .Y(_1775_));
 sky130_fd_sc_hd__mux2i_1 _5541_ (.A0(\dp.rf.rf[17][1] ),
    .A1(\dp.rf.rf[21][1] ),
    .S(net206),
    .Y(_1776_));
 sky130_fd_sc_hd__a221oi_1 _5542_ (.A1(_1775_),
    .A2(net203),
    .B1(_1776_),
    .B2(net209),
    .C1(net8),
    .Y(_1777_));
 sky130_fd_sc_hd__o22ai_2 _5543_ (.A1(\dp.rf.rf[16][1] ),
    .A2(net181),
    .B1(_1777_),
    .B2(net196),
    .Y(_1778_));
 sky130_fd_sc_hd__a22oi_4 _5544_ (.A1(_1762_),
    .A2(_1768_),
    .B1(_1774_),
    .B2(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand4_1 _5545_ (.A(\dp.rf.rf[10][1] ),
    .B(net1),
    .C(net12),
    .D(net23),
    .Y(_1780_));
 sky130_fd_sc_hd__o2bb2ai_1 _5546_ (.A1_N(\dp.rf.rf[10][1] ),
    .A2_N(_0245_),
    .B1(_0129_),
    .B2(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__and2_0 _5547_ (.A(\dp.rf.rf[11][1] ),
    .B(net209),
    .X(_1782_));
 sky130_fd_sc_hd__mux2i_1 _5548_ (.A0(\dp.rf.rf[14][1] ),
    .A1(\dp.rf.rf[15][1] ),
    .S(net209),
    .Y(_1783_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(net206),
    .B(_1783_),
    .Y(_1784_));
 sky130_fd_sc_hd__o311ai_4 _5550_ (.A1(_0221_),
    .A2(_1781_),
    .A3(_1782_),
    .B1(_1784_),
    .C1(net182),
    .Y(_1785_));
 sky130_fd_sc_hd__mux4_1 _5551_ (.A0(\dp.rf.rf[8][1] ),
    .A1(\dp.rf.rf[9][1] ),
    .A2(\dp.rf.rf[12][1] ),
    .A3(\dp.rf.rf[13][1] ),
    .S0(net209),
    .S1(net206),
    .X(_1786_));
 sky130_fd_sc_hd__a21oi_1 _5552_ (.A1(net205),
    .A2(_1786_),
    .B1(net199),
    .Y(_1787_));
 sky130_fd_sc_hd__mux4_1 _5553_ (.A0(\dp.rf.rf[2][1] ),
    .A1(\dp.rf.rf[3][1] ),
    .A2(\dp.rf.rf[6][1] ),
    .A3(\dp.rf.rf[7][1] ),
    .S0(net209),
    .S1(net206),
    .X(_1788_));
 sky130_fd_sc_hd__mux2i_1 _5554_ (.A0(\dp.rf.rf[1][1] ),
    .A1(\dp.rf.rf[5][1] ),
    .S(net206),
    .Y(_1789_));
 sky130_fd_sc_hd__a221oi_1 _5555_ (.A1(_1733_),
    .A2(net203),
    .B1(_1789_),
    .B2(net209),
    .C1(net8),
    .Y(_1790_));
 sky130_fd_sc_hd__a211oi_2 _5556_ (.A1(net8),
    .A2(_1788_),
    .B1(_1790_),
    .C1(net196),
    .Y(_1791_));
 sky130_fd_sc_hd__a211oi_4 _5557_ (.A1(_1785_),
    .A2(_1787_),
    .B1(_1791_),
    .C1(_0271_),
    .Y(_1792_));
 sky130_fd_sc_hd__nor2_4 _5558_ (.A(_1779_),
    .B(_1792_),
    .Y(_3525_));
 sky130_fd_sc_hd__inv_1 _5559_ (.A(net497),
    .Y(_3275_));
 sky130_fd_sc_hd__a21oi_4 _5560_ (.A1(net27),
    .A2(_0111_),
    .B1(_0108_),
    .Y(_1793_));
 sky130_fd_sc_hd__nor2_2 _5561_ (.A(_0121_),
    .B(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nand4b_4 _5562_ (.A_N(net4),
    .B(net5),
    .C(_1794_),
    .D(net6),
    .Y(_1795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_92 ();
 sky130_fd_sc_hd__or2_2 _5564_ (.A(net27),
    .B(_0108_),
    .X(_1797_));
 sky130_fd_sc_hd__nand2_2 _5565_ (.A(net5),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__nor2_1 _5566_ (.A(net6),
    .B(net4),
    .Y(_1799_));
 sky130_fd_sc_hd__a21oi_1 _5567_ (.A1(net6),
    .A2(net4),
    .B1(_1793_),
    .Y(_1800_));
 sky130_fd_sc_hd__nand2_2 _5568_ (.A(net6),
    .B(net4),
    .Y(_1801_));
 sky130_fd_sc_hd__a21oi_1 _5569_ (.A1(_1797_),
    .A2(_1801_),
    .B1(net5),
    .Y(_1802_));
 sky130_fd_sc_hd__a2111oi_4 _5570_ (.A1(_1798_),
    .A2(_1799_),
    .B1(_0121_),
    .C1(_1800_),
    .D1(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_91 ();
 sky130_fd_sc_hd__nor2_8 _5572_ (.A(net27),
    .B(_0108_),
    .Y(_1805_));
 sky130_fd_sc_hd__nand2b_4 _5573_ (.A_N(net5),
    .B(net4),
    .Y(_1806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__nor2b_1 _5575_ (.A(net6),
    .B_N(net24),
    .Y(_1808_));
 sky130_fd_sc_hd__nor4_4 _5576_ (.A(_0130_),
    .B(_1805_),
    .C(_1806_),
    .D(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_89 ();
 sky130_fd_sc_hd__a21oi_1 _5578_ (.A1(_3277_),
    .A2(net174),
    .B1(net176),
    .Y(_1811_));
 sky130_fd_sc_hd__o21ai_0 _5579_ (.A1(_3281_),
    .A2(_1795_),
    .B1(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(net6),
    .Y(_1813_));
 sky130_fd_sc_hd__and3_1 _5581_ (.A(_1813_),
    .B(_1797_),
    .C(_1793_),
    .X(_1814_));
 sky130_fd_sc_hd__o21ai_2 _5582_ (.A1(net5),
    .A2(_1814_),
    .B1(net4),
    .Y(_1815_));
 sky130_fd_sc_hd__nor2_1 _5583_ (.A(net4),
    .B(_1805_),
    .Y(_1816_));
 sky130_fd_sc_hd__o21ai_2 _5584_ (.A1(net5),
    .A2(_1816_),
    .B1(net6),
    .Y(_1817_));
 sky130_fd_sc_hd__a31o_4 _5585_ (.A1(_1798_),
    .A2(_1815_),
    .A3(_1817_),
    .B1(_0121_),
    .X(_1818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_88 ();
 sky130_fd_sc_hd__and3_4 _5587_ (.A(net6),
    .B(_0109_),
    .C(_1794_),
    .X(_1820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_86 ();
 sky130_fd_sc_hd__a21oi_1 _5590_ (.A1(_0122_),
    .A2(_1818_),
    .B1(_1820_),
    .Y(_1823_));
 sky130_fd_sc_hd__a31oi_4 _5591_ (.A1(_1798_),
    .A2(_1815_),
    .A3(_1817_),
    .B1(_0121_),
    .Y(_1824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_85 ();
 sky130_fd_sc_hd__nor2_1 _5593_ (.A(_0122_),
    .B(_1824_),
    .Y(_1826_));
 sky130_fd_sc_hd__nor2_1 _5594_ (.A(_3278_),
    .B(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__a21oi_1 _5595_ (.A1(_3278_),
    .A2(_1823_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor2b_1 _5596_ (.A(net6),
    .B_N(net5),
    .Y(_1829_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(net4),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__xor2_1 _5598_ (.A(_0274_),
    .B(_0300_),
    .X(_1831_));
 sky130_fd_sc_hd__o21ai_0 _5599_ (.A1(_1793_),
    .A2(_1830_),
    .B1(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hd__xnor2_1 _5600_ (.A(_0122_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__or3_1 _5601_ (.A(_3286_),
    .B(_3285_),
    .C(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_3285_),
    .B(_1833_),
    .Y(_1835_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_1794_),
    .B(_1829_),
    .Y(_1836_));
 sky130_fd_sc_hd__a21oi_1 _5604_ (.A1(_1834_),
    .A2(_1835_),
    .B1(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__nor3_1 _5605_ (.A(_1812_),
    .B(_1828_),
    .C(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__nor3_1 _5607_ (.A(_3357_),
    .B(_3373_),
    .C(_3365_),
    .Y(_1840_));
 sky130_fd_sc_hd__o21a_1 _5608_ (.A1(_3494_),
    .A2(_3493_),
    .B1(_3486_),
    .X(_1841_));
 sky130_fd_sc_hd__nor2_1 _5609_ (.A(_3485_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__a21o_1 _5610_ (.A1(_3518_),
    .A2(_3268_),
    .B1(_3517_),
    .X(_1843_));
 sky130_fd_sc_hd__a21o_1 _5611_ (.A1(_1843_),
    .A2(_3510_),
    .B1(_3509_),
    .X(_1844_));
 sky130_fd_sc_hd__a2111oi_4 _5612_ (.A1(_3502_),
    .A2(_1844_),
    .B1(_3493_),
    .C1(_3485_),
    .D1(_3501_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand4_2 _5613_ (.A(_3438_),
    .B(_3446_),
    .C(_3454_),
    .D(_3462_),
    .Y(_1846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_83 ();
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_3470_),
    .B(_3478_),
    .Y(_1848_));
 sky130_fd_sc_hd__nor4_4 _5616_ (.A(_1842_),
    .B(_1845_),
    .C(_1846_),
    .D(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__a21o_1 _5617_ (.A1(_3470_),
    .A2(_3477_),
    .B1(_3469_),
    .X(_1850_));
 sky130_fd_sc_hd__a21o_1 _5618_ (.A1(_3462_),
    .A2(_1850_),
    .B1(_3461_),
    .X(_1851_));
 sky130_fd_sc_hd__a2111oi_1 _5619_ (.A1(_3454_),
    .A2(_1851_),
    .B1(_3445_),
    .C1(_3437_),
    .D1(_3453_),
    .Y(_1852_));
 sky130_fd_sc_hd__or3_1 _5620_ (.A(_3437_),
    .B(_3446_),
    .C(_3445_),
    .X(_1853_));
 sky130_fd_sc_hd__o21ai_1 _5621_ (.A1(_3437_),
    .A2(_3438_),
    .B1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__nor2_1 _5622_ (.A(_3421_),
    .B(_3429_),
    .Y(_1855_));
 sky130_fd_sc_hd__o21ai_1 _5623_ (.A1(_1852_),
    .A2(_1854_),
    .B1(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__inv_1 _5624_ (.A(_3397_),
    .Y(_1857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__o21ai_0 _5626_ (.A1(_3405_),
    .A2(_3406_),
    .B1(_3398_),
    .Y(_1859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__nand2_1 _5628_ (.A(_3390_),
    .B(_3382_),
    .Y(_1861_));
 sky130_fd_sc_hd__a21oi_1 _5629_ (.A1(_1857_),
    .A2(_1859_),
    .B1(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__o21ai_0 _5630_ (.A1(_3430_),
    .A2(_3429_),
    .B1(_3422_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand2b_1 _5631_ (.A_N(_3421_),
    .B(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__and3_1 _5632_ (.A(_3414_),
    .B(_1862_),
    .C(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__o21ai_2 _5633_ (.A1(_1849_),
    .A2(_1856_),
    .B1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__inv_1 _5634_ (.A(_3382_),
    .Y(_1867_));
 sky130_fd_sc_hd__nand2_1 _5635_ (.A(_3405_),
    .B(_3398_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_1857_),
    .B(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__a21oi_1 _5637_ (.A1(_3390_),
    .A2(_1869_),
    .B1(_3389_),
    .Y(_1870_));
 sky130_fd_sc_hd__nor2_1 _5638_ (.A(_1867_),
    .B(_1870_),
    .Y(_1871_));
 sky130_fd_sc_hd__a211oi_1 _5639_ (.A1(_3413_),
    .A2(_1862_),
    .B1(_1871_),
    .C1(_3381_),
    .Y(_1872_));
 sky130_fd_sc_hd__nand3_2 _5640_ (.A(_1840_),
    .B(_1866_),
    .C(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__inv_1 _5641_ (.A(_3374_),
    .Y(_1874_));
 sky130_fd_sc_hd__o21a_1 _5642_ (.A1(_3366_),
    .A2(_3365_),
    .B1(_3358_),
    .X(_1875_));
 sky130_fd_sc_hd__o21ai_0 _5643_ (.A1(_3357_),
    .A2(_1875_),
    .B1(_3350_),
    .Y(_1876_));
 sky130_fd_sc_hd__a21oi_1 _5644_ (.A1(_1874_),
    .A2(_1840_),
    .B1(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__a2111oi_4 _5645_ (.A1(_1873_),
    .A2(_1877_),
    .B1(_3341_),
    .C1(_3333_),
    .D1(_3349_),
    .Y(_1878_));
 sky130_fd_sc_hd__or2_0 _5646_ (.A(_3341_),
    .B(_3342_),
    .X(_1879_));
 sky130_fd_sc_hd__a21oi_1 _5647_ (.A1(_3334_),
    .A2(_1879_),
    .B1(_3333_),
    .Y(_1880_));
 sky130_fd_sc_hd__nand2_1 _5648_ (.A(_3318_),
    .B(_3326_),
    .Y(_1881_));
 sky130_fd_sc_hd__a21oi_1 _5649_ (.A1(_3318_),
    .A2(_3325_),
    .B1(_3317_),
    .Y(_1882_));
 sky130_fd_sc_hd__o31ai_2 _5650_ (.A1(_1878_),
    .A2(_1880_),
    .A3(_1881_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__and2_0 _5651_ (.A(_3302_),
    .B(_3310_),
    .X(_1884_));
 sky130_fd_sc_hd__a221o_1 _5652_ (.A1(_3302_),
    .A2(_3309_),
    .B1(_1883_),
    .B2(_1884_),
    .C1(_3301_),
    .X(_1885_));
 sky130_fd_sc_hd__a21oi_2 _5653_ (.A1(_3294_),
    .A2(_1885_),
    .B1(_3293_),
    .Y(_1886_));
 sky130_fd_sc_hd__or4bb_1 _5654_ (.A(_1836_),
    .B(_1886_),
    .C_N(_1833_),
    .D_N(_3286_),
    .X(_1887_));
 sky130_fd_sc_hd__nor3_1 _5655_ (.A(_3285_),
    .B(_1836_),
    .C(_1833_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_2 _5656_ (.A(_1886_),
    .B(_1888_),
    .Y(_1889_));
 sky130_fd_sc_hd__mux2i_4 _5657_ (.A0(_3539_),
    .A1(net158),
    .S(net178),
    .Y(_1890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__o22ai_4 _5660_ (.A1(net179),
    .A2(_3530_),
    .B1(_0099_),
    .B2(net606),
    .Y(_1893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__inv_1 _5663_ (.A(_3495_),
    .Y(_3491_));
 sky130_fd_sc_hd__o21ai_4 _5664_ (.A1(net409),
    .A2(_0138_),
    .B1(_1753_),
    .Y(_1896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__nor2_1 _5668_ (.A(_3479_),
    .B(net407),
    .Y(_1900_));
 sky130_fd_sc_hd__a21oi_1 _5669_ (.A1(_3491_),
    .A2(net708),
    .B1(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__inv_1 _5670_ (.A(net515),
    .Y(_3483_));
 sky130_fd_sc_hd__nand2_1 _5671_ (.A(_3503_),
    .B(net709),
    .Y(_1902_));
 sky130_fd_sc_hd__o211ai_1 _5672_ (.A1(_3483_),
    .A2(net407),
    .B1(_1902_),
    .C1(net276),
    .Y(_1903_));
 sky130_fd_sc_hd__o21ai_1 _5673_ (.A1(net257),
    .A2(_1901_),
    .B1(_1903_),
    .Y(_1904_));
 sky130_fd_sc_hd__inv_1 _5674_ (.A(_1689_),
    .Y(_3507_));
 sky130_fd_sc_hd__nor2_1 _5675_ (.A(net265),
    .B(_3525_),
    .Y(_1905_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__a211oi_1 _5678_ (.A1(_3507_),
    .A2(net265),
    .B1(_1905_),
    .C1(net276),
    .Y(_1908_));
 sky130_fd_sc_hd__nor2_1 _5679_ (.A(net497),
    .B(net265),
    .Y(_1909_));
 sky130_fd_sc_hd__a211oi_1 _5680_ (.A1(_3515_),
    .A2(net265),
    .B1(_1909_),
    .C1(_0140_),
    .Y(_1910_));
 sky130_fd_sc_hd__nor3_1 _5681_ (.A(_1702_),
    .B(_1908_),
    .C(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__a21oi_1 _5682_ (.A1(net267),
    .A2(_1904_),
    .B1(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__mux2i_2 _5685_ (.A0(_3423_),
    .A1(_3439_),
    .S(net708),
    .Y(_1915_));
 sky130_fd_sc_hd__mux2i_2 _5686_ (.A0(_3415_),
    .A1(_3431_),
    .S(net708),
    .Y(_1916_));
 sky130_fd_sc_hd__mux2i_1 _5687_ (.A0(_1915_),
    .A1(_1916_),
    .S(_0140_),
    .Y(_1917_));
 sky130_fd_sc_hd__mux2i_2 _5688_ (.A0(_3447_),
    .A1(net855),
    .S(net708),
    .Y(_1918_));
 sky130_fd_sc_hd__mux2i_2 _5689_ (.A0(_3455_),
    .A1(_3471_),
    .S(net708),
    .Y(_1919_));
 sky130_fd_sc_hd__mux2i_2 _5690_ (.A0(_1918_),
    .A1(_1919_),
    .S(net257),
    .Y(_1920_));
 sky130_fd_sc_hd__o21ai_4 _5691_ (.A1(net178),
    .A2(_3535_),
    .B1(net432),
    .Y(_1921_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__mux2i_1 _5694_ (.A0(_1917_),
    .A1(_1920_),
    .S(_1921_),
    .Y(_1924_));
 sky130_fd_sc_hd__nor2_1 _5695_ (.A(net171),
    .B(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__a211oi_1 _5696_ (.A1(_1890_),
    .A2(_1912_),
    .B1(_1925_),
    .C1(net266),
    .Y(_1926_));
 sky130_fd_sc_hd__mux2_8 _5697_ (.A0(_1605_),
    .A1(net429),
    .S(net178),
    .X(_1927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__mux2i_4 _5700_ (.A0(_0371_),
    .A1(_3311_),
    .S(net167),
    .Y(_1930_));
 sky130_fd_sc_hd__mux2i_4 _5701_ (.A0(_0274_),
    .A1(_3303_),
    .S(net167),
    .Y(_1931_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(_1930_),
    .A1(_1931_),
    .S(_0140_),
    .X(_1932_));
 sky130_fd_sc_hd__mux2i_2 _5703_ (.A0(_0621_),
    .A1(_3343_),
    .S(net167),
    .Y(_1933_));
 sky130_fd_sc_hd__mux2i_2 _5704_ (.A0(_3319_),
    .A1(_3335_),
    .S(net167),
    .Y(_1934_));
 sky130_fd_sc_hd__mux2_2 _5705_ (.A0(_1933_),
    .A1(_1934_),
    .S(_0140_),
    .X(_1935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(_1932_),
    .A1(_1935_),
    .S(net165),
    .X(_1937_));
 sky130_fd_sc_hd__mux2i_4 _5708_ (.A0(_3359_),
    .A1(_3375_),
    .S(net167),
    .Y(_1938_));
 sky130_fd_sc_hd__mux2i_2 _5709_ (.A0(_3351_),
    .A1(_3367_),
    .S(net167),
    .Y(_1939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__mux2i_1 _5711_ (.A0(_1938_),
    .A1(_1939_),
    .S(_0140_),
    .Y(_1941_));
 sky130_fd_sc_hd__mux2i_2 _5712_ (.A0(_1031_),
    .A1(_3407_),
    .S(net167),
    .Y(_1942_));
 sky130_fd_sc_hd__mux2i_1 _5713_ (.A0(_3383_),
    .A1(_3399_),
    .S(net167),
    .Y(_1943_));
 sky130_fd_sc_hd__mux2i_1 _5714_ (.A0(_1942_),
    .A1(_1943_),
    .S(_0140_),
    .Y(_1944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__mux2i_1 _5716_ (.A0(_1941_),
    .A1(_1944_),
    .S(net165),
    .Y(_1946_));
 sky130_fd_sc_hd__mux2i_1 _5717_ (.A0(_1937_),
    .A1(_1946_),
    .S(_1890_),
    .Y(_1947_));
 sky130_fd_sc_hd__nor2_1 _5718_ (.A(_1927_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nor3_4 _5719_ (.A(net5),
    .B(_1805_),
    .C(_1801_),
    .Y(_1949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__o21ai_2 _5722_ (.A1(_1926_),
    .A2(_1948_),
    .B1(_1949_),
    .Y(_1952_));
 sky130_fd_sc_hd__nor3_2 _5723_ (.A(_0140_),
    .B(net497),
    .C(net265),
    .Y(_1953_));
 sky130_fd_sc_hd__nor2_4 _5724_ (.A(_1652_),
    .B(net421),
    .Y(_1954_));
 sky130_fd_sc_hd__nor2_8 _5725_ (.A(net438),
    .B(_1949_),
    .Y(_1955_));
 sky130_fd_sc_hd__or4_4 _5726_ (.A(_0130_),
    .B(_1805_),
    .C(_1806_),
    .D(_1808_),
    .X(_1956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__a31oi_4 _5729_ (.A1(_1953_),
    .A2(_1954_),
    .A3(_1955_),
    .B1(_1956_),
    .Y(_1959_));
 sky130_fd_sc_hd__a32oi_4 _5730_ (.A1(_1838_),
    .A2(_1887_),
    .A3(_1889_),
    .B1(_1952_),
    .B2(_1959_),
    .Y(net66));
 sky130_fd_sc_hd__or3_4 _5731_ (.A(net27),
    .B(net28),
    .C(_0108_),
    .X(_1960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__inv_12 _5733_ (.A(_1960_),
    .Y(net98));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__inv_1 _5736_ (.A(_3525_),
    .Y(_3266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__mux2i_2 _5739_ (.A0(_3311_),
    .A1(_0621_),
    .S(net167),
    .Y(_1966_));
 sky130_fd_sc_hd__mux2_2 _5740_ (.A0(_1934_),
    .A1(_1966_),
    .S(_0140_),
    .X(_1967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__nor3_1 _5742_ (.A(net253),
    .B(_0371_),
    .C(net265),
    .Y(_1969_));
 sky130_fd_sc_hd__a21o_2 _5743_ (.A1(net255),
    .A2(_1931_),
    .B1(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(_1967_),
    .A1(_1970_),
    .S(net425),
    .X(_1971_));
 sky130_fd_sc_hd__inv_1 _5745_ (.A(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__mux2i_2 _5747_ (.A0(_0371_),
    .A1(_3303_),
    .S(net252),
    .Y(_1974_));
 sky130_fd_sc_hd__nor2_1 _5748_ (.A(_0274_),
    .B(net167),
    .Y(_1975_));
 sky130_fd_sc_hd__a21o_2 _5749_ (.A1(net167),
    .A2(_1974_),
    .B1(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__mux2i_4 _5750_ (.A0(_1967_),
    .A1(_1976_),
    .S(net423),
    .Y(_1977_));
 sky130_fd_sc_hd__mux2i_2 _5751_ (.A0(_1972_),
    .A1(_1977_),
    .S(net24),
    .Y(_1978_));
 sky130_fd_sc_hd__nor2_1 _5752_ (.A(_0140_),
    .B(_1939_),
    .Y(_1979_));
 sky130_fd_sc_hd__mux2i_2 _5753_ (.A0(_3343_),
    .A1(_3359_),
    .S(net167),
    .Y(_1980_));
 sky130_fd_sc_hd__nor2_1 _5754_ (.A(net261),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__nor2_2 _5755_ (.A(_1979_),
    .B(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__mux2i_1 _5756_ (.A0(_3375_),
    .A1(_1031_),
    .S(net167),
    .Y(_1983_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_0140_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__nand2_1 _5759_ (.A(net169),
    .B(_1943_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_2 _5760_ (.A(_1984_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__mux2i_2 _5761_ (.A0(_1982_),
    .A1(_1987_),
    .S(net166),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5762_ (.A(net171),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__or3_4 _5763_ (.A(net5),
    .B(_1805_),
    .C(_1801_),
    .X(_1990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__nor2_2 _5766_ (.A(_1927_),
    .B(_1990_),
    .Y(_1993_));
 sky130_fd_sc_hd__o211ai_2 _5767_ (.A1(net171),
    .A2(_1978_),
    .B1(_1989_),
    .C1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__nor2_2 _5768_ (.A(net437),
    .B(_1990_),
    .Y(_1995_));
 sky130_fd_sc_hd__mux2i_2 _5769_ (.A0(_3407_),
    .A1(_3423_),
    .S(net707),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5770_ (.A(_0140_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _5771_ (.A(net257),
    .B(_1916_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__nor2_1 _5773_ (.A(_0140_),
    .B(_1918_),
    .Y(_2000_));
 sky130_fd_sc_hd__mux2i_1 _5774_ (.A0(_3439_),
    .A1(_3455_),
    .S(net708),
    .Y(_2001_));
 sky130_fd_sc_hd__nor2_1 _5775_ (.A(net257),
    .B(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nor2_1 _5776_ (.A(_2000_),
    .B(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__mux2i_2 _5778_ (.A0(_1999_),
    .A1(_2003_),
    .S(net932),
    .Y(_2005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__mux2i_1 _5781_ (.A0(_3471_),
    .A1(net517),
    .S(net407),
    .Y(_2008_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_0140_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__o21ai_1 _5783_ (.A1(_0140_),
    .A2(_1901_),
    .B1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__mux2i_1 _5784_ (.A0(_3503_),
    .A1(_1689_),
    .S(net257),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _5785_ (.A(net265),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__nand2_1 _5787_ (.A(net257),
    .B(_3525_),
    .Y(_2014_));
 sky130_fd_sc_hd__o211ai_1 _5788_ (.A1(net257),
    .A2(_3515_),
    .B1(net407),
    .C1(_2014_),
    .Y(_2015_));
 sky130_fd_sc_hd__nand3_1 _5789_ (.A(net932),
    .B(_2012_),
    .C(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__o211ai_1 _5790_ (.A1(net932),
    .A2(_2010_),
    .B1(_2016_),
    .C1(net171),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_0 _5791_ (.A1(net171),
    .A2(_2005_),
    .B1(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__nand2_1 _5792_ (.A(_1954_),
    .B(_1955_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _5793_ (.A(_0140_),
    .B(net497),
    .Y(_2020_));
 sky130_fd_sc_hd__nand3_2 _5794_ (.A(net709),
    .B(_2014_),
    .C(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__o21ai_0 _5795_ (.A1(_2019_),
    .A2(_2021_),
    .B1(net177),
    .Y(_2022_));
 sky130_fd_sc_hd__a21oi_1 _5796_ (.A1(_1995_),
    .A2(_2018_),
    .B1(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__nor2_1 _5797_ (.A(_3269_),
    .B(_1824_),
    .Y(_2024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__nand2_1 _5799_ (.A(_3524_),
    .B(_1820_),
    .Y(_2026_));
 sky130_fd_sc_hd__o21ai_0 _5800_ (.A1(_3527_),
    .A2(_1795_),
    .B1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__a2111oi_1 _5801_ (.A1(_3523_),
    .A2(net172),
    .B1(_2024_),
    .C1(_2027_),
    .D1(net177),
    .Y(_2028_));
 sky130_fd_sc_hd__a21oi_2 _5802_ (.A1(_1994_),
    .A2(_2023_),
    .B1(_2028_),
    .Y(net77));
 sky130_fd_sc_hd__mux2i_4 _5803_ (.A0(_3399_),
    .A1(_3415_),
    .S(net707),
    .Y(_2029_));
 sky130_fd_sc_hd__mux2i_2 _5804_ (.A0(_1996_),
    .A1(_2029_),
    .S(_0140_),
    .Y(_2030_));
 sky130_fd_sc_hd__mux2i_2 _5805_ (.A0(_3431_),
    .A1(_3447_),
    .S(net708),
    .Y(_2031_));
 sky130_fd_sc_hd__mux2i_1 _5806_ (.A0(_2001_),
    .A1(_2031_),
    .S(_0140_),
    .Y(_2032_));
 sky130_fd_sc_hd__mux2i_1 _5807_ (.A0(_2030_),
    .A1(_2032_),
    .S(_1921_),
    .Y(_2033_));
 sky130_fd_sc_hd__mux2i_2 _5808_ (.A0(net856),
    .A1(_3479_),
    .S(net407),
    .Y(_2034_));
 sky130_fd_sc_hd__mux2i_1 _5809_ (.A0(_2008_),
    .A1(_2034_),
    .S(_0140_),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_1689_),
    .B(net407),
    .Y(_2036_));
 sky130_fd_sc_hd__o21ai_0 _5811_ (.A1(_3491_),
    .A2(net407),
    .B1(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__a21oi_4 _5812_ (.A1(_1720_),
    .A2(_1731_),
    .B1(net466),
    .Y(_2038_));
 sky130_fd_sc_hd__a211oi_1 _5813_ (.A1(_3499_),
    .A2(net265),
    .B1(_2038_),
    .C1(_0140_),
    .Y(_2039_));
 sky130_fd_sc_hd__a21oi_1 _5814_ (.A1(_0140_),
    .A2(_2037_),
    .B1(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__nand2_1 _5815_ (.A(net932),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__o211ai_1 _5816_ (.A1(net932),
    .A2(_2035_),
    .B1(_2041_),
    .C1(net171),
    .Y(_2042_));
 sky130_fd_sc_hd__o21ai_0 _5817_ (.A1(net171),
    .A2(_2033_),
    .B1(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__mux2i_4 _5819_ (.A0(_3335_),
    .A1(_3351_),
    .S(net167),
    .Y(_2045_));
 sky130_fd_sc_hd__mux2i_4 _5820_ (.A0(_1980_),
    .A1(_2045_),
    .S(_0140_),
    .Y(_2046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__mux2i_2 _5822_ (.A0(_3367_),
    .A1(_3383_),
    .S(net167),
    .Y(_2048_));
 sky130_fd_sc_hd__mux2_1 _5823_ (.A0(_1983_),
    .A1(_2048_),
    .S(_0140_),
    .X(_2049_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(net165),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21ai_2 _5825_ (.A1(net165),
    .A2(_2046_),
    .B1(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__mux2i_4 _5826_ (.A0(_3303_),
    .A1(_3319_),
    .S(net167),
    .Y(_2052_));
 sky130_fd_sc_hd__mux2i_4 _5827_ (.A0(_1966_),
    .A1(_2052_),
    .S(_0140_),
    .Y(_2053_));
 sky130_fd_sc_hd__mux2i_1 _5828_ (.A0(_0274_),
    .A1(_0371_),
    .S(net253),
    .Y(_2054_));
 sky130_fd_sc_hd__a21oi_1 _5829_ (.A1(net167),
    .A2(_2054_),
    .B1(net165),
    .Y(_2055_));
 sky130_fd_sc_hd__a21oi_4 _5830_ (.A1(net165),
    .A2(_2053_),
    .B1(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_2 _5831_ (.A(net167),
    .B(_2054_),
    .Y(_2057_));
 sky130_fd_sc_hd__nor2_1 _5832_ (.A(net165),
    .B(_1975_),
    .Y(_2058_));
 sky130_fd_sc_hd__a22oi_4 _5833_ (.A1(net165),
    .A2(_2053_),
    .B1(_2057_),
    .B2(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__mux2i_1 _5834_ (.A0(_2056_),
    .A1(_2059_),
    .S(net24),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5835_ (.A(net465),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__o211ai_1 _5836_ (.A1(net431),
    .A2(_2051_),
    .B1(_2061_),
    .C1(net437),
    .Y(_2062_));
 sky130_fd_sc_hd__o21a_1 _5837_ (.A1(net266),
    .A2(_2043_),
    .B1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__nor2_2 _5838_ (.A(net499),
    .B(_1896_),
    .Y(_2064_));
 sky130_fd_sc_hd__o21ai_1 _5839_ (.A1(net466),
    .A2(_3525_),
    .B1(_0140_),
    .Y(_2065_));
 sky130_fd_sc_hd__o31ai_4 _5840_ (.A1(_0140_),
    .A2(_2038_),
    .A3(_2064_),
    .B1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__nor2_1 _5841_ (.A(_2019_),
    .B(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nor2_1 _5842_ (.A(_1956_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__xor2_1 _5845_ (.A(net605),
    .B(net271),
    .X(_2071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_3518_),
    .B(_1820_),
    .Y(_2073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__o211ai_1 _5849_ (.A1(_3521_),
    .A2(_1795_),
    .B1(_2073_),
    .C1(_1956_),
    .Y(_2075_));
 sky130_fd_sc_hd__a221oi_2 _5850_ (.A1(_3517_),
    .A2(net172),
    .B1(_1818_),
    .B2(_2071_),
    .C1(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__o22ai_2 _5851_ (.A1(_1990_),
    .A2(_2063_),
    .B1(_2068_),
    .B2(_2076_),
    .Y(net88));
 sky130_fd_sc_hd__nand2_4 _5852_ (.A(_0122_),
    .B(net168),
    .Y(_2077_));
 sky130_fd_sc_hd__and2_4 _5853_ (.A(_2077_),
    .B(_2020_),
    .X(_3265_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__mux2i_4 _5855_ (.A0(_1930_),
    .A1(_2052_),
    .S(net253),
    .Y(_2079_));
 sky130_fd_sc_hd__nor3_2 _5856_ (.A(_0140_),
    .B(_0274_),
    .C(net265),
    .Y(_2080_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(net422),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__o21ai_2 _5858_ (.A1(net267),
    .A2(_2079_),
    .B1(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__inv_2 _5859_ (.A(_0274_),
    .Y(_3284_));
 sky130_fd_sc_hd__nor2_1 _5860_ (.A(_3284_),
    .B(net165),
    .Y(_2083_));
 sky130_fd_sc_hd__a21oi_1 _5861_ (.A1(net165),
    .A2(_2079_),
    .B1(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__mux2i_1 _5862_ (.A0(_2082_),
    .A1(_2084_),
    .S(net24),
    .Y(_2085_));
 sky130_fd_sc_hd__mux2i_4 _5863_ (.A0(_1933_),
    .A1(_2045_),
    .S(net248),
    .Y(_2086_));
 sky130_fd_sc_hd__mux2i_4 _5864_ (.A0(_1938_),
    .A1(_2048_),
    .S(net261),
    .Y(_2087_));
 sky130_fd_sc_hd__mux2i_4 _5865_ (.A0(_2086_),
    .A1(_2087_),
    .S(net166),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(net171),
    .B(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__o21ai_0 _5867_ (.A1(net171),
    .A2(_2085_),
    .B1(_2089_),
    .Y(_2090_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_1993_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__nor2_1 _5869_ (.A(net257),
    .B(net518),
    .Y(_2092_));
 sky130_fd_sc_hd__a21oi_1 _5870_ (.A1(net257),
    .A2(_3491_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(net407),
    .B(_2011_),
    .Y(_2094_));
 sky130_fd_sc_hd__o21ai_0 _5872_ (.A1(net407),
    .A2(_2093_),
    .B1(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__mux2i_2 _5873_ (.A0(_1919_),
    .A1(_2034_),
    .S(net257),
    .Y(_2096_));
 sky130_fd_sc_hd__nor2_1 _5874_ (.A(net932),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__a21oi_1 _5875_ (.A1(net932),
    .A2(_2095_),
    .B1(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__mux2i_4 _5876_ (.A0(_1942_),
    .A1(_2029_),
    .S(net261),
    .Y(_2099_));
 sky130_fd_sc_hd__mux2i_2 _5877_ (.A0(_1915_),
    .A1(_2031_),
    .S(net257),
    .Y(_2100_));
 sky130_fd_sc_hd__mux2i_2 _5878_ (.A0(_2099_),
    .A1(_2100_),
    .S(_1921_),
    .Y(_2101_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(net431),
    .B(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__o21ai_0 _5880_ (.A1(net431),
    .A2(_2098_),
    .B1(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__o221ai_1 _5882_ (.A1(_0138_),
    .A2(net411),
    .B1(_1779_),
    .B2(_1792_),
    .C1(_1753_),
    .Y(_2105_));
 sky130_fd_sc_hd__o211ai_2 _5883_ (.A1(_1689_),
    .A2(net265),
    .B1(_2105_),
    .C1(net261),
    .Y(_2106_));
 sky130_fd_sc_hd__o31ai_4 _5884_ (.A1(net261),
    .A2(_2038_),
    .A3(_2064_),
    .B1(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__o21ai_0 _5886_ (.A1(_2019_),
    .A2(_2107_),
    .B1(net177),
    .Y(_2109_));
 sky130_fd_sc_hd__a21oi_1 _5887_ (.A1(_1995_),
    .A2(_2103_),
    .B1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__and3_1 _5890_ (.A(_3524_),
    .B(_2077_),
    .C(_2020_),
    .X(_2113_));
 sky130_fd_sc_hd__o21a_1 _5891_ (.A1(_3523_),
    .A2(_2113_),
    .B1(net270),
    .X(_2114_));
 sky130_fd_sc_hd__nor2_1 _5892_ (.A(_3517_),
    .B(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__xnor2_1 _5893_ (.A(net435),
    .B(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(net435),
    .B(_1820_),
    .Y(_2119_));
 sky130_fd_sc_hd__o211ai_1 _5897_ (.A1(_3513_),
    .A2(_1795_),
    .B1(_2119_),
    .C1(_1956_),
    .Y(_2120_));
 sky130_fd_sc_hd__a221oi_2 _5898_ (.A1(_3509_),
    .A2(net172),
    .B1(_1818_),
    .B2(_2116_),
    .C1(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a21oi_1 _5899_ (.A1(_2091_),
    .A2(_2110_),
    .B1(_2121_),
    .Y(net91));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_1927_),
    .B(net177),
    .Y(_2122_));
 sky130_fd_sc_hd__o211ai_2 _5901_ (.A1(_3515_),
    .A2(net407),
    .B1(_1902_),
    .C1(net257),
    .Y(_2123_));
 sky130_fd_sc_hd__o211ai_2 _5902_ (.A1(net407),
    .A2(_3266_),
    .B1(_2036_),
    .C1(_0140_),
    .Y(_2124_));
 sky130_fd_sc_hd__nor2_1 _5903_ (.A(net166),
    .B(_1953_),
    .Y(_2125_));
 sky130_fd_sc_hd__a31oi_2 _5904_ (.A1(net166),
    .A2(_2123_),
    .A3(_2124_),
    .B1(_2125_),
    .Y(_2126_));
 sky130_fd_sc_hd__nor2_1 _5905_ (.A(_1949_),
    .B(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__nor2_1 _5906_ (.A(_1921_),
    .B(_1920_),
    .Y(_2128_));
 sky130_fd_sc_hd__a211oi_1 _5907_ (.A1(net932),
    .A2(_1904_),
    .B1(_2128_),
    .C1(_1990_),
    .Y(_2129_));
 sky130_fd_sc_hd__nor3_1 _5908_ (.A(net431),
    .B(_2127_),
    .C(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__nor2_1 _5909_ (.A(net165),
    .B(_1944_),
    .Y(_2131_));
 sky130_fd_sc_hd__nor2_1 _5910_ (.A(net267),
    .B(_1917_),
    .Y(_2132_));
 sky130_fd_sc_hd__nor2_1 _5911_ (.A(_2131_),
    .B(_2132_),
    .Y(_2133_));
 sky130_fd_sc_hd__nor3_1 _5912_ (.A(net171),
    .B(_1990_),
    .C(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__or3_1 _5913_ (.A(_2122_),
    .B(_2130_),
    .C(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_1818_),
    .B(net279),
    .Y(_2136_));
 sky130_fd_sc_hd__nor2_1 _5915_ (.A(_1824_),
    .B(_1844_),
    .Y(_2137_));
 sky130_fd_sc_hd__o21ai_0 _5916_ (.A1(_1820_),
    .A2(_2137_),
    .B1(_3502_),
    .Y(_2138_));
 sky130_fd_sc_hd__o21ai_0 _5917_ (.A1(_3505_),
    .A2(_1795_),
    .B1(_1956_),
    .Y(_2139_));
 sky130_fd_sc_hd__a21oi_1 _5918_ (.A1(_3501_),
    .A2(net172),
    .B1(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hd__o211ai_1 _5919_ (.A1(_3502_),
    .A2(_2136_),
    .B1(_2138_),
    .C1(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__nor2_1 _5920_ (.A(net431),
    .B(_1935_),
    .Y(_2142_));
 sky130_fd_sc_hd__and2_2 _5921_ (.A(net24),
    .B(_1949_),
    .X(_2143_));
 sky130_fd_sc_hd__nand2_2 _5922_ (.A(_3284_),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__mux2i_4 _5923_ (.A0(_1930_),
    .A1(_1931_),
    .S(_0140_),
    .Y(_2145_));
 sky130_fd_sc_hd__nand2_2 _5924_ (.A(_1652_),
    .B(net166),
    .Y(_2146_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(_1938_),
    .A1(_1939_),
    .S(_0140_),
    .X(_2147_));
 sky130_fd_sc_hd__mux2i_2 _5926_ (.A0(_1935_),
    .A1(_2147_),
    .S(net165),
    .Y(_2148_));
 sky130_fd_sc_hd__o22ai_1 _5927_ (.A1(_2145_),
    .A2(_2146_),
    .B1(_2148_),
    .B2(net465),
    .Y(_2149_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(_1949_),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__nor2_2 _5929_ (.A(_1927_),
    .B(_1956_),
    .Y(_2151_));
 sky130_fd_sc_hd__o311ai_1 _5930_ (.A1(net166),
    .A2(_2142_),
    .A3(_2144_),
    .B1(_2150_),
    .C1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__and3_1 _5931_ (.A(_2135_),
    .B(_2141_),
    .C(_2152_),
    .X(net92));
 sky130_fd_sc_hd__nor2_1 _5932_ (.A(_3497_),
    .B(_1795_),
    .Y(_2153_));
 sky130_fd_sc_hd__a221o_1 _5933_ (.A1(_3493_),
    .A2(net172),
    .B1(_1820_),
    .B2(_3494_),
    .C1(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__a21oi_1 _5934_ (.A1(_3523_),
    .A2(net270),
    .B1(_3517_),
    .Y(_2155_));
 sky130_fd_sc_hd__nor2b_1 _5935_ (.A(_2155_),
    .B_N(_3510_),
    .Y(_2156_));
 sky130_fd_sc_hd__o21ai_1 _5936_ (.A1(_3509_),
    .A2(_2156_),
    .B1(_3502_),
    .Y(_2157_));
 sky130_fd_sc_hd__nand2b_1 _5937_ (.A_N(_3501_),
    .B(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__a41oi_1 _5938_ (.A1(_3502_),
    .A2(_3510_),
    .A3(_3518_),
    .A4(_2113_),
    .B1(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__xor2_1 _5939_ (.A(_3494_),
    .B(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__nor2_1 _5940_ (.A(_1824_),
    .B(_2160_),
    .Y(_2161_));
 sky130_fd_sc_hd__mux2i_2 _5941_ (.A0(net519),
    .A1(_1689_),
    .S(_1754_),
    .Y(_2162_));
 sky130_fd_sc_hd__o211a_1 _5942_ (.A1(_3515_),
    .A2(net709),
    .B1(_1902_),
    .C1(_0140_),
    .X(_2163_));
 sky130_fd_sc_hd__a21oi_2 _5943_ (.A1(net276),
    .A2(_2162_),
    .B1(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hd__mux2i_4 _5944_ (.A0(_2021_),
    .A1(_2164_),
    .S(_1921_),
    .Y(_2165_));
 sky130_fd_sc_hd__nor2_1 _5945_ (.A(net932),
    .B(_2003_),
    .Y(_2166_));
 sky130_fd_sc_hd__nor2_1 _5946_ (.A(net267),
    .B(_2010_),
    .Y(_2167_));
 sky130_fd_sc_hd__o21ai_0 _5947_ (.A1(_2166_),
    .A2(_2167_),
    .B1(_1949_),
    .Y(_2168_));
 sky130_fd_sc_hd__o211ai_1 _5948_ (.A1(_1949_),
    .A2(_2165_),
    .B1(_2168_),
    .C1(net171),
    .Y(_2169_));
 sky130_fd_sc_hd__nor2_1 _5949_ (.A(net171),
    .B(_1990_),
    .Y(_2170_));
 sky130_fd_sc_hd__nor2_1 _5950_ (.A(_1921_),
    .B(_1987_),
    .Y(_2171_));
 sky130_fd_sc_hd__a31oi_2 _5951_ (.A1(_1921_),
    .A2(_1997_),
    .A3(_1998_),
    .B1(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand2_1 _5952_ (.A(_2170_),
    .B(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__a21oi_1 _5953_ (.A1(_2169_),
    .A2(_2173_),
    .B1(net266),
    .Y(_2174_));
 sky130_fd_sc_hd__mux2i_2 _5954_ (.A0(_1982_),
    .A1(_1967_),
    .S(net426),
    .Y(_2175_));
 sky130_fd_sc_hd__nor2_1 _5955_ (.A(net431),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__a21oi_1 _5956_ (.A1(_0274_),
    .A2(net424),
    .B1(net170),
    .Y(_2177_));
 sky130_fd_sc_hd__o21ai_2 _5957_ (.A1(net267),
    .A2(_1976_),
    .B1(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__nor2_2 _5958_ (.A(net171),
    .B(net426),
    .Y(_2179_));
 sky130_fd_sc_hd__a21oi_1 _5959_ (.A1(_1970_),
    .A2(_2179_),
    .B1(net24),
    .Y(_2180_));
 sky130_fd_sc_hd__a21oi_1 _5960_ (.A1(net24),
    .A2(_2178_),
    .B1(_2180_),
    .Y(_2181_));
 sky130_fd_sc_hd__o21ai_1 _5961_ (.A1(_2176_),
    .A2(_2181_),
    .B1(_1993_),
    .Y(_2182_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(net177),
    .B(_2182_),
    .Y(_2183_));
 sky130_fd_sc_hd__o32a_1 _5963_ (.A1(net177),
    .A2(_2154_),
    .A3(_2161_),
    .B1(_2174_),
    .B2(_2183_),
    .X(net93));
 sky130_fd_sc_hd__mux2i_2 _5964_ (.A0(_2046_),
    .A1(_2053_),
    .S(net426),
    .Y(_2184_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(net171),
    .B(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__o21ai_0 _5966_ (.A1(_2057_),
    .A2(_2146_),
    .B1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hd__nand2_1 _5967_ (.A(_1949_),
    .B(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hd__nand2_4 _5968_ (.A(net24),
    .B(_1949_),
    .Y(_2188_));
 sky130_fd_sc_hd__nor2_4 _5969_ (.A(_0274_),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__a21oi_1 _5970_ (.A1(net166),
    .A2(net407),
    .B1(net171),
    .Y(_2190_));
 sky130_fd_sc_hd__nand2_1 _5971_ (.A(_2189_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__a21o_1 _5972_ (.A1(_3502_),
    .A2(net279),
    .B1(_3501_),
    .X(_2192_));
 sky130_fd_sc_hd__a21oi_2 _5973_ (.A1(_2192_),
    .A2(_3494_),
    .B1(_3493_),
    .Y(_2193_));
 sky130_fd_sc_hd__xnor2_2 _5974_ (.A(_2193_),
    .B(_3486_),
    .Y(_2194_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_3486_),
    .B(_1820_),
    .Y(_2195_));
 sky130_fd_sc_hd__o211ai_2 _5976_ (.A1(_3489_),
    .A2(_1795_),
    .B1(_2195_),
    .C1(_1956_),
    .Y(_2196_));
 sky130_fd_sc_hd__a221oi_4 _5977_ (.A1(_3485_),
    .A2(net172),
    .B1(_2194_),
    .B2(_1818_),
    .C1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hd__mux2i_4 _5978_ (.A0(net517),
    .A1(_3503_),
    .S(_1754_),
    .Y(_2198_));
 sky130_fd_sc_hd__mux2i_1 _5979_ (.A0(_2162_),
    .A1(_2198_),
    .S(net168),
    .Y(_2199_));
 sky130_fd_sc_hd__mux2_1 _5980_ (.A0(_2066_),
    .A1(_2199_),
    .S(net166),
    .X(_2200_));
 sky130_fd_sc_hd__nand2_1 _5981_ (.A(net267),
    .B(_2032_),
    .Y(_2201_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(net932),
    .B(_2035_),
    .Y(_2202_));
 sky130_fd_sc_hd__nand3_1 _5983_ (.A(_1949_),
    .B(_2201_),
    .C(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hd__o21ai_0 _5984_ (.A1(_1949_),
    .A2(_2200_),
    .B1(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(net267),
    .B(_2049_),
    .Y(_2205_));
 sky130_fd_sc_hd__o21ai_1 _5986_ (.A1(_1702_),
    .A2(_2030_),
    .B1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__a221oi_2 _5987_ (.A1(net171),
    .A2(_2204_),
    .B1(_2206_),
    .B2(_2170_),
    .C1(_2122_),
    .Y(_2207_));
 sky130_fd_sc_hd__a311oi_4 _5988_ (.A1(_2151_),
    .A2(_2187_),
    .A3(_2191_),
    .B1(_2197_),
    .C1(_2207_),
    .Y(net94));
 sky130_fd_sc_hd__inv_1 _5989_ (.A(_3479_),
    .Y(_3475_));
 sky130_fd_sc_hd__mux2i_4 _5990_ (.A0(_2086_),
    .A1(_2079_),
    .S(net267),
    .Y(_2208_));
 sky130_fd_sc_hd__a31oi_1 _5991_ (.A1(net254),
    .A2(net165),
    .A3(net167),
    .B1(net24),
    .Y(_2209_));
 sky130_fd_sc_hd__o21ai_1 _5992_ (.A1(_0274_),
    .A2(_2209_),
    .B1(net465),
    .Y(_2210_));
 sky130_fd_sc_hd__o211ai_4 _5993_ (.A1(net431),
    .A2(_2208_),
    .B1(_2210_),
    .C1(_1949_),
    .Y(_2211_));
 sky130_fd_sc_hd__nor2_1 _5994_ (.A(net166),
    .B(_2107_),
    .Y(_2212_));
 sky130_fd_sc_hd__mux2i_4 _5995_ (.A0(_3479_),
    .A1(net520),
    .S(net265),
    .Y(_2213_));
 sky130_fd_sc_hd__mux2i_4 _5996_ (.A0(_2198_),
    .A1(_2213_),
    .S(net276),
    .Y(_2214_));
 sky130_fd_sc_hd__nor2_1 _5997_ (.A(net427),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__nor2_1 _5998_ (.A(_2212_),
    .B(_2215_),
    .Y(_2216_));
 sky130_fd_sc_hd__nand2_1 _5999_ (.A(net267),
    .B(_2100_),
    .Y(_2217_));
 sky130_fd_sc_hd__nand2_1 _6000_ (.A(net932),
    .B(_2096_),
    .Y(_2218_));
 sky130_fd_sc_hd__nand3_1 _6001_ (.A(_1949_),
    .B(_2217_),
    .C(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__o21ai_0 _6002_ (.A1(_1949_),
    .A2(_2216_),
    .B1(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__mux2i_2 _6003_ (.A0(_2087_),
    .A1(_2099_),
    .S(net166),
    .Y(_2221_));
 sky130_fd_sc_hd__a221oi_2 _6004_ (.A1(net171),
    .A2(_2220_),
    .B1(_2221_),
    .B2(_2170_),
    .C1(_2122_),
    .Y(_2222_));
 sky130_fd_sc_hd__and4_1 _6005_ (.A(_3494_),
    .B(_3502_),
    .C(_3510_),
    .D(_3518_),
    .X(_2223_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(_3524_),
    .B(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hd__nor3_1 _6007_ (.A(net168),
    .B(net501),
    .C(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__a21oi_2 _6008_ (.A1(_3494_),
    .A2(_2158_),
    .B1(_3493_),
    .Y(_2226_));
 sky130_fd_sc_hd__o31ai_2 _6009_ (.A1(_0122_),
    .A2(_0140_),
    .A3(_2224_),
    .B1(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__o21a_1 _6010_ (.A1(_2225_),
    .A2(_2227_),
    .B1(_3486_),
    .X(_2228_));
 sky130_fd_sc_hd__nor2_1 _6011_ (.A(_3485_),
    .B(_2228_),
    .Y(_2229_));
 sky130_fd_sc_hd__xnor2_1 _6012_ (.A(_3478_),
    .B(_2229_),
    .Y(_2230_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_3478_),
    .B(_1820_),
    .Y(_2231_));
 sky130_fd_sc_hd__o211ai_2 _6014_ (.A1(_3481_),
    .A2(_1795_),
    .B1(_2231_),
    .C1(_1956_),
    .Y(_2232_));
 sky130_fd_sc_hd__a221oi_4 _6015_ (.A1(_3477_),
    .A2(net172),
    .B1(_1818_),
    .B2(_2230_),
    .C1(_2232_),
    .Y(_2233_));
 sky130_fd_sc_hd__a211oi_4 _6016_ (.A1(_2151_),
    .A2(_2211_),
    .B1(_2233_),
    .C1(_2222_),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _6017_ (.A(_3471_),
    .Y(_3467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__mux2i_1 _6019_ (.A0(_3471_),
    .A1(net517),
    .S(net466),
    .Y(_2235_));
 sky130_fd_sc_hd__mux2i_2 _6020_ (.A0(_2213_),
    .A1(_2235_),
    .S(net276),
    .Y(_2236_));
 sky130_fd_sc_hd__nand2_1 _6021_ (.A(net166),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__nand3_1 _6022_ (.A(net426),
    .B(_2123_),
    .C(_2124_),
    .Y(_2238_));
 sky130_fd_sc_hd__a32oi_2 _6023_ (.A1(net171),
    .A2(_2237_),
    .A3(_2238_),
    .B1(_1953_),
    .B2(_2179_),
    .Y(_2239_));
 sky130_fd_sc_hd__mux2i_1 _6024_ (.A0(_1924_),
    .A1(_1946_),
    .S(net465),
    .Y(_2240_));
 sky130_fd_sc_hd__mux2i_1 _6025_ (.A0(_2239_),
    .A1(_2240_),
    .S(_1949_),
    .Y(_2241_));
 sky130_fd_sc_hd__nand2_1 _6026_ (.A(net24),
    .B(_3284_),
    .Y(_2242_));
 sky130_fd_sc_hd__nor2_1 _6027_ (.A(net170),
    .B(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__a21oi_1 _6028_ (.A1(_1890_),
    .A2(_1937_),
    .B1(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__o21ai_0 _6029_ (.A1(_1990_),
    .A2(_2244_),
    .B1(net266),
    .Y(_2245_));
 sky130_fd_sc_hd__o21ai_2 _6030_ (.A1(net266),
    .A2(_2241_),
    .B1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__nor3b_2 _6031_ (.A(_1842_),
    .B(net288),
    .C_N(_3478_),
    .Y(_2247_));
 sky130_fd_sc_hd__o21a_1 _6032_ (.A1(_3477_),
    .A2(_2247_),
    .B1(_3470_),
    .X(_2248_));
 sky130_fd_sc_hd__o31ai_1 _6033_ (.A1(_3470_),
    .A2(_3477_),
    .A3(_2247_),
    .B1(_1818_),
    .Y(_2249_));
 sky130_fd_sc_hd__nor2_1 _6034_ (.A(_3473_),
    .B(_1795_),
    .Y(_2250_));
 sky130_fd_sc_hd__a221oi_1 _6035_ (.A1(_3469_),
    .A2(net175),
    .B1(_1820_),
    .B2(_3470_),
    .C1(_2250_),
    .Y(_2251_));
 sky130_fd_sc_hd__o211a_1 _6036_ (.A1(_2248_),
    .A2(_2249_),
    .B1(_1956_),
    .C1(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__a21oi_4 _6037_ (.A1(_1809_),
    .A2(_2246_),
    .B1(_2252_),
    .Y(net96));
 sky130_fd_sc_hd__inv_1 _6038_ (.A(net852),
    .Y(_3459_));
 sky130_fd_sc_hd__nand2_8 _6039_ (.A(_1927_),
    .B(_1990_),
    .Y(_2253_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__mux2i_1 _6041_ (.A0(net855),
    .A1(_3479_),
    .S(_1754_),
    .Y(_2255_));
 sky130_fd_sc_hd__mux2_1 _6042_ (.A0(_2235_),
    .A1(_2255_),
    .S(net168),
    .X(_2256_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(net166),
    .B(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__o21ai_2 _6044_ (.A1(net166),
    .A2(_2164_),
    .B1(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__o2bb2ai_1 _6045_ (.A1_N(net171),
    .A2_N(_2258_),
    .B1(_2146_),
    .B2(_2021_),
    .Y(_2259_));
 sky130_fd_sc_hd__mux2i_2 _6046_ (.A0(_1988_),
    .A1(_2005_),
    .S(net171),
    .Y(_2260_));
 sky130_fd_sc_hd__nand2_2 _6047_ (.A(_1927_),
    .B(_1949_),
    .Y(_2261_));
 sky130_fd_sc_hd__mux2_1 _6048_ (.A0(_0274_),
    .A1(_1977_),
    .S(net170),
    .X(_2262_));
 sky130_fd_sc_hd__nor3_4 _6049_ (.A(net24),
    .B(_1652_),
    .C(_1990_),
    .Y(_2263_));
 sky130_fd_sc_hd__inv_1 _6050_ (.A(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__o221ai_4 _6051_ (.A1(_2188_),
    .A2(_2262_),
    .B1(_2264_),
    .B2(_1972_),
    .C1(net440),
    .Y(_2265_));
 sky130_fd_sc_hd__o221ai_4 _6052_ (.A1(_2253_),
    .A2(_2259_),
    .B1(_2260_),
    .B2(_2261_),
    .C1(_2265_),
    .Y(_2266_));
 sky130_fd_sc_hd__and3_1 _6053_ (.A(_3470_),
    .B(_3478_),
    .C(_3486_),
    .X(_2267_));
 sky130_fd_sc_hd__o21ai_2 _6054_ (.A1(_2227_),
    .A2(_2225_),
    .B1(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__a21o_1 _6055_ (.A1(_3485_),
    .A2(_3478_),
    .B1(_3477_),
    .X(_2269_));
 sky130_fd_sc_hd__a21oi_1 _6056_ (.A1(_3470_),
    .A2(_2269_),
    .B1(_3469_),
    .Y(_2270_));
 sky130_fd_sc_hd__nand2_2 _6057_ (.A(net305),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__xor2_1 _6058_ (.A(_3462_),
    .B(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__a22oi_1 _6059_ (.A1(_3461_),
    .A2(net175),
    .B1(_1820_),
    .B2(_3462_),
    .Y(_2273_));
 sky130_fd_sc_hd__o21ai_0 _6060_ (.A1(_3465_),
    .A2(_1795_),
    .B1(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__a211oi_2 _6061_ (.A1(_2272_),
    .A2(_1818_),
    .B1(_2274_),
    .C1(_1809_),
    .Y(_2275_));
 sky130_fd_sc_hd__a21oi_2 _6062_ (.A1(_1809_),
    .A2(_2266_),
    .B1(_2275_),
    .Y(net97));
 sky130_fd_sc_hd__mux2i_1 _6063_ (.A0(_3455_),
    .A1(_3471_),
    .S(_1754_),
    .Y(_2276_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(_2255_),
    .A1(_2276_),
    .S(net168),
    .X(_2277_));
 sky130_fd_sc_hd__nor2_1 _6065_ (.A(net166),
    .B(_2199_),
    .Y(_2278_));
 sky130_fd_sc_hd__a21oi_1 _6066_ (.A1(net166),
    .A2(_2277_),
    .B1(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__o22a_1 _6067_ (.A1(_2066_),
    .A2(_2146_),
    .B1(_2279_),
    .B2(_1652_),
    .X(_2280_));
 sky130_fd_sc_hd__nand2b_1 _6068_ (.A_N(_2033_),
    .B(net171),
    .Y(_2281_));
 sky130_fd_sc_hd__o211ai_1 _6069_ (.A1(net170),
    .A2(_2051_),
    .B1(_2281_),
    .C1(_1949_),
    .Y(_2282_));
 sky130_fd_sc_hd__o21ai_1 _6070_ (.A1(_1949_),
    .A2(_2280_),
    .B1(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__nor2_1 _6071_ (.A(_1652_),
    .B(net265),
    .Y(_2284_));
 sky130_fd_sc_hd__o22ai_2 _6072_ (.A1(_1652_),
    .A2(_2055_),
    .B1(_2284_),
    .B2(_0274_),
    .Y(_2285_));
 sky130_fd_sc_hd__a21oi_1 _6073_ (.A1(_1954_),
    .A2(_2053_),
    .B1(_2188_),
    .Y(_2286_));
 sky130_fd_sc_hd__a22oi_4 _6074_ (.A1(_2056_),
    .A2(_2263_),
    .B1(_2285_),
    .B2(_2286_),
    .Y(_2287_));
 sky130_fd_sc_hd__nand2_1 _6075_ (.A(net266),
    .B(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__o21ai_4 _6076_ (.A1(net266),
    .A2(_2283_),
    .B1(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__o21a_1 _6077_ (.A1(_3469_),
    .A2(_2248_),
    .B1(_3462_),
    .X(_2290_));
 sky130_fd_sc_hd__nor3_1 _6078_ (.A(_3454_),
    .B(_3461_),
    .C(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__o21ai_1 _6079_ (.A1(_3461_),
    .A2(_2290_),
    .B1(_3454_),
    .Y(_2292_));
 sky130_fd_sc_hd__nor3b_2 _6080_ (.A(_1824_),
    .B(_2291_),
    .C_N(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2_1 _6081_ (.A(_3454_),
    .B(_1820_),
    .Y(_2294_));
 sky130_fd_sc_hd__o21ai_0 _6082_ (.A1(_3457_),
    .A2(_1795_),
    .B1(_2294_),
    .Y(_2295_));
 sky130_fd_sc_hd__a2111oi_4 _6083_ (.A1(_3453_),
    .A2(net175),
    .B1(_2295_),
    .C1(_2293_),
    .D1(_1809_),
    .Y(_2296_));
 sky130_fd_sc_hd__a21oi_4 _6084_ (.A1(_1809_),
    .A2(_2289_),
    .B1(_2296_),
    .Y(net67));
 sky130_fd_sc_hd__a21o_1 _6085_ (.A1(_3462_),
    .A2(_2271_),
    .B1(_3461_),
    .X(_2297_));
 sky130_fd_sc_hd__a21oi_2 _6086_ (.A1(_3454_),
    .A2(_2297_),
    .B1(_3453_),
    .Y(_2298_));
 sky130_fd_sc_hd__xnor2_1 _6087_ (.A(_2298_),
    .B(_3446_),
    .Y(_2299_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_3446_),
    .B(_1820_),
    .Y(_2300_));
 sky130_fd_sc_hd__o21ai_1 _6089_ (.A1(_3449_),
    .A2(_1795_),
    .B1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__a221oi_4 _6090_ (.A1(_3445_),
    .A2(net175),
    .B1(_2299_),
    .B2(_1818_),
    .C1(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__nand2_1 _6091_ (.A(net170),
    .B(net165),
    .Y(_2303_));
 sky130_fd_sc_hd__a21oi_1 _6092_ (.A1(_0274_),
    .A2(_2303_),
    .B1(_2188_),
    .Y(_2304_));
 sky130_fd_sc_hd__nand2_1 _6093_ (.A(_1954_),
    .B(_2079_),
    .Y(_2305_));
 sky130_fd_sc_hd__a221o_1 _6094_ (.A1(_2082_),
    .A2(_2263_),
    .B1(_2304_),
    .B2(_2305_),
    .C1(_1927_),
    .X(_2306_));
 sky130_fd_sc_hd__mux2i_2 _6095_ (.A0(_3447_),
    .A1(net855),
    .S(_1754_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux2_1 _6096_ (.A0(_2276_),
    .A1(_2307_),
    .S(net168),
    .X(_2308_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(net165),
    .B(_2308_),
    .Y(_2309_));
 sky130_fd_sc_hd__o21ai_2 _6098_ (.A1(net165),
    .A2(_2214_),
    .B1(_2309_),
    .Y(_2310_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(net171),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__nand2b_1 _6100_ (.A_N(_2107_),
    .B(_2179_),
    .Y(_2312_));
 sky130_fd_sc_hd__mux2i_1 _6101_ (.A0(_2088_),
    .A1(_2101_),
    .S(net171),
    .Y(_2313_));
 sky130_fd_sc_hd__a32oi_1 _6102_ (.A1(_1955_),
    .A2(_2311_),
    .A3(_2312_),
    .B1(_1995_),
    .B2(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__a21oi_2 _6103_ (.A1(_2306_),
    .A2(_2314_),
    .B1(_1956_),
    .Y(_2315_));
 sky130_fd_sc_hd__a21oi_2 _6104_ (.A1(_2302_),
    .A2(_1956_),
    .B1(_2315_),
    .Y(net68));
 sky130_fd_sc_hd__nor2_1 _6105_ (.A(net170),
    .B(_2148_),
    .Y(_2316_));
 sky130_fd_sc_hd__nor2_1 _6106_ (.A(net431),
    .B(_2133_),
    .Y(_2317_));
 sky130_fd_sc_hd__mux2i_2 _6107_ (.A0(_3439_),
    .A1(_3455_),
    .S(net466),
    .Y(_2318_));
 sky130_fd_sc_hd__mux2i_2 _6108_ (.A0(_2307_),
    .A1(_2318_),
    .S(net276),
    .Y(_2319_));
 sky130_fd_sc_hd__mux2i_4 _6109_ (.A0(_2236_),
    .A1(_2319_),
    .S(_1921_),
    .Y(_2320_));
 sky130_fd_sc_hd__mux2i_2 _6110_ (.A0(_2126_),
    .A1(_2320_),
    .S(net170),
    .Y(_2321_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_1990_),
    .B(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__o311ai_4 _6112_ (.A1(_1990_),
    .A2(_2316_),
    .A3(_2317_),
    .B1(_2322_),
    .C1(_1927_),
    .Y(_2323_));
 sky130_fd_sc_hd__nand2_1 _6113_ (.A(_1932_),
    .B(_1954_),
    .Y(_2324_));
 sky130_fd_sc_hd__o21ai_1 _6114_ (.A1(_1954_),
    .A2(_2242_),
    .B1(_2324_),
    .Y(_2325_));
 sky130_fd_sc_hd__a21oi_2 _6115_ (.A1(_1993_),
    .A2(_2325_),
    .B1(_1956_),
    .Y(_2326_));
 sky130_fd_sc_hd__nand2b_1 _6116_ (.A_N(_3453_),
    .B(_2292_),
    .Y(_2327_));
 sky130_fd_sc_hd__a21oi_1 _6117_ (.A1(_3446_),
    .A2(_2327_),
    .B1(_3445_),
    .Y(_2328_));
 sky130_fd_sc_hd__xnor2_1 _6118_ (.A(_3438_),
    .B(_2328_),
    .Y(_2329_));
 sky130_fd_sc_hd__nand2_1 _6119_ (.A(_3438_),
    .B(_1820_),
    .Y(_2330_));
 sky130_fd_sc_hd__o211ai_2 _6120_ (.A1(_3441_),
    .A2(_1795_),
    .B1(_2330_),
    .C1(_1956_),
    .Y(_2331_));
 sky130_fd_sc_hd__a221oi_4 _6121_ (.A1(_3437_),
    .A2(net175),
    .B1(_2329_),
    .B2(_1818_),
    .C1(_2331_),
    .Y(_2332_));
 sky130_fd_sc_hd__a21oi_4 _6122_ (.A1(_2323_),
    .A2(_2326_),
    .B1(_2332_),
    .Y(net69));
 sky130_fd_sc_hd__a21o_1 _6123_ (.A1(_3454_),
    .A2(_3461_),
    .B1(_3453_),
    .X(_2333_));
 sky130_fd_sc_hd__a21o_1 _6124_ (.A1(_3446_),
    .A2(_2333_),
    .B1(_3445_),
    .X(_2334_));
 sky130_fd_sc_hd__a21oi_4 _6125_ (.A1(_3438_),
    .A2(_2334_),
    .B1(_3437_),
    .Y(_2335_));
 sky130_fd_sc_hd__a21o_2 _6126_ (.A1(_2270_),
    .A2(_2268_),
    .B1(_1846_),
    .X(_2336_));
 sky130_fd_sc_hd__and2_1 _6127_ (.A(_2335_),
    .B(net304),
    .X(_2337_));
 sky130_fd_sc_hd__xnor2_1 _6128_ (.A(_3430_),
    .B(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__nand2_1 _6129_ (.A(_1818_),
    .B(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__nor2_1 _6130_ (.A(_3433_),
    .B(_1795_),
    .Y(_2340_));
 sky130_fd_sc_hd__a21oi_1 _6131_ (.A1(_3430_),
    .A2(_1820_),
    .B1(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__a21oi_1 _6132_ (.A1(_3429_),
    .A2(net175),
    .B1(_1809_),
    .Y(_2342_));
 sky130_fd_sc_hd__o21ai_2 _6133_ (.A1(_2303_),
    .A2(_1976_),
    .B1(_2304_),
    .Y(_2343_));
 sky130_fd_sc_hd__nand3_1 _6134_ (.A(net166),
    .B(_1970_),
    .C(_2263_),
    .Y(_2344_));
 sky130_fd_sc_hd__nor2_1 _6135_ (.A(net171),
    .B(_2175_),
    .Y(_2345_));
 sky130_fd_sc_hd__a211oi_1 _6136_ (.A1(net171),
    .A2(_2172_),
    .B1(_2345_),
    .C1(_2261_),
    .Y(_2346_));
 sky130_fd_sc_hd__mux2i_2 _6137_ (.A0(_3435_),
    .A1(_3451_),
    .S(net466),
    .Y(_2347_));
 sky130_fd_sc_hd__mux2i_4 _6138_ (.A0(_3427_),
    .A1(_3443_),
    .S(_1754_),
    .Y(_2348_));
 sky130_fd_sc_hd__mux2i_4 _6139_ (.A0(_2347_),
    .A1(_2348_),
    .S(net259),
    .Y(_2349_));
 sky130_fd_sc_hd__mux2i_2 _6140_ (.A0(_2256_),
    .A1(_2349_),
    .S(net166),
    .Y(_2350_));
 sky130_fd_sc_hd__nand2_1 _6141_ (.A(net171),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__o21a_1 _6142_ (.A1(net171),
    .A2(_2165_),
    .B1(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__nor2_1 _6143_ (.A(_2253_),
    .B(_2352_),
    .Y(_2353_));
 sky130_fd_sc_hd__a311o_4 _6144_ (.A1(net266),
    .A2(_2343_),
    .A3(_2344_),
    .B1(_2346_),
    .C1(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__a32oi_4 _6145_ (.A1(_2339_),
    .A2(_2341_),
    .A3(_2342_),
    .B1(_2354_),
    .B2(_1809_),
    .Y(net70));
 sky130_fd_sc_hd__nand2_1 _6146_ (.A(net431),
    .B(_2184_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(net171),
    .B(_2206_),
    .Y(_2356_));
 sky130_fd_sc_hd__and3_1 _6148_ (.A(_1995_),
    .B(_2355_),
    .C(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__nor3_1 _6149_ (.A(_0140_),
    .B(net265),
    .C(_2303_),
    .Y(_2358_));
 sky130_fd_sc_hd__nand2_1 _6150_ (.A(_0371_),
    .B(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__o211ai_1 _6151_ (.A1(_3284_),
    .A2(_2358_),
    .B1(_2359_),
    .C1(_2143_),
    .Y(_2360_));
 sky130_fd_sc_hd__o311a_1 _6152_ (.A1(net421),
    .A2(_2057_),
    .A3(_2264_),
    .B1(_2360_),
    .C1(net266),
    .X(_2361_));
 sky130_fd_sc_hd__mux2i_4 _6153_ (.A0(_3419_),
    .A1(_3435_),
    .S(_1754_),
    .Y(_2362_));
 sky130_fd_sc_hd__mux2i_4 _6154_ (.A0(_2348_),
    .A1(_2362_),
    .S(net258),
    .Y(_2363_));
 sky130_fd_sc_hd__mux2i_2 _6155_ (.A0(_2277_),
    .A1(_2363_),
    .S(net166),
    .Y(_2364_));
 sky130_fd_sc_hd__mux2i_2 _6156_ (.A0(_2200_),
    .A1(_2364_),
    .S(net171),
    .Y(_2365_));
 sky130_fd_sc_hd__nor2_1 _6157_ (.A(_2253_),
    .B(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__nor2_1 _6158_ (.A(_1852_),
    .B(_1854_),
    .Y(_2367_));
 sky130_fd_sc_hd__o21ai_0 _6159_ (.A1(_1849_),
    .A2(_2367_),
    .B1(_3430_),
    .Y(_2368_));
 sky130_fd_sc_hd__nand2b_1 _6160_ (.A_N(_3429_),
    .B(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__xnor2_1 _6161_ (.A(_3422_),
    .B(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hd__a22oi_1 _6162_ (.A1(_3421_),
    .A2(net175),
    .B1(_1820_),
    .B2(_3422_),
    .Y(_2371_));
 sky130_fd_sc_hd__o221ai_1 _6163_ (.A1(_3425_),
    .A2(_1795_),
    .B1(_1824_),
    .B2(_2370_),
    .C1(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__nand2_2 _6164_ (.A(_1956_),
    .B(_2372_),
    .Y(_2373_));
 sky130_fd_sc_hd__o41ai_4 _6165_ (.A1(_1956_),
    .A2(_2357_),
    .A3(_2361_),
    .A4(_2366_),
    .B1(_2373_),
    .Y(net71));
 sky130_fd_sc_hd__inv_1 _6166_ (.A(_3414_),
    .Y(_2374_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_3422_),
    .B(_3430_),
    .Y(_2375_));
 sky130_fd_sc_hd__a21oi_1 _6168_ (.A1(_3422_),
    .A2(_3429_),
    .B1(_3421_),
    .Y(_2376_));
 sky130_fd_sc_hd__o21ai_0 _6169_ (.A1(_2337_),
    .A2(_2375_),
    .B1(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__xnor2_1 _6170_ (.A(_2374_),
    .B(_2377_),
    .Y(_2378_));
 sky130_fd_sc_hd__nand2_1 _6171_ (.A(_1818_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__nor2_1 _6172_ (.A(_3417_),
    .B(_1795_),
    .Y(_2380_));
 sky130_fd_sc_hd__a21oi_1 _6173_ (.A1(_3414_),
    .A2(_1820_),
    .B1(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__a21oi_1 _6174_ (.A1(_3413_),
    .A2(net175),
    .B1(_1809_),
    .Y(_2382_));
 sky130_fd_sc_hd__nand2_1 _6175_ (.A(net431),
    .B(_2208_),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_1 _6176_ (.A(net170),
    .B(_2221_),
    .Y(_2384_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(_2261_),
    .B(_2144_),
    .Y(_2385_));
 sky130_fd_sc_hd__a31oi_1 _6178_ (.A1(net166),
    .A2(_2080_),
    .A3(_2263_),
    .B1(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__a31oi_1 _6179_ (.A1(_1927_),
    .A2(_2383_),
    .A3(_2384_),
    .B1(_2386_),
    .Y(_2387_));
 sky130_fd_sc_hd__mux2i_2 _6180_ (.A0(_2107_),
    .A1(_2214_),
    .S(net165),
    .Y(_2388_));
 sky130_fd_sc_hd__mux2i_4 _6181_ (.A0(_3411_),
    .A1(_3427_),
    .S(net466),
    .Y(_2389_));
 sky130_fd_sc_hd__mux2i_4 _6182_ (.A0(_2362_),
    .A1(_2389_),
    .S(net258),
    .Y(_2390_));
 sky130_fd_sc_hd__mux2_1 _6183_ (.A0(_2308_),
    .A1(_2390_),
    .S(net165),
    .X(_2391_));
 sky130_fd_sc_hd__mux2i_4 _6184_ (.A0(_2388_),
    .A1(_2391_),
    .S(net170),
    .Y(_2392_));
 sky130_fd_sc_hd__o21ai_0 _6185_ (.A1(_2253_),
    .A2(_2392_),
    .B1(net176),
    .Y(_2393_));
 sky130_fd_sc_hd__nor2_2 _6186_ (.A(_2387_),
    .B(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__a31oi_4 _6187_ (.A1(_2379_),
    .A2(_2381_),
    .A3(_2382_),
    .B1(_2394_),
    .Y(net72));
 sky130_fd_sc_hd__nor2_1 _6188_ (.A(_3409_),
    .B(_1795_),
    .Y(_2395_));
 sky130_fd_sc_hd__a21oi_1 _6189_ (.A1(_3406_),
    .A2(_1820_),
    .B1(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__a21oi_1 _6190_ (.A1(_3405_),
    .A2(_1803_),
    .B1(net177),
    .Y(_2397_));
 sky130_fd_sc_hd__o21a_1 _6191_ (.A1(_1849_),
    .A2(_1856_),
    .B1(_1864_),
    .X(_2398_));
 sky130_fd_sc_hd__a21oi_2 _6192_ (.A1(_2398_),
    .A2(_3414_),
    .B1(_3413_),
    .Y(_2399_));
 sky130_fd_sc_hd__xnor2_1 _6193_ (.A(_2399_),
    .B(_3406_),
    .Y(_2400_));
 sky130_fd_sc_hd__nand2_1 _6194_ (.A(_1818_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__mux2_1 _6195_ (.A0(_2307_),
    .A1(_2318_),
    .S(net168),
    .X(_2402_));
 sky130_fd_sc_hd__mux2i_4 _6196_ (.A0(_3403_),
    .A1(_3419_),
    .S(net466),
    .Y(_2403_));
 sky130_fd_sc_hd__mux2i_1 _6197_ (.A0(_2389_),
    .A1(_2403_),
    .S(net169),
    .Y(_2404_));
 sky130_fd_sc_hd__mux2i_1 _6198_ (.A0(_2402_),
    .A1(_2404_),
    .S(_1921_),
    .Y(_2405_));
 sky130_fd_sc_hd__nor2_1 _6199_ (.A(net431),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__a31o_1 _6200_ (.A1(net465),
    .A2(_2237_),
    .A3(_2238_),
    .B1(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__nor2_4 _6201_ (.A(_1927_),
    .B(_1949_),
    .Y(_2408_));
 sky130_fd_sc_hd__and3_1 _6202_ (.A(_1953_),
    .B(_1954_),
    .C(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__nor2_2 _6203_ (.A(_1995_),
    .B(_2189_),
    .Y(_2410_));
 sky130_fd_sc_hd__a21oi_1 _6204_ (.A1(_1927_),
    .A2(_1947_),
    .B1(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__a2111oi_2 _6205_ (.A1(_1955_),
    .A2(_2407_),
    .B1(_2409_),
    .C1(_2411_),
    .D1(_1956_),
    .Y(_2412_));
 sky130_fd_sc_hd__a31oi_4 _6206_ (.A1(_2396_),
    .A2(_2401_),
    .A3(_2397_),
    .B1(_2412_),
    .Y(net73));
 sky130_fd_sc_hd__mux2i_4 _6207_ (.A0(_3395_),
    .A1(_3411_),
    .S(net466),
    .Y(_2413_));
 sky130_fd_sc_hd__mux2i_4 _6208_ (.A0(_2403_),
    .A1(_2413_),
    .S(net261),
    .Y(_2414_));
 sky130_fd_sc_hd__mux2i_1 _6209_ (.A0(_2349_),
    .A1(_2414_),
    .S(net166),
    .Y(_2415_));
 sky130_fd_sc_hd__nand2_1 _6210_ (.A(net170),
    .B(_2415_),
    .Y(_2416_));
 sky130_fd_sc_hd__o211ai_2 _6211_ (.A1(net170),
    .A2(_2258_),
    .B1(_2416_),
    .C1(_1955_),
    .Y(_2417_));
 sky130_fd_sc_hd__a21oi_4 _6212_ (.A1(_0274_),
    .A2(net440),
    .B1(_2188_),
    .Y(_2418_));
 sky130_fd_sc_hd__o21ai_0 _6213_ (.A1(net170),
    .A2(_1977_),
    .B1(_1927_),
    .Y(_2419_));
 sky130_fd_sc_hd__nand2_1 _6214_ (.A(_1954_),
    .B(_2408_),
    .Y(_2420_));
 sky130_fd_sc_hd__o21ai_0 _6215_ (.A1(_2021_),
    .A2(_2420_),
    .B1(net177),
    .Y(_2421_));
 sky130_fd_sc_hd__a21oi_1 _6216_ (.A1(_2418_),
    .A2(_2419_),
    .B1(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__nor3_2 _6217_ (.A(net24),
    .B(net437),
    .C(_1990_),
    .Y(_2423_));
 sky130_fd_sc_hd__nor3_1 _6218_ (.A(net465),
    .B(_1988_),
    .C(_2410_),
    .Y(_2424_));
 sky130_fd_sc_hd__a31oi_2 _6219_ (.A1(net431),
    .A2(_1971_),
    .A3(_2423_),
    .B1(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__nand2_1 _6220_ (.A(_3470_),
    .B(_2269_),
    .Y(_2426_));
 sky130_fd_sc_hd__nand4_4 _6221_ (.A(_3406_),
    .B(_3414_),
    .C(_3422_),
    .D(_3430_),
    .Y(_2427_));
 sky130_fd_sc_hd__nor2_1 _6222_ (.A(_1846_),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__a21boi_2 _6223_ (.A1(_2268_),
    .A2(_2426_),
    .B1_N(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__nand2_1 _6224_ (.A(_3469_),
    .B(_2428_),
    .Y(_2430_));
 sky130_fd_sc_hd__o21ai_0 _6225_ (.A1(_2335_),
    .A2(_2427_),
    .B1(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__o21bai_1 _6226_ (.A1(_2374_),
    .A2(_2376_),
    .B1_N(_3413_),
    .Y(_2432_));
 sky130_fd_sc_hd__a21oi_2 _6227_ (.A1(_3406_),
    .A2(_2432_),
    .B1(_3405_),
    .Y(_2433_));
 sky130_fd_sc_hd__nor3b_2 _6228_ (.A(_2431_),
    .B(_2429_),
    .C_N(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__xnor2_1 _6229_ (.A(_3398_),
    .B(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__nand2_1 _6230_ (.A(_3398_),
    .B(_1820_),
    .Y(_2436_));
 sky130_fd_sc_hd__o211ai_2 _6231_ (.A1(_3401_),
    .A2(_1795_),
    .B1(_2436_),
    .C1(_1956_),
    .Y(_2437_));
 sky130_fd_sc_hd__a221oi_4 _6232_ (.A1(_3397_),
    .A2(_1803_),
    .B1(_2435_),
    .B2(_1818_),
    .C1(_2437_),
    .Y(_2438_));
 sky130_fd_sc_hd__a31oi_4 _6233_ (.A1(_2417_),
    .A2(_2422_),
    .A3(_2425_),
    .B1(_2438_),
    .Y(net74));
 sky130_fd_sc_hd__inv_1 _6234_ (.A(_1031_),
    .Y(_3387_));
 sky130_fd_sc_hd__and2_0 _6235_ (.A(net431),
    .B(_2059_),
    .X(_2439_));
 sky130_fd_sc_hd__o21ai_1 _6236_ (.A1(net266),
    .A2(_2439_),
    .B1(_2418_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor2_2 _6237_ (.A(net465),
    .B(_2410_),
    .Y(_2441_));
 sky130_fd_sc_hd__nand3_1 _6238_ (.A(net431),
    .B(_2056_),
    .C(_2423_),
    .Y(_2442_));
 sky130_fd_sc_hd__o211ai_1 _6239_ (.A1(_2066_),
    .A2(_2420_),
    .B1(_2442_),
    .C1(net177),
    .Y(_2443_));
 sky130_fd_sc_hd__a21oi_1 _6240_ (.A1(_2051_),
    .A2(_2441_),
    .B1(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__nand2_1 _6241_ (.A(net431),
    .B(_2279_),
    .Y(_2445_));
 sky130_fd_sc_hd__mux2_1 _6242_ (.A0(_1031_),
    .A1(_3407_),
    .S(net466),
    .X(_2446_));
 sky130_fd_sc_hd__mux2i_2 _6243_ (.A0(_2413_),
    .A1(_2446_),
    .S(net169),
    .Y(_2447_));
 sky130_fd_sc_hd__mux2i_1 _6244_ (.A0(_2363_),
    .A1(_2447_),
    .S(net165),
    .Y(_2448_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(net170),
    .B(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__nand3_1 _6246_ (.A(_1955_),
    .B(_2445_),
    .C(_2449_),
    .Y(_2450_));
 sky130_fd_sc_hd__inv_1 _6247_ (.A(_3406_),
    .Y(_2451_));
 sky130_fd_sc_hd__o21bai_1 _6248_ (.A1(_2451_),
    .A2(_2399_),
    .B1_N(_3405_),
    .Y(_2452_));
 sky130_fd_sc_hd__a21oi_1 _6249_ (.A1(_2452_),
    .A2(_3398_),
    .B1(_3397_),
    .Y(_2453_));
 sky130_fd_sc_hd__xnor2_1 _6250_ (.A(_3390_),
    .B(_2453_),
    .Y(_2454_));
 sky130_fd_sc_hd__nand2_1 _6251_ (.A(_3390_),
    .B(_1820_),
    .Y(_2455_));
 sky130_fd_sc_hd__o211ai_2 _6252_ (.A1(_3393_),
    .A2(_1795_),
    .B1(_2455_),
    .C1(_1956_),
    .Y(_2456_));
 sky130_fd_sc_hd__a221oi_4 _6253_ (.A1(_3389_),
    .A2(net174),
    .B1(_2454_),
    .B2(_1818_),
    .C1(_2456_),
    .Y(_2457_));
 sky130_fd_sc_hd__a31oi_4 _6254_ (.A1(_2440_),
    .A2(_2444_),
    .A3(_2450_),
    .B1(_2457_),
    .Y(net75));
 sky130_fd_sc_hd__inv_1 _6255_ (.A(_3383_),
    .Y(_3379_));
 sky130_fd_sc_hd__nand2_1 _6256_ (.A(_3390_),
    .B(_3398_),
    .Y(_2458_));
 sky130_fd_sc_hd__a21oi_1 _6257_ (.A1(_3390_),
    .A2(_3397_),
    .B1(_3389_),
    .Y(_2459_));
 sky130_fd_sc_hd__o21ai_1 _6258_ (.A1(_2458_),
    .A2(_2434_),
    .B1(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__xnor2_1 _6259_ (.A(_1867_),
    .B(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__nand2_1 _6260_ (.A(_3382_),
    .B(_1820_),
    .Y(_2462_));
 sky130_fd_sc_hd__o211ai_2 _6261_ (.A1(_3385_),
    .A2(_1795_),
    .B1(_2462_),
    .C1(_1956_),
    .Y(_2463_));
 sky130_fd_sc_hd__a221oi_4 _6262_ (.A1(_3381_),
    .A2(net174),
    .B1(_2461_),
    .B2(_1818_),
    .C1(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__mux2i_1 _6263_ (.A0(_1031_),
    .A1(_3407_),
    .S(net265),
    .Y(_2465_));
 sky130_fd_sc_hd__mux2i_1 _6264_ (.A0(_3383_),
    .A1(_3399_),
    .S(net466),
    .Y(_2466_));
 sky130_fd_sc_hd__mux2i_2 _6265_ (.A0(_2465_),
    .A1(_2466_),
    .S(net261),
    .Y(_2467_));
 sky130_fd_sc_hd__nand2_1 _6266_ (.A(net267),
    .B(_2390_),
    .Y(_2468_));
 sky130_fd_sc_hd__o21ai_2 _6267_ (.A1(net267),
    .A2(_2467_),
    .B1(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__mux2i_1 _6268_ (.A0(_2310_),
    .A1(_2469_),
    .S(net170),
    .Y(_2470_));
 sky130_fd_sc_hd__a221oi_1 _6269_ (.A1(_2084_),
    .A2(_2418_),
    .B1(_2423_),
    .B2(_2082_),
    .C1(_2441_),
    .Y(_2471_));
 sky130_fd_sc_hd__nor2_1 _6270_ (.A(net431),
    .B(_2088_),
    .Y(_2472_));
 sky130_fd_sc_hd__a21oi_4 _6271_ (.A1(net439),
    .A2(_2189_),
    .B1(_1956_),
    .Y(_2473_));
 sky130_fd_sc_hd__o21a_1 _6272_ (.A1(_2107_),
    .A2(_2420_),
    .B1(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__o221a_1 _6273_ (.A1(_2253_),
    .A2(_2470_),
    .B1(_2471_),
    .B2(_2472_),
    .C1(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__nor2_1 _6274_ (.A(_2464_),
    .B(_2475_),
    .Y(net76));
 sky130_fd_sc_hd__inv_1 _6275_ (.A(_3375_),
    .Y(_3371_));
 sky130_fd_sc_hd__mux2i_2 _6276_ (.A0(_3375_),
    .A1(_1031_),
    .S(net466),
    .Y(_2476_));
 sky130_fd_sc_hd__mux2_1 _6277_ (.A0(_2466_),
    .A1(_2476_),
    .S(net169),
    .X(_2477_));
 sky130_fd_sc_hd__nor2_1 _6278_ (.A(net421),
    .B(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__nor2_1 _6279_ (.A(_1921_),
    .B(_2404_),
    .Y(_2479_));
 sky130_fd_sc_hd__nor3_1 _6280_ (.A(_2253_),
    .B(_2478_),
    .C(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(_2126_),
    .B(_2408_),
    .Y(_2481_));
 sky130_fd_sc_hd__o21ai_0 _6282_ (.A1(_2148_),
    .A2(_2410_),
    .B1(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__o21ai_0 _6283_ (.A1(_2480_),
    .A2(_2482_),
    .B1(net170),
    .Y(_2483_));
 sky130_fd_sc_hd__nand2_1 _6284_ (.A(net267),
    .B(_1935_),
    .Y(_2484_));
 sky130_fd_sc_hd__o21ai_0 _6285_ (.A1(net267),
    .A2(_1932_),
    .B1(net465),
    .Y(_2485_));
 sky130_fd_sc_hd__a21oi_1 _6286_ (.A1(_2484_),
    .A2(_2485_),
    .B1(_2144_),
    .Y(_2486_));
 sky130_fd_sc_hd__o31ai_1 _6287_ (.A1(_2145_),
    .A2(_2261_),
    .A3(_2146_),
    .B1(_2473_),
    .Y(_2487_));
 sky130_fd_sc_hd__a311oi_1 _6288_ (.A1(net431),
    .A2(_1955_),
    .A3(_2320_),
    .B1(_2486_),
    .C1(_2487_),
    .Y(_2488_));
 sky130_fd_sc_hd__nand2_1 _6289_ (.A(_1866_),
    .B(_1872_),
    .Y(_2489_));
 sky130_fd_sc_hd__xnor2_2 _6290_ (.A(_1874_),
    .B(_2489_),
    .Y(_2490_));
 sky130_fd_sc_hd__nand2_1 _6291_ (.A(_3374_),
    .B(_1820_),
    .Y(_2491_));
 sky130_fd_sc_hd__o211ai_2 _6292_ (.A1(_3377_),
    .A2(_1795_),
    .B1(_2491_),
    .C1(_1956_),
    .Y(_2492_));
 sky130_fd_sc_hd__a221oi_4 _6293_ (.A1(_3373_),
    .A2(net174),
    .B1(_2490_),
    .B2(_1818_),
    .C1(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__a21oi_4 _6294_ (.A1(_2483_),
    .A2(_2488_),
    .B1(_2493_),
    .Y(net78));
 sky130_fd_sc_hd__inv_1 _6295_ (.A(_3367_),
    .Y(_3363_));
 sky130_fd_sc_hd__nand2b_1 _6296_ (.A_N(_2175_),
    .B(_2441_),
    .Y(_2494_));
 sky130_fd_sc_hd__nand2_1 _6297_ (.A(net166),
    .B(_2423_),
    .Y(_2495_));
 sky130_fd_sc_hd__nor2b_1 _6298_ (.A(_2495_),
    .B_N(_1970_),
    .Y(_2496_));
 sky130_fd_sc_hd__nor2_1 _6299_ (.A(_2253_),
    .B(_2350_),
    .Y(_2497_));
 sky130_fd_sc_hd__o21ai_0 _6300_ (.A1(_2496_),
    .A2(_2497_),
    .B1(net431),
    .Y(_2498_));
 sky130_fd_sc_hd__nand2b_1 _6301_ (.A_N(_2178_),
    .B(_2418_),
    .Y(_2499_));
 sky130_fd_sc_hd__and3_1 _6302_ (.A(_2473_),
    .B(_2498_),
    .C(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__mux2i_2 _6303_ (.A0(_3367_),
    .A1(_3383_),
    .S(_1754_),
    .Y(_2501_));
 sky130_fd_sc_hd__mux2i_4 _6304_ (.A0(_2476_),
    .A1(_2501_),
    .S(net251),
    .Y(_2502_));
 sky130_fd_sc_hd__nor2_1 _6305_ (.A(net166),
    .B(_2414_),
    .Y(_2503_));
 sky130_fd_sc_hd__a211oi_2 _6306_ (.A1(net166),
    .A2(_2502_),
    .B1(_2503_),
    .C1(_2253_),
    .Y(_2504_));
 sky130_fd_sc_hd__a21o_1 _6307_ (.A1(_2165_),
    .A2(_2408_),
    .B1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__nand2_1 _6308_ (.A(net171),
    .B(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__nand2_1 _6309_ (.A(_3366_),
    .B(_1820_),
    .Y(_2507_));
 sky130_fd_sc_hd__o211ai_2 _6310_ (.A1(_3369_),
    .A2(_1795_),
    .B1(_2507_),
    .C1(_1956_),
    .Y(_2508_));
 sky130_fd_sc_hd__a21oi_4 _6311_ (.A1(_3365_),
    .A2(net173),
    .B1(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand4_1 _6312_ (.A(_3390_),
    .B(_3374_),
    .C(_3382_),
    .D(_3398_),
    .Y(_2510_));
 sky130_fd_sc_hd__o21bai_1 _6313_ (.A1(_1867_),
    .A2(_2459_),
    .B1_N(_3381_),
    .Y(_2511_));
 sky130_fd_sc_hd__a21oi_1 _6314_ (.A1(_3374_),
    .A2(_2511_),
    .B1(_3373_),
    .Y(_2512_));
 sky130_fd_sc_hd__o21ai_1 _6315_ (.A1(_2433_),
    .A2(_2510_),
    .B1(_2512_),
    .Y(_2513_));
 sky130_fd_sc_hd__a211oi_2 _6316_ (.A1(_2336_),
    .A2(_2335_),
    .B1(_2427_),
    .C1(_2510_),
    .Y(_2514_));
 sky130_fd_sc_hd__nor3_1 _6317_ (.A(_3366_),
    .B(_2513_),
    .C(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__o21ai_0 _6318_ (.A1(_2513_),
    .A2(_2514_),
    .B1(_3366_),
    .Y(_2516_));
 sky130_fd_sc_hd__or3b_4 _6319_ (.A(_1824_),
    .B(_2515_),
    .C_N(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__a32oi_4 _6320_ (.A1(_2494_),
    .A2(_2500_),
    .A3(_2506_),
    .B1(_2517_),
    .B2(_2509_),
    .Y(net79));
 sky130_fd_sc_hd__inv_1 _6321_ (.A(_3359_),
    .Y(_3355_));
 sky130_fd_sc_hd__a31oi_1 _6322_ (.A1(_1927_),
    .A2(net166),
    .A3(net407),
    .B1(_2144_),
    .Y(_2518_));
 sky130_fd_sc_hd__o21ai_1 _6323_ (.A1(_2441_),
    .A2(_2518_),
    .B1(_2184_),
    .Y(_2519_));
 sky130_fd_sc_hd__o21ai_0 _6324_ (.A1(net437),
    .A2(_2190_),
    .B1(_2189_),
    .Y(_2520_));
 sky130_fd_sc_hd__o21ai_0 _6325_ (.A1(_2057_),
    .A2(_2146_),
    .B1(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__nor3_1 _6326_ (.A(net171),
    .B(_2253_),
    .C(_2364_),
    .Y(_2522_));
 sky130_fd_sc_hd__a21oi_1 _6327_ (.A1(_2385_),
    .A2(_2521_),
    .B1(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__nor2_1 _6328_ (.A(net165),
    .B(_2447_),
    .Y(_2524_));
 sky130_fd_sc_hd__mux2i_1 _6329_ (.A0(_3359_),
    .A1(_3375_),
    .S(_1754_),
    .Y(_2525_));
 sky130_fd_sc_hd__mux2_1 _6330_ (.A0(_2501_),
    .A1(_2525_),
    .S(net169),
    .X(_2526_));
 sky130_fd_sc_hd__nor2_1 _6331_ (.A(net421),
    .B(_2526_),
    .Y(_2527_));
 sky130_fd_sc_hd__nor3_2 _6332_ (.A(net441),
    .B(_2524_),
    .C(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__nor2_1 _6333_ (.A(_1927_),
    .B(_2200_),
    .Y(_2529_));
 sky130_fd_sc_hd__o211ai_2 _6334_ (.A1(_2528_),
    .A2(_2529_),
    .B1(net171),
    .C1(_1990_),
    .Y(_2530_));
 sky130_fd_sc_hd__a21oi_1 _6335_ (.A1(_2489_),
    .A2(_3374_),
    .B1(_3373_),
    .Y(_2531_));
 sky130_fd_sc_hd__nor2b_1 _6336_ (.A(_2531_),
    .B_N(_3366_),
    .Y(_2532_));
 sky130_fd_sc_hd__nor2_1 _6337_ (.A(_3365_),
    .B(_2532_),
    .Y(_2533_));
 sky130_fd_sc_hd__xnor2_1 _6338_ (.A(_2533_),
    .B(_3358_),
    .Y(_2534_));
 sky130_fd_sc_hd__nand2_1 _6339_ (.A(_3358_),
    .B(_1820_),
    .Y(_2535_));
 sky130_fd_sc_hd__o211ai_2 _6340_ (.A1(_3361_),
    .A2(_1795_),
    .B1(_2535_),
    .C1(_1956_),
    .Y(_2536_));
 sky130_fd_sc_hd__a221oi_4 _6341_ (.A1(_3357_),
    .A2(net173),
    .B1(_2534_),
    .B2(_1818_),
    .C1(_2536_),
    .Y(_2537_));
 sky130_fd_sc_hd__a41oi_4 _6342_ (.A1(net177),
    .A2(_2519_),
    .A3(_2523_),
    .A4(_2530_),
    .B1(_2537_),
    .Y(net80));
 sky130_fd_sc_hd__inv_1 _6343_ (.A(_3351_),
    .Y(_3347_));
 sky130_fd_sc_hd__nor2_1 _6344_ (.A(_3353_),
    .B(_1795_),
    .Y(_2538_));
 sky130_fd_sc_hd__a21oi_1 _6345_ (.A1(_3350_),
    .A2(_1820_),
    .B1(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__a21oi_1 _6346_ (.A1(_3349_),
    .A2(net174),
    .B1(net176),
    .Y(_2540_));
 sky130_fd_sc_hd__a21o_1 _6347_ (.A1(_3366_),
    .A2(_2513_),
    .B1(_3365_),
    .X(_2541_));
 sky130_fd_sc_hd__a21oi_2 _6348_ (.A1(_3358_),
    .A2(_2541_),
    .B1(_3357_),
    .Y(_2542_));
 sky130_fd_sc_hd__nand2_1 _6349_ (.A(_3358_),
    .B(_3366_),
    .Y(_2543_));
 sky130_fd_sc_hd__a2111o_1 _6350_ (.A1(_2336_),
    .A2(_2335_),
    .B1(_2427_),
    .C1(_2510_),
    .D1(_2543_),
    .X(_2544_));
 sky130_fd_sc_hd__a21oi_1 _6351_ (.A1(_2542_),
    .A2(_2544_),
    .B1(_3350_),
    .Y(_2545_));
 sky130_fd_sc_hd__and3_1 _6352_ (.A(_3350_),
    .B(_2542_),
    .C(_2544_),
    .X(_2546_));
 sky130_fd_sc_hd__o21ai_1 _6353_ (.A1(_2545_),
    .A2(_2546_),
    .B1(_1818_),
    .Y(_2547_));
 sky130_fd_sc_hd__a31oi_1 _6354_ (.A1(net166),
    .A2(_2080_),
    .A3(_2423_),
    .B1(net170),
    .Y(_2548_));
 sky130_fd_sc_hd__o21ai_0 _6355_ (.A1(_2261_),
    .A2(_2548_),
    .B1(_2144_),
    .Y(_2549_));
 sky130_fd_sc_hd__o21a_1 _6356_ (.A1(net431),
    .A2(_2208_),
    .B1(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__mux2i_2 _6357_ (.A0(_3351_),
    .A1(_3367_),
    .S(net265),
    .Y(_2551_));
 sky130_fd_sc_hd__mux2i_2 _6358_ (.A0(_2525_),
    .A1(_2551_),
    .S(net250),
    .Y(_2552_));
 sky130_fd_sc_hd__mux2i_2 _6359_ (.A0(_2467_),
    .A1(_2552_),
    .S(net165),
    .Y(_2553_));
 sky130_fd_sc_hd__mux2i_1 _6360_ (.A0(_2391_),
    .A1(_2553_),
    .S(net170),
    .Y(_2554_));
 sky130_fd_sc_hd__nand2_1 _6361_ (.A(net170),
    .B(_2408_),
    .Y(_2555_));
 sky130_fd_sc_hd__o221ai_1 _6362_ (.A1(_2253_),
    .A2(_2554_),
    .B1(_2555_),
    .B2(_2216_),
    .C1(_2473_),
    .Y(_2556_));
 sky130_fd_sc_hd__nor2_1 _6363_ (.A(_2550_),
    .B(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__a31oi_4 _6364_ (.A1(_2539_),
    .A2(_2547_),
    .A3(_2540_),
    .B1(_2557_),
    .Y(net81));
 sky130_fd_sc_hd__inv_1 _6365_ (.A(_3343_),
    .Y(_3339_));
 sky130_fd_sc_hd__nor2_1 _6366_ (.A(_1890_),
    .B(_2405_),
    .Y(_2558_));
 sky130_fd_sc_hd__mux2i_2 _6367_ (.A0(_3343_),
    .A1(_3359_),
    .S(net466),
    .Y(_2559_));
 sky130_fd_sc_hd__mux2i_2 _6368_ (.A0(_2551_),
    .A1(_2559_),
    .S(net263),
    .Y(_2560_));
 sky130_fd_sc_hd__nor2_1 _6369_ (.A(net165),
    .B(_2477_),
    .Y(_2561_));
 sky130_fd_sc_hd__a211oi_1 _6370_ (.A1(net165),
    .A2(_2560_),
    .B1(_2561_),
    .C1(_1652_),
    .Y(_2562_));
 sky130_fd_sc_hd__o21ai_0 _6371_ (.A1(_2558_),
    .A2(_2562_),
    .B1(_1990_),
    .Y(_2563_));
 sky130_fd_sc_hd__o21ai_0 _6372_ (.A1(_1990_),
    .A2(_2244_),
    .B1(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__o21ai_0 _6373_ (.A1(_1949_),
    .A2(_2239_),
    .B1(net266),
    .Y(_2565_));
 sky130_fd_sc_hd__o21ai_2 _6374_ (.A1(net266),
    .A2(_2564_),
    .B1(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__a21oi_1 _6375_ (.A1(_1873_),
    .A2(_1877_),
    .B1(_3349_),
    .Y(_2567_));
 sky130_fd_sc_hd__xnor2_1 _6376_ (.A(_3342_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__nand2_1 _6377_ (.A(_3341_),
    .B(net173),
    .Y(_2569_));
 sky130_fd_sc_hd__o211ai_2 _6378_ (.A1(_3345_),
    .A2(_1795_),
    .B1(_2569_),
    .C1(_1956_),
    .Y(_2570_));
 sky130_fd_sc_hd__a221oi_4 _6379_ (.A1(_3342_),
    .A2(_1820_),
    .B1(_1818_),
    .B2(_2568_),
    .C1(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__a21oi_4 _6380_ (.A1(_2473_),
    .A2(_2566_),
    .B1(_2571_),
    .Y(net82));
 sky130_fd_sc_hd__inv_1 _6381_ (.A(_3335_),
    .Y(_3331_));
 sky130_fd_sc_hd__nand2_1 _6382_ (.A(_2259_),
    .B(_2408_),
    .Y(_2572_));
 sky130_fd_sc_hd__a21oi_1 _6383_ (.A1(_1927_),
    .A2(net170),
    .B1(_0274_),
    .Y(_2573_));
 sky130_fd_sc_hd__nor3_1 _6384_ (.A(net443),
    .B(net465),
    .C(_1977_),
    .Y(_2574_));
 sky130_fd_sc_hd__o21ai_1 _6385_ (.A1(_2573_),
    .A2(_2574_),
    .B1(_2143_),
    .Y(_2575_));
 sky130_fd_sc_hd__nand2_1 _6386_ (.A(net267),
    .B(_2502_),
    .Y(_2576_));
 sky130_fd_sc_hd__mux2i_1 _6387_ (.A0(_3335_),
    .A1(_3351_),
    .S(_1754_),
    .Y(_2577_));
 sky130_fd_sc_hd__mux2i_2 _6388_ (.A0(_2559_),
    .A1(_2577_),
    .S(net249),
    .Y(_2578_));
 sky130_fd_sc_hd__nand2_1 _6389_ (.A(net165),
    .B(_2578_),
    .Y(_2579_));
 sky130_fd_sc_hd__nor2_1 _6390_ (.A(net170),
    .B(_2415_),
    .Y(_2580_));
 sky130_fd_sc_hd__a31oi_1 _6391_ (.A1(net170),
    .A2(_2576_),
    .A3(_2579_),
    .B1(_2580_),
    .Y(_2581_));
 sky130_fd_sc_hd__o22ai_1 _6392_ (.A1(_1972_),
    .A2(_2264_),
    .B1(_2581_),
    .B2(_1949_),
    .Y(_2582_));
 sky130_fd_sc_hd__nand2_1 _6393_ (.A(_1927_),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__inv_1 _6394_ (.A(_3334_),
    .Y(_2584_));
 sky130_fd_sc_hd__nand2_1 _6395_ (.A(_3342_),
    .B(_3350_),
    .Y(_2585_));
 sky130_fd_sc_hd__nor2_1 _6396_ (.A(_2543_),
    .B(_2585_),
    .Y(_2586_));
 sky130_fd_sc_hd__o21ai_1 _6397_ (.A1(_2513_),
    .A2(_2514_),
    .B1(_2586_),
    .Y(_2587_));
 sky130_fd_sc_hd__a21o_1 _6398_ (.A1(_3358_),
    .A2(_3365_),
    .B1(_3357_),
    .X(_2588_));
 sky130_fd_sc_hd__a21o_1 _6399_ (.A1(_3350_),
    .A2(_2588_),
    .B1(_3349_),
    .X(_2589_));
 sky130_fd_sc_hd__a21oi_1 _6400_ (.A1(_3342_),
    .A2(_2589_),
    .B1(_3341_),
    .Y(_2590_));
 sky130_fd_sc_hd__nand3_1 _6401_ (.A(_2584_),
    .B(_2587_),
    .C(_2590_),
    .Y(_2591_));
 sky130_fd_sc_hd__a21o_1 _6402_ (.A1(_2587_),
    .A2(_2590_),
    .B1(_2584_),
    .X(_2592_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(_3334_),
    .B(_1820_),
    .Y(_2593_));
 sky130_fd_sc_hd__a21oi_1 _6404_ (.A1(_3333_),
    .A2(net173),
    .B1(net176),
    .Y(_2594_));
 sky130_fd_sc_hd__o211ai_2 _6405_ (.A1(_3337_),
    .A2(_1795_),
    .B1(_2593_),
    .C1(_2594_),
    .Y(_2595_));
 sky130_fd_sc_hd__a31oi_4 _6406_ (.A1(_1818_),
    .A2(_2591_),
    .A3(_2592_),
    .B1(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__a41oi_4 _6407_ (.A1(net177),
    .A2(_2572_),
    .A3(_2575_),
    .A4(_2583_),
    .B1(_2596_),
    .Y(net83));
 sky130_fd_sc_hd__inv_1 _6408_ (.A(_0621_),
    .Y(_3323_));
 sky130_fd_sc_hd__mux2i_1 _6409_ (.A0(_0621_),
    .A1(_3343_),
    .S(_1754_),
    .Y(_2597_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(_2577_),
    .A1(_2597_),
    .S(net247),
    .X(_2598_));
 sky130_fd_sc_hd__mux2i_1 _6411_ (.A0(_2526_),
    .A1(_2598_),
    .S(net165),
    .Y(_2599_));
 sky130_fd_sc_hd__mux2_1 _6412_ (.A0(_2448_),
    .A1(_2599_),
    .S(net170),
    .X(_2600_));
 sky130_fd_sc_hd__o21ai_0 _6413_ (.A1(_1949_),
    .A2(_2600_),
    .B1(_2287_),
    .Y(_2601_));
 sky130_fd_sc_hd__nand2_1 _6414_ (.A(_1927_),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__nand2b_1 _6415_ (.A_N(_2280_),
    .B(_2408_),
    .Y(_2603_));
 sky130_fd_sc_hd__nor3_1 _6416_ (.A(_3326_),
    .B(_1878_),
    .C(_1880_),
    .Y(_2604_));
 sky130_fd_sc_hd__o21ai_0 _6417_ (.A1(_1878_),
    .A2(_1880_),
    .B1(_3326_),
    .Y(_2605_));
 sky130_fd_sc_hd__nand2b_4 _6418_ (.A_N(_2604_),
    .B(_2605_),
    .Y(_2606_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(_3326_),
    .B(_1820_),
    .Y(_2607_));
 sky130_fd_sc_hd__o211ai_2 _6420_ (.A1(_3329_),
    .A2(_1795_),
    .B1(_2607_),
    .C1(_1956_),
    .Y(_2608_));
 sky130_fd_sc_hd__a221oi_4 _6421_ (.A1(_3325_),
    .A2(net174),
    .B1(_2606_),
    .B2(_1818_),
    .C1(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__a31oi_4 _6422_ (.A1(_2473_),
    .A2(_2602_),
    .A3(_2603_),
    .B1(_2609_),
    .Y(net84));
 sky130_fd_sc_hd__nand2_1 _6423_ (.A(_3318_),
    .B(_1820_),
    .Y(_2610_));
 sky130_fd_sc_hd__a21oi_1 _6424_ (.A1(_3317_),
    .A2(net173),
    .B1(net176),
    .Y(_2611_));
 sky130_fd_sc_hd__o211ai_1 _6425_ (.A1(_3321_),
    .A2(_1795_),
    .B1(_2610_),
    .C1(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__a21oi_1 _6426_ (.A1(_3342_),
    .A2(_3349_),
    .B1(_3341_),
    .Y(_2613_));
 sky130_fd_sc_hd__nor2_1 _6427_ (.A(_2584_),
    .B(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__nand3_1 _6428_ (.A(_3342_),
    .B(_3334_),
    .C(_3350_),
    .Y(_2615_));
 sky130_fd_sc_hd__a21oi_1 _6429_ (.A1(_2542_),
    .A2(_2544_),
    .B1(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__o31ai_1 _6430_ (.A1(_3333_),
    .A2(_2614_),
    .A3(_2616_),
    .B1(_3326_),
    .Y(_2617_));
 sky130_fd_sc_hd__nor2_1 _6431_ (.A(_3318_),
    .B(_3325_),
    .Y(_2618_));
 sky130_fd_sc_hd__a211oi_4 _6432_ (.A1(_2544_),
    .A2(_2542_),
    .B1(_2615_),
    .C1(_1881_),
    .Y(_2619_));
 sky130_fd_sc_hd__nor2_1 _6433_ (.A(_3333_),
    .B(_2614_),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _6434_ (.A(_3318_),
    .B(_3325_),
    .Y(_2621_));
 sky130_fd_sc_hd__o21ai_1 _6435_ (.A1(_1881_),
    .A2(_2620_),
    .B1(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__or3_1 _6436_ (.A(_1824_),
    .B(_2619_),
    .C(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__a21oi_2 _6437_ (.A1(_2617_),
    .A2(_2618_),
    .B1(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__mux2i_1 _6438_ (.A0(_3319_),
    .A1(_3335_),
    .S(net265),
    .Y(_2625_));
 sky130_fd_sc_hd__mux2i_1 _6439_ (.A0(_2597_),
    .A1(_2625_),
    .S(net263),
    .Y(_2626_));
 sky130_fd_sc_hd__nand2_1 _6440_ (.A(net165),
    .B(_2626_),
    .Y(_2627_));
 sky130_fd_sc_hd__nand2_1 _6441_ (.A(net267),
    .B(_2552_),
    .Y(_2628_));
 sky130_fd_sc_hd__and3_1 _6442_ (.A(net170),
    .B(_2627_),
    .C(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__a21oi_1 _6443_ (.A1(net465),
    .A2(_2469_),
    .B1(_2629_),
    .Y(_2630_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(net170),
    .B(_2308_),
    .Y(_2631_));
 sky130_fd_sc_hd__o21ai_0 _6445_ (.A1(net170),
    .A2(_2107_),
    .B1(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__nor2_1 _6446_ (.A(_2214_),
    .B(_2555_),
    .Y(_2633_));
 sky130_fd_sc_hd__a31oi_1 _6447_ (.A1(_1927_),
    .A2(_2080_),
    .A3(_2263_),
    .B1(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__nor2_1 _6448_ (.A(net165),
    .B(_2634_),
    .Y(_2635_));
 sky130_fd_sc_hd__a31oi_2 _6449_ (.A1(net165),
    .A2(_2408_),
    .A3(_2632_),
    .B1(_2635_),
    .Y(_2636_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_1927_),
    .B(_1954_),
    .Y(_2637_));
 sky130_fd_sc_hd__nor3_1 _6451_ (.A(_1990_),
    .B(_2079_),
    .C(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__a21oi_1 _6452_ (.A1(_2189_),
    .A2(_2637_),
    .B1(_2638_),
    .Y(_2639_));
 sky130_fd_sc_hd__o2111ai_4 _6453_ (.A1(_2253_),
    .A2(_2630_),
    .B1(_2636_),
    .C1(_2639_),
    .D1(net176),
    .Y(_2640_));
 sky130_fd_sc_hd__o21a_4 _6454_ (.A1(_2612_),
    .A2(_2624_),
    .B1(_2640_),
    .X(net85));
 sky130_fd_sc_hd__inv_1 _6455_ (.A(_3311_),
    .Y(_3307_));
 sky130_fd_sc_hd__nor2_1 _6456_ (.A(_3313_),
    .B(_1795_),
    .Y(_2641_));
 sky130_fd_sc_hd__a21oi_1 _6457_ (.A1(_3310_),
    .A2(_1820_),
    .B1(_2641_),
    .Y(_2642_));
 sky130_fd_sc_hd__a21oi_1 _6458_ (.A1(_3309_),
    .A2(net173),
    .B1(net176),
    .Y(_2643_));
 sky130_fd_sc_hd__xor2_1 _6459_ (.A(_3310_),
    .B(_1883_),
    .X(_2644_));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(_1818_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__mux2i_1 _6461_ (.A0(_3311_),
    .A1(_0621_),
    .S(net265),
    .Y(_2646_));
 sky130_fd_sc_hd__nor2_1 _6462_ (.A(_0140_),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__nor2_1 _6463_ (.A(net263),
    .B(_2625_),
    .Y(_2648_));
 sky130_fd_sc_hd__nor2_1 _6464_ (.A(_2647_),
    .B(_2648_),
    .Y(_2649_));
 sky130_fd_sc_hd__nor2_1 _6465_ (.A(net165),
    .B(_2560_),
    .Y(_2650_));
 sky130_fd_sc_hd__a21oi_1 _6466_ (.A1(net165),
    .A2(_2649_),
    .B1(_2650_),
    .Y(_2651_));
 sky130_fd_sc_hd__o22ai_2 _6467_ (.A1(_2145_),
    .A2(_2495_),
    .B1(_2651_),
    .B2(_2253_),
    .Y(_2652_));
 sky130_fd_sc_hd__nand2_1 _6468_ (.A(net442),
    .B(_1990_),
    .Y(_2653_));
 sky130_fd_sc_hd__nor2_1 _6469_ (.A(_2321_),
    .B(_2653_),
    .Y(_2654_));
 sky130_fd_sc_hd__mux2i_1 _6470_ (.A0(_2145_),
    .A1(_0274_),
    .S(_2637_),
    .Y(_2655_));
 sky130_fd_sc_hd__a221o_1 _6471_ (.A1(net465),
    .A2(_2480_),
    .B1(_2655_),
    .B2(_2143_),
    .C1(_1956_),
    .X(_2656_));
 sky130_fd_sc_hd__a211oi_4 _6472_ (.A1(net170),
    .A2(_2652_),
    .B1(_2654_),
    .C1(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__a31oi_4 _6473_ (.A1(_2642_),
    .A2(_2645_),
    .A3(_2643_),
    .B1(_2657_),
    .Y(net86));
 sky130_fd_sc_hd__inv_1 _6474_ (.A(_3303_),
    .Y(_3299_));
 sky130_fd_sc_hd__nand3b_1 _6475_ (.A_N(_3302_),
    .B(_3310_),
    .C(_1818_),
    .Y(_2658_));
 sky130_fd_sc_hd__nand3b_1 _6476_ (.A_N(_3309_),
    .B(_1818_),
    .C(_3302_),
    .Y(_2659_));
 sky130_fd_sc_hd__nor3_2 _6477_ (.A(_3317_),
    .B(_2619_),
    .C(_2622_),
    .Y(_2660_));
 sky130_fd_sc_hd__mux2i_2 _6478_ (.A0(_2658_),
    .A1(_2659_),
    .S(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__nor2_1 _6479_ (.A(_3310_),
    .B(_3309_),
    .Y(_2662_));
 sky130_fd_sc_hd__mux2i_1 _6480_ (.A0(_3309_),
    .A1(_2662_),
    .S(_3302_),
    .Y(_2663_));
 sky130_fd_sc_hd__a21oi_1 _6481_ (.A1(_3301_),
    .A2(net173),
    .B1(net176),
    .Y(_2664_));
 sky130_fd_sc_hd__nor2_1 _6482_ (.A(_3305_),
    .B(_1795_),
    .Y(_2665_));
 sky130_fd_sc_hd__a21oi_1 _6483_ (.A1(_3302_),
    .A2(_1820_),
    .B1(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__o211ai_2 _6484_ (.A1(_1824_),
    .A2(_2663_),
    .B1(_2664_),
    .C1(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__mux2i_1 _6485_ (.A0(_2496_),
    .A1(_2504_),
    .S(net431),
    .Y(_2668_));
 sky130_fd_sc_hd__o21ai_0 _6486_ (.A1(net265),
    .A2(_2637_),
    .B1(_0274_),
    .Y(_2669_));
 sky130_fd_sc_hd__o311ai_0 _6487_ (.A1(net265),
    .A2(_1974_),
    .A3(_2637_),
    .B1(_2669_),
    .C1(_2143_),
    .Y(_2670_));
 sky130_fd_sc_hd__nand2_1 _6488_ (.A(net267),
    .B(_2578_),
    .Y(_2671_));
 sky130_fd_sc_hd__mux2i_1 _6489_ (.A0(_3303_),
    .A1(_3319_),
    .S(net265),
    .Y(_2672_));
 sky130_fd_sc_hd__nand2_1 _6490_ (.A(net252),
    .B(_2672_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_0140_),
    .B(_2646_),
    .Y(_2674_));
 sky130_fd_sc_hd__nand3_1 _6492_ (.A(net165),
    .B(_2673_),
    .C(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__nand4_1 _6493_ (.A(net170),
    .B(_1955_),
    .C(_2671_),
    .D(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__nand3_1 _6494_ (.A(net176),
    .B(_2670_),
    .C(_2676_),
    .Y(_2677_));
 sky130_fd_sc_hd__a21oi_1 _6495_ (.A1(_2352_),
    .A2(_2408_),
    .B1(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__nand2_2 _6496_ (.A(_2668_),
    .B(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__o21ai_4 _6497_ (.A1(_2667_),
    .A2(_2661_),
    .B1(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__inv_1 _6498_ (.A(_2680_),
    .Y(net87));
 sky130_fd_sc_hd__inv_1 _6499_ (.A(_0371_),
    .Y(_3291_));
 sky130_fd_sc_hd__a21oi_1 _6500_ (.A1(_1990_),
    .A2(_2365_),
    .B1(_2418_),
    .Y(_2681_));
 sky130_fd_sc_hd__a21oi_1 _6501_ (.A1(_1927_),
    .A2(_2360_),
    .B1(_2681_),
    .Y(_2682_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_2524_),
    .B(_2527_),
    .Y(_2683_));
 sky130_fd_sc_hd__nand2_1 _6503_ (.A(_1652_),
    .B(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand2_1 _6504_ (.A(_0140_),
    .B(_2672_),
    .Y(_2685_));
 sky130_fd_sc_hd__mux2i_1 _6505_ (.A0(_0371_),
    .A1(_3311_),
    .S(net265),
    .Y(_2686_));
 sky130_fd_sc_hd__nand2_1 _6506_ (.A(net263),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__nor2_1 _6507_ (.A(net165),
    .B(_2598_),
    .Y(_2688_));
 sky130_fd_sc_hd__a311o_1 _6508_ (.A1(net165),
    .A2(_2685_),
    .A3(_2687_),
    .B1(_2688_),
    .C1(_1652_),
    .X(_2689_));
 sky130_fd_sc_hd__a21oi_1 _6509_ (.A1(_2684_),
    .A2(_2689_),
    .B1(_2253_),
    .Y(_2690_));
 sky130_fd_sc_hd__nor3_1 _6510_ (.A(net431),
    .B(_2057_),
    .C(_2495_),
    .Y(_2691_));
 sky130_fd_sc_hd__or4_2 _6511_ (.A(_1956_),
    .B(_2682_),
    .C(_2690_),
    .D(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__xnor2_1 _6512_ (.A(_1885_),
    .B(_3294_),
    .Y(_2693_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(_3294_),
    .B(_1820_),
    .Y(_2694_));
 sky130_fd_sc_hd__o21ai_0 _6514_ (.A1(_3297_),
    .A2(_1795_),
    .B1(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__a211oi_1 _6515_ (.A1(_3293_),
    .A2(net174),
    .B1(_2695_),
    .C1(net176),
    .Y(_2696_));
 sky130_fd_sc_hd__o21ai_1 _6516_ (.A1(_1824_),
    .A2(_2693_),
    .B1(_2696_),
    .Y(_2697_));
 sky130_fd_sc_hd__and2_4 _6517_ (.A(_2692_),
    .B(_2697_),
    .X(net89));
 sky130_fd_sc_hd__a21o_1 _6518_ (.A1(_3310_),
    .A2(_3317_),
    .B1(_3309_),
    .X(_2698_));
 sky130_fd_sc_hd__a21oi_1 _6519_ (.A1(_3302_),
    .A2(_2698_),
    .B1(_3301_),
    .Y(_2699_));
 sky130_fd_sc_hd__nand3b_1 _6520_ (.A_N(_3293_),
    .B(_2699_),
    .C(_3286_),
    .Y(_2700_));
 sky130_fd_sc_hd__nor3_2 _6521_ (.A(_2619_),
    .B(_2622_),
    .C(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__nand2_1 _6522_ (.A(_3302_),
    .B(_3310_),
    .Y(_2702_));
 sky130_fd_sc_hd__nand2_1 _6523_ (.A(_2702_),
    .B(_2699_),
    .Y(_2703_));
 sky130_fd_sc_hd__a21o_1 _6524_ (.A1(_3294_),
    .A2(_2703_),
    .B1(_3293_),
    .X(_2704_));
 sky130_fd_sc_hd__nor2b_1 _6525_ (.A(_2699_),
    .B_N(_3294_),
    .Y(_2705_));
 sky130_fd_sc_hd__nor3_1 _6526_ (.A(_3286_),
    .B(_3293_),
    .C(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__a21oi_1 _6527_ (.A1(_3286_),
    .A2(_2704_),
    .B1(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__nor3b_1 _6528_ (.A(_2702_),
    .B(_3286_),
    .C_N(_3294_),
    .Y(_2708_));
 sky130_fd_sc_hd__o21a_1 _6529_ (.A1(_2619_),
    .A2(_2622_),
    .B1(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__nor3_1 _6530_ (.A(_2701_),
    .B(_2707_),
    .C(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(_1824_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_1 _6532_ (.A(_3286_),
    .B(_1820_),
    .Y(_2712_));
 sky130_fd_sc_hd__a21oi_1 _6533_ (.A1(_3285_),
    .A2(net174),
    .B1(net176),
    .Y(_2713_));
 sky130_fd_sc_hd__o211ai_1 _6534_ (.A1(_3289_),
    .A2(_1795_),
    .B1(_2712_),
    .C1(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__mux2i_1 _6535_ (.A0(_0274_),
    .A1(_3303_),
    .S(net265),
    .Y(_2715_));
 sky130_fd_sc_hd__mux2i_1 _6536_ (.A0(_2686_),
    .A1(_2715_),
    .S(net256),
    .Y(_2716_));
 sky130_fd_sc_hd__mux2i_1 _6537_ (.A0(_2626_),
    .A1(_2716_),
    .S(net165),
    .Y(_2717_));
 sky130_fd_sc_hd__mux2i_2 _6538_ (.A0(_2553_),
    .A1(_2717_),
    .S(net170),
    .Y(_2718_));
 sky130_fd_sc_hd__o41ai_1 _6539_ (.A1(_0140_),
    .A2(_1652_),
    .A3(net265),
    .A4(_2495_),
    .B1(_2188_),
    .Y(_2719_));
 sky130_fd_sc_hd__a21oi_1 _6540_ (.A1(_3284_),
    .A2(_2719_),
    .B1(_1956_),
    .Y(_2720_));
 sky130_fd_sc_hd__o221ai_4 _6541_ (.A1(_2392_),
    .A2(_2653_),
    .B1(_2718_),
    .B2(_2253_),
    .C1(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__o21a_2 _6542_ (.A1(_2714_),
    .A2(_2711_),
    .B1(_2721_),
    .X(net90));
 sky130_fd_sc_hd__or2_4 _6543_ (.A(net31),
    .B(net30),
    .X(_2722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__a311oi_4 _6545_ (.A1(_0035_),
    .A2(_0037_),
    .A3(_0041_),
    .B1(_0130_),
    .C1(net202),
    .Y(_2724_));
 sky130_fd_sc_hd__nor2b_4 _6546_ (.A(_2724_),
    .B_N(net32),
    .Y(_2725_));
 sky130_fd_sc_hd__nand3b_4 _6547_ (.A_N(net2),
    .B(_2725_),
    .C(net3),
    .Y(_2726_));
 sky130_fd_sc_hd__nor2_8 _6548_ (.A(_2722_),
    .B(_2726_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2b_4 _6549_ (.A_N(net30),
    .B(net31),
    .Y(_2727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__nor2_4 _6551_ (.A(net32),
    .B(_2724_),
    .Y(_2729_));
 sky130_fd_sc_hd__nor2_2 _6552_ (.A(net3),
    .B(net2),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_4 _6553_ (.A(_2729_),
    .B(_2730_),
    .Y(_2731_));
 sky130_fd_sc_hd__nor2_8 _6554_ (.A(_2727_),
    .B(_2731_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand2_8 _6555_ (.A(net31),
    .B(net30),
    .Y(_2732_));
 sky130_fd_sc_hd__nand3b_4 _6556_ (.A_N(net3),
    .B(net2),
    .C(_2729_),
    .Y(_2733_));
 sky130_fd_sc_hd__nor2_8 _6557_ (.A(_2732_),
    .B(_2733_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor2_8 _6558_ (.A(_2727_),
    .B(_2733_),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2b_4 _6559_ (.A_N(net31),
    .B(net30),
    .Y(_2734_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__nor2_8 _6561_ (.A(_2733_),
    .B(_2734_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand3b_4 _6562_ (.A_N(net2),
    .B(_2729_),
    .C(net3),
    .Y(_2736_));
 sky130_fd_sc_hd__nor2_8 _6563_ (.A(_2732_),
    .B(_2736_),
    .Y(_0009_));
 sky130_fd_sc_hd__nor2_8 _6564_ (.A(_2722_),
    .B(_2733_),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_8 _6565_ (.A(_2727_),
    .B(_2736_),
    .Y(_0008_));
 sky130_fd_sc_hd__nor2_8 _6566_ (.A(_2734_),
    .B(_2736_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_8 _6567_ (.A(_2725_),
    .B(_2730_),
    .Y(_2737_));
 sky130_fd_sc_hd__nor2_8 _6568_ (.A(_2732_),
    .B(_2737_),
    .Y(_0028_));
 sky130_fd_sc_hd__nor2_8 _6569_ (.A(_2722_),
    .B(_2736_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor2_8 _6570_ (.A(_2727_),
    .B(_2737_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_8 _6571_ (.A(_2734_),
    .B(_2737_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand3b_4 _6572_ (.A_N(net3),
    .B(net2),
    .C(_2725_),
    .Y(_2738_));
 sky130_fd_sc_hd__nor2_8 _6573_ (.A(_2732_),
    .B(_2738_),
    .Y(_0005_));
 sky130_fd_sc_hd__nor2_8 _6574_ (.A(_2722_),
    .B(_2737_),
    .Y(_0025_));
 sky130_fd_sc_hd__nor2_8 _6575_ (.A(_2727_),
    .B(_2738_),
    .Y(_0004_));
 sky130_fd_sc_hd__nor2_8 _6576_ (.A(_2734_),
    .B(_2738_),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_8 _6577_ (.A(_2731_),
    .B(_2732_),
    .Y(_0024_));
 sky130_fd_sc_hd__nor2_8 _6578_ (.A(_2722_),
    .B(_2738_),
    .Y(_0002_));
 sky130_fd_sc_hd__nor2_8 _6579_ (.A(_2731_),
    .B(_2734_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand3_4 _6580_ (.A(net3),
    .B(net2),
    .C(_2725_),
    .Y(_2739_));
 sky130_fd_sc_hd__nor2_8 _6581_ (.A(_2732_),
    .B(_2739_),
    .Y(_0023_));
 sky130_fd_sc_hd__nor2_8 _6582_ (.A(_2727_),
    .B(_2739_),
    .Y(_0022_));
 sky130_fd_sc_hd__nor2_8 _6583_ (.A(_2734_),
    .B(_2739_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand3_4 _6584_ (.A(net3),
    .B(net2),
    .C(_2729_),
    .Y(_2740_));
 sky130_fd_sc_hd__nor2_8 _6585_ (.A(_2734_),
    .B(_2740_),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_8 _6586_ (.A(_2722_),
    .B(_2739_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_8 _6587_ (.A(_2727_),
    .B(_2740_),
    .Y(_0017_));
 sky130_fd_sc_hd__nor2_8 _6588_ (.A(_2732_),
    .B(_2740_),
    .Y(_0018_));
 sky130_fd_sc_hd__nor2_8 _6589_ (.A(_2722_),
    .B(_2740_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_8 _6590_ (.A(_2726_),
    .B(_2732_),
    .Y(_0014_));
 sky130_fd_sc_hd__nor2_8 _6591_ (.A(_2726_),
    .B(_2734_),
    .Y(_0012_));
 sky130_fd_sc_hd__nor2_8 _6592_ (.A(_2726_),
    .B(_2727_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkinv_16 _6593_ (.A(net65),
    .Y(_0031_));
 sky130_fd_sc_hd__or3_4 _6594_ (.A(net28),
    .B(_0126_),
    .C(_0129_),
    .X(_2741_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__nand3_4 _6596_ (.A(_0120_),
    .B(_0913_),
    .C(_2741_),
    .Y(_2743_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__nand2_1 _6599_ (.A(net100),
    .B(_2743_),
    .Y(_2746_));
 sky130_fd_sc_hd__o21ai_0 _6600_ (.A1(net502),
    .A2(_2743_),
    .B1(_2746_),
    .Y(_3529_));
 sky130_fd_sc_hd__nand2_1 _6601_ (.A(net111),
    .B(_2743_),
    .Y(_2747_));
 sky130_fd_sc_hd__o21ai_1 _6602_ (.A1(_3525_),
    .A2(_2743_),
    .B1(_2747_),
    .Y(_3271_));
 sky130_fd_sc_hd__nand2_1 _6603_ (.A(net122),
    .B(_2743_),
    .Y(_2748_));
 sky130_fd_sc_hd__o21ai_0 _6604_ (.A1(_3519_),
    .A2(_2743_),
    .B1(_2748_),
    .Y(_3534_));
 sky130_fd_sc_hd__nand2_1 _6605_ (.A(net125),
    .B(_2743_),
    .Y(_2749_));
 sky130_fd_sc_hd__o21ai_0 _6606_ (.A1(_1689_),
    .A2(_2743_),
    .B1(_2749_),
    .Y(_3538_));
 sky130_fd_sc_hd__nand2_1 _6607_ (.A(net126),
    .B(_2743_),
    .Y(_2750_));
 sky130_fd_sc_hd__o21ai_0 _6608_ (.A1(_3503_),
    .A2(_2743_),
    .B1(_2750_),
    .Y(_3544_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(net127),
    .B(_2743_),
    .Y(_2751_));
 sky130_fd_sc_hd__o21ai_0 _6610_ (.A1(_3495_),
    .A2(_2743_),
    .B1(_2751_),
    .Y(_3548_));
 sky130_fd_sc_hd__nand2_1 _6611_ (.A(net128),
    .B(_2743_),
    .Y(_2752_));
 sky130_fd_sc_hd__o21ai_0 _6612_ (.A1(net516),
    .A2(_2743_),
    .B1(_2752_),
    .Y(_3552_));
 sky130_fd_sc_hd__nand2_1 _6613_ (.A(net129),
    .B(_2743_),
    .Y(_2753_));
 sky130_fd_sc_hd__o21ai_0 _6614_ (.A1(_3479_),
    .A2(_2743_),
    .B1(_2753_),
    .Y(_3556_));
 sky130_fd_sc_hd__nand2_1 _6615_ (.A(net130),
    .B(_2743_),
    .Y(_2754_));
 sky130_fd_sc_hd__o21ai_0 _6616_ (.A1(_3471_),
    .A2(_2743_),
    .B1(_2754_),
    .Y(_3560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__nand2_1 _6618_ (.A(net131),
    .B(_2743_),
    .Y(_2756_));
 sky130_fd_sc_hd__o21ai_0 _6619_ (.A1(net854),
    .A2(_2743_),
    .B1(_2756_),
    .Y(_3564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__nand2_1 _6621_ (.A(net101),
    .B(_2743_),
    .Y(_2758_));
 sky130_fd_sc_hd__o21ai_0 _6622_ (.A1(_3455_),
    .A2(_2743_),
    .B1(_2758_),
    .Y(_3568_));
 sky130_fd_sc_hd__nand2_1 _6623_ (.A(net102),
    .B(_2743_),
    .Y(_2759_));
 sky130_fd_sc_hd__o21ai_0 _6624_ (.A1(_3447_),
    .A2(_2743_),
    .B1(_2759_),
    .Y(_3572_));
 sky130_fd_sc_hd__nand2_1 _6625_ (.A(net103),
    .B(_2743_),
    .Y(_2760_));
 sky130_fd_sc_hd__o21ai_0 _6626_ (.A1(_3439_),
    .A2(_2743_),
    .B1(_2760_),
    .Y(_3576_));
 sky130_fd_sc_hd__nand2_1 _6627_ (.A(net104),
    .B(_2743_),
    .Y(_2761_));
 sky130_fd_sc_hd__o21ai_0 _6628_ (.A1(_3431_),
    .A2(_2743_),
    .B1(_2761_),
    .Y(_3580_));
 sky130_fd_sc_hd__nand2_1 _6629_ (.A(net105),
    .B(_2743_),
    .Y(_2762_));
 sky130_fd_sc_hd__o21ai_0 _6630_ (.A1(_3423_),
    .A2(_2743_),
    .B1(_2762_),
    .Y(_3584_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(net106),
    .B(_2743_),
    .Y(_2763_));
 sky130_fd_sc_hd__o21ai_0 _6632_ (.A1(_3415_),
    .A2(_2743_),
    .B1(_2763_),
    .Y(_3588_));
 sky130_fd_sc_hd__nand2_1 _6633_ (.A(net107),
    .B(_2743_),
    .Y(_2764_));
 sky130_fd_sc_hd__o21ai_0 _6634_ (.A1(_3407_),
    .A2(_2743_),
    .B1(_2764_),
    .Y(_3592_));
 sky130_fd_sc_hd__nand2_1 _6635_ (.A(net108),
    .B(_2743_),
    .Y(_2765_));
 sky130_fd_sc_hd__o21ai_0 _6636_ (.A1(_3399_),
    .A2(_2743_),
    .B1(_2765_),
    .Y(_3596_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(net109),
    .B(_2743_),
    .Y(_2766_));
 sky130_fd_sc_hd__o21ai_0 _6638_ (.A1(_1031_),
    .A2(_2743_),
    .B1(_2766_),
    .Y(_3600_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__nand2_1 _6640_ (.A(net110),
    .B(_2743_),
    .Y(_2768_));
 sky130_fd_sc_hd__o21ai_0 _6641_ (.A1(_3383_),
    .A2(_2743_),
    .B1(_2768_),
    .Y(_3604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__nand2_1 _6643_ (.A(net112),
    .B(_2743_),
    .Y(_2770_));
 sky130_fd_sc_hd__o21ai_0 _6644_ (.A1(_3375_),
    .A2(_2743_),
    .B1(_2770_),
    .Y(_3608_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(net113),
    .B(_2743_),
    .Y(_2771_));
 sky130_fd_sc_hd__o21ai_0 _6646_ (.A1(_3367_),
    .A2(_2743_),
    .B1(_2771_),
    .Y(_3612_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(net114),
    .B(_2743_),
    .Y(_2772_));
 sky130_fd_sc_hd__o21ai_0 _6648_ (.A1(_3359_),
    .A2(_2743_),
    .B1(_2772_),
    .Y(_3616_));
 sky130_fd_sc_hd__nand2_1 _6649_ (.A(net115),
    .B(_2743_),
    .Y(_2773_));
 sky130_fd_sc_hd__o21ai_0 _6650_ (.A1(_3351_),
    .A2(_2743_),
    .B1(_2773_),
    .Y(_3620_));
 sky130_fd_sc_hd__nand2_1 _6651_ (.A(net116),
    .B(_2743_),
    .Y(_2774_));
 sky130_fd_sc_hd__o21ai_0 _6652_ (.A1(_3343_),
    .A2(_2743_),
    .B1(_2774_),
    .Y(_3624_));
 sky130_fd_sc_hd__nand2_1 _6653_ (.A(net117),
    .B(_2743_),
    .Y(_2775_));
 sky130_fd_sc_hd__o21ai_0 _6654_ (.A1(_3335_),
    .A2(_2743_),
    .B1(_2775_),
    .Y(_3628_));
 sky130_fd_sc_hd__nand2_1 _6655_ (.A(net118),
    .B(_2743_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21ai_0 _6656_ (.A1(_0621_),
    .A2(_2743_),
    .B1(_2776_),
    .Y(_3632_));
 sky130_fd_sc_hd__nand2_1 _6657_ (.A(net119),
    .B(_2743_),
    .Y(_2777_));
 sky130_fd_sc_hd__o21ai_0 _6658_ (.A1(_3319_),
    .A2(_2743_),
    .B1(_2777_),
    .Y(_3636_));
 sky130_fd_sc_hd__nand2_1 _6659_ (.A(net120),
    .B(_2743_),
    .Y(_2778_));
 sky130_fd_sc_hd__o21ai_0 _6660_ (.A1(_3311_),
    .A2(_2743_),
    .B1(_2778_),
    .Y(_3640_));
 sky130_fd_sc_hd__nand2_1 _6661_ (.A(net121),
    .B(_2743_),
    .Y(_2779_));
 sky130_fd_sc_hd__o21ai_0 _6662_ (.A1(_3303_),
    .A2(_2743_),
    .B1(_2779_),
    .Y(_3644_));
 sky130_fd_sc_hd__nand2_1 _6663_ (.A(net123),
    .B(_2743_),
    .Y(_2780_));
 sky130_fd_sc_hd__o21ai_0 _6664_ (.A1(_0371_),
    .A2(_2743_),
    .B1(_2780_),
    .Y(_3648_));
 sky130_fd_sc_hd__or3_4 _6665_ (.A(net27),
    .B(_0126_),
    .C(_0127_),
    .X(_2781_));
 sky130_fd_sc_hd__nor4_1 _6666_ (.A(net6),
    .B(net4),
    .C(net5),
    .D(_0120_),
    .Y(_2782_));
 sky130_fd_sc_hd__nor4b_1 _6667_ (.A(net6),
    .B(net5),
    .C(_0120_),
    .D_N(net4),
    .Y(_2783_));
 sky130_fd_sc_hd__nand2_1 _6668_ (.A(_0950_),
    .B(_3383_),
    .Y(_2784_));
 sky130_fd_sc_hd__nor2_1 _6669_ (.A(_0401_),
    .B(_0747_),
    .Y(_2785_));
 sky130_fd_sc_hd__nor2b_1 _6670_ (.A(_0794_),
    .B_N(_3359_),
    .Y(_2786_));
 sky130_fd_sc_hd__maj3_1 _6671_ (.A(_2785_),
    .B(_3351_),
    .C(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__inv_1 _6672_ (.A(_0838_),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2b_1 _6673_ (.A(_0881_),
    .B_N(_3375_),
    .Y(_2789_));
 sky130_fd_sc_hd__maj3_1 _6674_ (.A(_2788_),
    .B(_3367_),
    .C(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__nor2_1 _6675_ (.A(_2787_),
    .B(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__inv_1 _6676_ (.A(_1002_),
    .Y(_2792_));
 sky130_fd_sc_hd__nor3_1 _6677_ (.A(_1127_),
    .B(_1144_),
    .C(_1159_),
    .Y(_2793_));
 sky130_fd_sc_hd__maj3_1 _6678_ (.A(_1059_),
    .B(_3399_),
    .C(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__maj3_1 _6679_ (.A(_2792_),
    .B(_1031_),
    .C(_2794_),
    .X(_2795_));
 sky130_fd_sc_hd__o21ai_1 _6680_ (.A1(_0950_),
    .A2(_3383_),
    .B1(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__nand2b_1 _6681_ (.A_N(_3375_),
    .B(_0881_),
    .Y(_2797_));
 sky130_fd_sc_hd__maj3_1 _6682_ (.A(_2788_),
    .B(_3367_),
    .C(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2b_1 _6683_ (.A_N(_3359_),
    .B(_0794_),
    .Y(_2799_));
 sky130_fd_sc_hd__maj3_1 _6684_ (.A(_2785_),
    .B(_3351_),
    .C(_2799_),
    .X(_2800_));
 sky130_fd_sc_hd__o21ai_1 _6685_ (.A1(_2787_),
    .A2(_2798_),
    .B1(_2800_),
    .Y(_2801_));
 sky130_fd_sc_hd__a31oi_1 _6686_ (.A1(_2784_),
    .A2(_2791_),
    .A3(_2796_),
    .B1(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__a21oi_2 _6687_ (.A1(_0628_),
    .A2(_0634_),
    .B1(_0401_),
    .Y(_2803_));
 sky130_fd_sc_hd__nand2_1 _6688_ (.A(_2803_),
    .B(_3335_),
    .Y(_2804_));
 sky130_fd_sc_hd__nor2_1 _6689_ (.A(_2803_),
    .B(_3335_),
    .Y(_2805_));
 sky130_fd_sc_hd__a31oi_1 _6690_ (.A1(_0694_),
    .A2(_3339_),
    .A3(_2804_),
    .B1(_2805_),
    .Y(_2806_));
 sky130_fd_sc_hd__a21oi_1 _6691_ (.A1(_0516_),
    .A2(_3315_),
    .B1(_0571_),
    .Y(_2807_));
 sky130_fd_sc_hd__o21ai_0 _6692_ (.A1(_0621_),
    .A2(_2806_),
    .B1(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__nand2_1 _6693_ (.A(_0516_),
    .B(_3315_),
    .Y(_2809_));
 sky130_fd_sc_hd__nor2_1 _6694_ (.A(_0516_),
    .B(_3315_),
    .Y(_2810_));
 sky130_fd_sc_hd__a31oi_1 _6695_ (.A1(_0621_),
    .A2(_2809_),
    .A3(_2806_),
    .B1(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__nand2_2 _6696_ (.A(net5),
    .B(_1341_),
    .Y(_2812_));
 sky130_fd_sc_hd__nor2b_1 _6697_ (.A(_0274_),
    .B_N(_0298_),
    .Y(_2813_));
 sky130_fd_sc_hd__xnor2_1 _6698_ (.A(_0274_),
    .B(_0298_),
    .Y(_2814_));
 sky130_fd_sc_hd__inv_2 _6699_ (.A(_0324_),
    .Y(_2815_));
 sky130_fd_sc_hd__and2_0 _6700_ (.A(_2815_),
    .B(_0371_),
    .X(_2816_));
 sky130_fd_sc_hd__nor3b_1 _6701_ (.A(_0298_),
    .B(_2812_),
    .C_N(_0274_),
    .Y(_2817_));
 sky130_fd_sc_hd__a221oi_2 _6702_ (.A1(_2812_),
    .A2(_2813_),
    .B1(_2814_),
    .B2(_2816_),
    .C1(_2817_),
    .Y(_2818_));
 sky130_fd_sc_hd__o21ai_0 _6703_ (.A1(_0481_),
    .A2(_0495_),
    .B1(_0458_),
    .Y(_2819_));
 sky130_fd_sc_hd__maj3_1 _6704_ (.A(_0404_),
    .B(_3303_),
    .C(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__o211ai_1 _6705_ (.A1(_2815_),
    .A2(_0371_),
    .B1(_2814_),
    .C1(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__and2_2 _6706_ (.A(_2818_),
    .B(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__a21oi_1 _6707_ (.A1(_2808_),
    .A2(_2811_),
    .B1(_2822_),
    .Y(_2823_));
 sky130_fd_sc_hd__nor3_1 _6708_ (.A(_0694_),
    .B(_0720_),
    .C(_0735_),
    .Y(_2824_));
 sky130_fd_sc_hd__maj3_1 _6709_ (.A(_2803_),
    .B(_3335_),
    .C(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__a21o_1 _6710_ (.A1(_0621_),
    .A2(_2809_),
    .B1(_2807_),
    .X(_2826_));
 sky130_fd_sc_hd__a221oi_1 _6711_ (.A1(_0621_),
    .A2(_2807_),
    .B1(_2825_),
    .B2(_2826_),
    .C1(_2810_),
    .Y(_2827_));
 sky130_fd_sc_hd__nor2_1 _6712_ (.A(_2822_),
    .B(_2827_),
    .Y(_2828_));
 sky130_fd_sc_hd__nor3_1 _6713_ (.A(_0458_),
    .B(_0481_),
    .C(_0495_),
    .Y(_2829_));
 sky130_fd_sc_hd__maj3_1 _6714_ (.A(_0404_),
    .B(_3303_),
    .C(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__o211ai_1 _6715_ (.A1(_2815_),
    .A2(_0371_),
    .B1(_2814_),
    .C1(_2830_),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6716_ (.A(_2818_),
    .B(_2831_),
    .Y(_2832_));
 sky130_fd_sc_hd__a211o_2 _6717_ (.A1(_2802_),
    .A2(_2823_),
    .B1(_2828_),
    .C1(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__nand2_1 _6718_ (.A(_2808_),
    .B(_2811_),
    .Y(_2834_));
 sky130_fd_sc_hd__o21ai_0 _6719_ (.A1(_1144_),
    .A2(_1159_),
    .B1(_1127_),
    .Y(_2835_));
 sky130_fd_sc_hd__maj3_1 _6720_ (.A(_1059_),
    .B(_3399_),
    .C(_2835_),
    .X(_2836_));
 sky130_fd_sc_hd__a21oi_1 _6721_ (.A1(_1031_),
    .A2(_2836_),
    .B1(_2792_),
    .Y(_2837_));
 sky130_fd_sc_hd__nor3b_1 _6722_ (.A(_1031_),
    .B(_2836_),
    .C_N(_2784_),
    .Y(_2838_));
 sky130_fd_sc_hd__nor2_1 _6723_ (.A(_0950_),
    .B(_3383_),
    .Y(_2839_));
 sky130_fd_sc_hd__a211o_1 _6724_ (.A1(_2784_),
    .A2(_2837_),
    .B1(_2838_),
    .C1(_2839_),
    .X(_2840_));
 sky130_fd_sc_hd__a21oi_1 _6725_ (.A1(_2791_),
    .A2(_2840_),
    .B1(_2801_),
    .Y(_2841_));
 sky130_fd_sc_hd__nand3_1 _6726_ (.A(_2818_),
    .B(_2831_),
    .C(_2827_),
    .Y(_2842_));
 sky130_fd_sc_hd__nand2_1 _6727_ (.A(_1218_),
    .B(_3423_),
    .Y(_2843_));
 sky130_fd_sc_hd__maj3_1 _6728_ (.A(_1174_),
    .B(_3411_),
    .C(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__nand2_1 _6729_ (.A(_1299_),
    .B(_3435_),
    .Y(_2845_));
 sky130_fd_sc_hd__o21ai_0 _6730_ (.A1(_3431_),
    .A2(_2845_),
    .B1(_1264_),
    .Y(_2846_));
 sky130_fd_sc_hd__nand2_1 _6731_ (.A(_3431_),
    .B(_2845_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _6732_ (.A(_1218_),
    .B(_3423_),
    .Y(_2848_));
 sky130_fd_sc_hd__maj3_1 _6733_ (.A(_1174_),
    .B(_3411_),
    .C(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__a21o_1 _6734_ (.A1(_2846_),
    .A2(_2847_),
    .B1(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__a21oi_4 _6735_ (.A1(_2844_),
    .A2(_2850_),
    .B1(_2822_),
    .Y(_2851_));
 sky130_fd_sc_hd__o221ai_4 _6736_ (.A1(_2832_),
    .A2(_2834_),
    .B1(_2841_),
    .B2(_2842_),
    .C1(_2851_),
    .Y(_2852_));
 sky130_fd_sc_hd__nor2_1 _6737_ (.A(_1299_),
    .B(_3435_),
    .Y(_2853_));
 sky130_fd_sc_hd__nor2_1 _6738_ (.A(_3431_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__a21oi_1 _6739_ (.A1(_3431_),
    .A2(_2853_),
    .B1(_1264_),
    .Y(_2855_));
 sky130_fd_sc_hd__nor3_1 _6740_ (.A(_0401_),
    .B(_1340_),
    .C(_3443_),
    .Y(_2856_));
 sky130_fd_sc_hd__a21oi_4 _6741_ (.A1(_1411_),
    .A2(_1417_),
    .B1(_0401_),
    .Y(_2857_));
 sky130_fd_sc_hd__a221oi_1 _6742_ (.A1(_1462_),
    .A2(_1469_),
    .B1(_1474_),
    .B2(_1482_),
    .C1(_1455_),
    .Y(_2858_));
 sky130_fd_sc_hd__maj3_1 _6743_ (.A(_2857_),
    .B(net852),
    .C(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__maj3_1 _6744_ (.A(_1378_),
    .B(_3455_),
    .C(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__o21ai_1 _6745_ (.A1(_0401_),
    .A2(_1340_),
    .B1(_3443_),
    .Y(_2861_));
 sky130_fd_sc_hd__o21ai_1 _6746_ (.A1(_2856_),
    .A2(_2860_),
    .B1(_2861_),
    .Y(_2862_));
 sky130_fd_sc_hd__o311a_1 _6747_ (.A1(_2849_),
    .A2(_2854_),
    .A3(_2855_),
    .B1(_2862_),
    .C1(_2844_),
    .X(_2863_));
 sky130_fd_sc_hd__nand2b_1 _6748_ (.A_N(_3471_),
    .B(_1455_),
    .Y(_2864_));
 sky130_fd_sc_hd__maj3_1 _6749_ (.A(_2857_),
    .B(net852),
    .C(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__maj3_1 _6750_ (.A(_1378_),
    .B(_3455_),
    .C(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__o21ai_2 _6751_ (.A1(_2856_),
    .A2(_2866_),
    .B1(_2861_),
    .Y(_2867_));
 sky130_fd_sc_hd__nor2_1 _6752_ (.A(_1502_),
    .B(_3475_),
    .Y(_2868_));
 sky130_fd_sc_hd__nor2_1 _6753_ (.A(_1618_),
    .B(_3499_),
    .Y(_2869_));
 sky130_fd_sc_hd__maj3_1 _6754_ (.A(net160),
    .B(net521),
    .C(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__maj3_1 _6755_ (.A(net161),
    .B(net515),
    .C(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__nand2_1 _6756_ (.A(_1502_),
    .B(_3475_),
    .Y(_2872_));
 sky130_fd_sc_hd__o21a_1 _6757_ (.A1(_2868_),
    .A2(_2871_),
    .B1(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__nor2_1 _6758_ (.A(net412),
    .B(_3525_),
    .Y(_2874_));
 sky130_fd_sc_hd__nand2_1 _6759_ (.A(net412),
    .B(_3525_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor2b_1 _6760_ (.A(_2874_),
    .B_N(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__nand2_1 _6761_ (.A(_2872_),
    .B(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__nor2_1 _6762_ (.A(net158),
    .B(_1689_),
    .Y(_2878_));
 sky130_fd_sc_hd__nand2_1 _6763_ (.A(net158),
    .B(_1689_),
    .Y(_2879_));
 sky130_fd_sc_hd__a21oi_1 _6764_ (.A1(_1720_),
    .A2(_1731_),
    .B1(net155),
    .Y(_2880_));
 sky130_fd_sc_hd__nor2_1 _6765_ (.A(_1700_),
    .B(_3515_),
    .Y(_2881_));
 sky130_fd_sc_hd__xnor2_1 _6766_ (.A(net133),
    .B(net500),
    .Y(_2882_));
 sky130_fd_sc_hd__nor3_1 _6767_ (.A(_2880_),
    .B(_2881_),
    .C(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__or4bb_1 _6768_ (.A(_2877_),
    .B(_2878_),
    .C_N(_2879_),
    .D_N(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__nand2_1 _6769_ (.A(_1618_),
    .B(_3499_),
    .Y(_2885_));
 sky130_fd_sc_hd__maj3_1 _6770_ (.A(net160),
    .B(net522),
    .C(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__maj3_1 _6771_ (.A(net161),
    .B(net515),
    .C(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__nor2_1 _6772_ (.A(_2868_),
    .B(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__nor4_1 _6773_ (.A(_2867_),
    .B(_2873_),
    .C(_2884_),
    .D(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__nand4bb_1 _6774_ (.A_N(_2833_),
    .B_N(_2852_),
    .C(_2863_),
    .D(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__mux2i_2 _6775_ (.A0(_2782_),
    .A1(_2783_),
    .S(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__nor2_1 _6776_ (.A(_0120_),
    .B(_1801_),
    .Y(_2892_));
 sky130_fd_sc_hd__nor3_1 _6777_ (.A(_1813_),
    .B(net4),
    .C(_0120_),
    .Y(_2893_));
 sky130_fd_sc_hd__nand2_1 _6778_ (.A(net133),
    .B(net500),
    .Y(_2894_));
 sky130_fd_sc_hd__o211a_1 _6779_ (.A1(_2874_),
    .A2(_2894_),
    .B1(_2875_),
    .C1(_3515_),
    .X(_2895_));
 sky130_fd_sc_hd__o211a_1 _6780_ (.A1(_2874_),
    .A2(_2894_),
    .B1(_2875_),
    .C1(_1700_),
    .X(_2896_));
 sky130_fd_sc_hd__o41ai_1 _6781_ (.A1(_2878_),
    .A2(_2895_),
    .A3(_2880_),
    .A4(_2896_),
    .B1(_2879_),
    .Y(_2897_));
 sky130_fd_sc_hd__a31oi_1 _6782_ (.A1(_2872_),
    .A2(_2887_),
    .A3(_2897_),
    .B1(_2873_),
    .Y(_2898_));
 sky130_fd_sc_hd__o21a_1 _6783_ (.A1(_2867_),
    .A2(_2898_),
    .B1(_2863_),
    .X(_2899_));
 sky130_fd_sc_hd__o21bai_1 _6784_ (.A1(_2852_),
    .A2(_2899_),
    .B1_N(_2833_),
    .Y(_2900_));
 sky130_fd_sc_hd__mux2i_2 _6785_ (.A0(_2892_),
    .A1(_2893_),
    .S(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__nand3_4 _6786_ (.A(_2781_),
    .B(_2891_),
    .C(_2901_),
    .Y(_2902_));
 sky130_fd_sc_hd__mux2_1 _6787_ (.A0(net100),
    .A1(_3531_),
    .S(_2902_),
    .X(_0032_));
 sky130_fd_sc_hd__inv_1 _6788_ (.A(net111),
    .Y(_2903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__mux2i_1 _6790_ (.A0(_2903_),
    .A1(_3274_),
    .S(_2902_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _6791_ (.A(net129),
    .Y(_2905_));
 sky130_fd_sc_hd__nand3_1 _6792_ (.A(net126),
    .B(net127),
    .C(net128),
    .Y(_2906_));
 sky130_fd_sc_hd__nor2_1 _6793_ (.A(_2905_),
    .B(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__nand4_1 _6794_ (.A(_3542_),
    .B(net130),
    .C(net131),
    .D(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__xor2_2 _6795_ (.A(net101),
    .B(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__a21o_1 _6796_ (.A1(_3563_),
    .A2(_3558_),
    .B1(_3562_),
    .X(_2910_));
 sky130_fd_sc_hd__a21oi_4 _6797_ (.A1(_3567_),
    .A2(_2910_),
    .B1(_3566_),
    .Y(_2911_));
 sky130_fd_sc_hd__clkinvlp_4 _6798_ (.A(_3547_),
    .Y(_2912_));
 sky130_fd_sc_hd__a21o_1 _6799_ (.A1(_3273_),
    .A2(_3537_),
    .B1(_3536_),
    .X(_2913_));
 sky130_fd_sc_hd__a21oi_4 _6800_ (.A1(_2913_),
    .A2(_3541_),
    .B1(_3540_),
    .Y(_2914_));
 sky130_fd_sc_hd__nor3_2 _6801_ (.A(_3546_),
    .B(_3550_),
    .C(_3554_),
    .Y(_2915_));
 sky130_fd_sc_hd__o21ai_2 _6802_ (.A1(_2912_),
    .A2(_2914_),
    .B1(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__o21a_1 _6803_ (.A1(_3551_),
    .A2(_3550_),
    .B1(_3555_),
    .X(_2917_));
 sky130_fd_sc_hd__o21a_1 _6804_ (.A1(_3554_),
    .A2(_2917_),
    .B1(_3559_),
    .X(_2918_));
 sky130_fd_sc_hd__and3_1 _6805_ (.A(_3563_),
    .B(_3567_),
    .C(_2918_),
    .X(_2919_));
 sky130_fd_sc_hd__nand2_1 _6806_ (.A(_2916_),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__nand2_1 _6807_ (.A(_2911_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__xnor2_1 _6808_ (.A(_3571_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__mux2i_1 _6809_ (.A0(_2909_),
    .A1(_2922_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[10] ));
 sky130_fd_sc_hd__nand2_1 _6810_ (.A(net122),
    .B(net125),
    .Y(_2923_));
 sky130_fd_sc_hd__nor3_2 _6811_ (.A(_2905_),
    .B(_2906_),
    .C(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__nand4_1 _6812_ (.A(net130),
    .B(net131),
    .C(net101),
    .D(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__xor2_1 _6813_ (.A(net102),
    .B(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__a21o_1 _6814_ (.A1(_3270_),
    .A2(_3533_),
    .B1(_3532_),
    .X(_2927_));
 sky130_fd_sc_hd__a21o_1 _6815_ (.A1(_3537_),
    .A2(_2927_),
    .B1(_3536_),
    .X(_2928_));
 sky130_fd_sc_hd__a21oi_2 _6816_ (.A1(_3541_),
    .A2(_2928_),
    .B1(_3540_),
    .Y(_2929_));
 sky130_fd_sc_hd__nor2_1 _6817_ (.A(_2912_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__nor2b_1 _6818_ (.A(_2930_),
    .B_N(_2915_),
    .Y(_2931_));
 sky130_fd_sc_hd__inv_1 _6819_ (.A(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__nand2_1 _6820_ (.A(_2919_),
    .B(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _6821_ (.A(_2911_),
    .B(_2933_),
    .Y(_2934_));
 sky130_fd_sc_hd__a21oi_1 _6822_ (.A1(_3571_),
    .A2(_2934_),
    .B1(_3570_),
    .Y(_2935_));
 sky130_fd_sc_hd__xor2_1 _6823_ (.A(_3575_),
    .B(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__mux2i_1 _6824_ (.A0(_2926_),
    .A1(_2936_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[11] ));
 sky130_fd_sc_hd__nand2_2 _6825_ (.A(_3542_),
    .B(_2907_),
    .Y(_2937_));
 sky130_fd_sc_hd__nand4_1 _6826_ (.A(net130),
    .B(net131),
    .C(net101),
    .D(net102),
    .Y(_2938_));
 sky130_fd_sc_hd__nor2_1 _6827_ (.A(_2937_),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__xnor2_4 _6828_ (.A(net103),
    .B(_2939_),
    .Y(_2940_));
 sky130_fd_sc_hd__inv_1 _6829_ (.A(_3574_),
    .Y(_2941_));
 sky130_fd_sc_hd__o21ai_1 _6830_ (.A1(_3571_),
    .A2(_3570_),
    .B1(_3575_),
    .Y(_2942_));
 sky130_fd_sc_hd__nor2_1 _6831_ (.A(_3570_),
    .B(_3574_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_1 _6832_ (.A(_2911_),
    .B(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21oi_4 _6833_ (.A1(_2919_),
    .A2(_2916_),
    .B1(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__a21oi_1 _6834_ (.A1(_2941_),
    .A2(_2942_),
    .B1(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__xnor2_2 _6835_ (.A(_3579_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__mux2i_1 _6836_ (.A0(_2940_),
    .A1(_2947_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[12] ));
 sky130_fd_sc_hd__inv_1 _6837_ (.A(net103),
    .Y(_2948_));
 sky130_fd_sc_hd__nor2_1 _6838_ (.A(_2948_),
    .B(_2938_),
    .Y(_2949_));
 sky130_fd_sc_hd__nand2_1 _6839_ (.A(_2924_),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__xor2_1 _6840_ (.A(net104),
    .B(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__a21boi_2 _6841_ (.A1(_2941_),
    .A2(_2942_),
    .B1_N(_3579_),
    .Y(_2952_));
 sky130_fd_sc_hd__or2_1 _6842_ (.A(_2919_),
    .B(_2944_),
    .X(_2953_));
 sky130_fd_sc_hd__o2111ai_4 _6843_ (.A1(_2912_),
    .A2(_2929_),
    .B1(_2943_),
    .C1(_2911_),
    .D1(_2915_),
    .Y(_2954_));
 sky130_fd_sc_hd__a31oi_2 _6844_ (.A1(_2952_),
    .A2(_2953_),
    .A3(_2954_),
    .B1(_3578_),
    .Y(_2955_));
 sky130_fd_sc_hd__xor2_2 _6845_ (.A(_3583_),
    .B(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__mux2i_1 _6846_ (.A0(_2951_),
    .A1(_2956_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[13] ));
 sky130_fd_sc_hd__nand4_1 _6847_ (.A(_3542_),
    .B(net104),
    .C(_2907_),
    .D(_2949_),
    .Y(_2957_));
 sky130_fd_sc_hd__xor2_1 _6848_ (.A(net105),
    .B(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__inv_1 _6849_ (.A(_2952_),
    .Y(_2959_));
 sky130_fd_sc_hd__o21bai_1 _6850_ (.A1(_2945_),
    .A2(_2959_),
    .B1_N(_3578_),
    .Y(_2960_));
 sky130_fd_sc_hd__a21oi_2 _6851_ (.A1(_3583_),
    .A2(_2960_),
    .B1(_3582_),
    .Y(_2961_));
 sky130_fd_sc_hd__xor2_4 _6852_ (.A(_3587_),
    .B(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__mux2i_1 _6853_ (.A0(_2958_),
    .A1(_2962_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[14] ));
 sky130_fd_sc_hd__nand4_1 _6854_ (.A(net104),
    .B(net105),
    .C(_2924_),
    .D(_2949_),
    .Y(_2963_));
 sky130_fd_sc_hd__xor2_1 _6855_ (.A(net106),
    .B(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__o211a_1 _6856_ (.A1(_3587_),
    .A2(_3586_),
    .B1(_2952_),
    .C1(_3583_),
    .X(_2965_));
 sky130_fd_sc_hd__a21o_1 _6857_ (.A1(_3583_),
    .A2(_3578_),
    .B1(_3582_),
    .X(_2966_));
 sky130_fd_sc_hd__a21o_1 _6858_ (.A1(_3587_),
    .A2(_2966_),
    .B1(_3586_),
    .X(_2967_));
 sky130_fd_sc_hd__a31oi_4 _6859_ (.A1(_2953_),
    .A2(_2954_),
    .A3(_2965_),
    .B1(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__xor2_1 _6860_ (.A(_3591_),
    .B(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__mux2i_1 _6861_ (.A0(_2964_),
    .A1(_2969_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[15] ));
 sky130_fd_sc_hd__and4_1 _6862_ (.A(net104),
    .B(net105),
    .C(net106),
    .D(_2949_),
    .X(_2970_));
 sky130_fd_sc_hd__nor2b_4 _6863_ (.A(_2937_),
    .B_N(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__xnor2_1 _6864_ (.A(net107),
    .B(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__nand4_1 _6865_ (.A(_3583_),
    .B(_3587_),
    .C(_3591_),
    .D(_2952_),
    .Y(_2973_));
 sky130_fd_sc_hd__a21oi_1 _6866_ (.A1(_3591_),
    .A2(_2967_),
    .B1(_3590_),
    .Y(_2974_));
 sky130_fd_sc_hd__o21ai_4 _6867_ (.A1(_2945_),
    .A2(_2973_),
    .B1(_2974_),
    .Y(_2975_));
 sky130_fd_sc_hd__xnor2_2 _6868_ (.A(_3595_),
    .B(_2975_),
    .Y(_2976_));
 sky130_fd_sc_hd__mux2i_1 _6869_ (.A0(_2972_),
    .A1(_2976_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[16] ));
 sky130_fd_sc_hd__and3_4 _6870_ (.A(net107),
    .B(_2924_),
    .C(_2970_),
    .X(_2977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__xnor2_1 _6872_ (.A(net108),
    .B(_2977_),
    .Y(_2979_));
 sky130_fd_sc_hd__nand2_1 _6873_ (.A(_3591_),
    .B(_3595_),
    .Y(_2980_));
 sky130_fd_sc_hd__a21oi_1 _6874_ (.A1(_3595_),
    .A2(_3590_),
    .B1(_3594_),
    .Y(_2981_));
 sky130_fd_sc_hd__o21ai_4 _6875_ (.A1(_2968_),
    .A2(_2980_),
    .B1(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__xnor2_4 _6876_ (.A(_3599_),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__mux2i_1 _6877_ (.A0(_2979_),
    .A1(_2983_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[17] ));
 sky130_fd_sc_hd__nand3_1 _6878_ (.A(net107),
    .B(net108),
    .C(_2971_),
    .Y(_2984_));
 sky130_fd_sc_hd__xor2_1 _6879_ (.A(net109),
    .B(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__a21o_1 _6880_ (.A1(_3595_),
    .A2(_2975_),
    .B1(_3594_),
    .X(_2986_));
 sky130_fd_sc_hd__a21oi_2 _6881_ (.A1(_3599_),
    .A2(_2986_),
    .B1(_3598_),
    .Y(_2987_));
 sky130_fd_sc_hd__xor2_4 _6882_ (.A(_3603_),
    .B(_2987_),
    .X(_2988_));
 sky130_fd_sc_hd__mux2i_1 _6883_ (.A0(_2985_),
    .A1(_2988_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[18] ));
 sky130_fd_sc_hd__nand3_1 _6884_ (.A(net108),
    .B(net109),
    .C(_2977_),
    .Y(_2989_));
 sky130_fd_sc_hd__xor2_1 _6885_ (.A(net110),
    .B(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__inv_1 _6886_ (.A(_3602_),
    .Y(_2991_));
 sky130_fd_sc_hd__o21ai_1 _6887_ (.A1(_3599_),
    .A2(_3598_),
    .B1(_3603_),
    .Y(_2992_));
 sky130_fd_sc_hd__nand2_1 _6888_ (.A(_2991_),
    .B(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__o31a_2 _6889_ (.A1(_3598_),
    .A2(_3602_),
    .A3(_2982_),
    .B1(_2993_),
    .X(_2994_));
 sky130_fd_sc_hd__xnor2_4 _6890_ (.A(_3607_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__mux2i_1 _6892_ (.A0(_2990_),
    .A1(_2995_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[19] ));
 sky130_fd_sc_hd__nand2_1 _6893_ (.A(net107),
    .B(_2971_),
    .Y(_2997_));
 sky130_fd_sc_hd__nand3_1 _6894_ (.A(net108),
    .B(net109),
    .C(net110),
    .Y(_2998_));
 sky130_fd_sc_hd__nor2_1 _6895_ (.A(_2997_),
    .B(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__xnor2_2 _6896_ (.A(net112),
    .B(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hd__a211oi_4 _6897_ (.A1(_2975_),
    .A2(_3595_),
    .B1(_3598_),
    .C1(_3594_),
    .Y(_3001_));
 sky130_fd_sc_hd__o21ai_0 _6898_ (.A1(_3001_),
    .A2(_2992_),
    .B1(_2991_),
    .Y(_3002_));
 sky130_fd_sc_hd__a21oi_1 _6899_ (.A1(_3607_),
    .A2(_3002_),
    .B1(_3606_),
    .Y(_3003_));
 sky130_fd_sc_hd__xor2_2 _6900_ (.A(_3611_),
    .B(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__mux2i_1 _6901_ (.A0(_3000_),
    .A1(_3004_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[20] ));
 sky130_fd_sc_hd__inv_1 _6902_ (.A(net112),
    .Y(_3005_));
 sky130_fd_sc_hd__nor2_1 _6903_ (.A(_3005_),
    .B(_2998_),
    .Y(_3006_));
 sky130_fd_sc_hd__nand2_1 _6904_ (.A(_2977_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__xor2_1 _6905_ (.A(net113),
    .B(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__a21o_1 _6906_ (.A1(_3607_),
    .A2(_2994_),
    .B1(_3606_),
    .X(_3009_));
 sky130_fd_sc_hd__a21oi_1 _6907_ (.A1(_3611_),
    .A2(_3009_),
    .B1(_3610_),
    .Y(_3010_));
 sky130_fd_sc_hd__xor2_2 _6908_ (.A(_3615_),
    .B(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__mux2i_1 _6909_ (.A0(_3008_),
    .A1(_3011_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[21] ));
 sky130_fd_sc_hd__nand4_1 _6910_ (.A(net107),
    .B(net113),
    .C(_2971_),
    .D(_3006_),
    .Y(_3012_));
 sky130_fd_sc_hd__xor2_1 _6911_ (.A(net114),
    .B(_3012_),
    .X(_3013_));
 sky130_fd_sc_hd__nor3_1 _6912_ (.A(_3602_),
    .B(_3606_),
    .C(_3610_),
    .Y(_3014_));
 sky130_fd_sc_hd__o21ai_2 _6913_ (.A1(_3001_),
    .A2(_2992_),
    .B1(_3014_),
    .Y(_3015_));
 sky130_fd_sc_hd__nor3_1 _6914_ (.A(_3607_),
    .B(_3606_),
    .C(_3610_),
    .Y(_3016_));
 sky130_fd_sc_hd__nor2_1 _6915_ (.A(_3611_),
    .B(_3610_),
    .Y(_3017_));
 sky130_fd_sc_hd__nor2_1 _6916_ (.A(_3016_),
    .B(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__a31oi_2 _6917_ (.A1(_3615_),
    .A2(_3015_),
    .A3(_3018_),
    .B1(_3614_),
    .Y(_3019_));
 sky130_fd_sc_hd__xor2_2 _6918_ (.A(_3619_),
    .B(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__mux2i_1 _6919_ (.A0(_3013_),
    .A1(_3020_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[22] ));
 sky130_fd_sc_hd__and3_1 _6920_ (.A(net113),
    .B(net114),
    .C(_3006_),
    .X(_3021_));
 sky130_fd_sc_hd__nand2_1 _6921_ (.A(_2977_),
    .B(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__xor2_1 _6922_ (.A(net115),
    .B(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__and3_1 _6923_ (.A(_3607_),
    .B(_3611_),
    .C(_3615_),
    .X(_3024_));
 sky130_fd_sc_hd__o311ai_4 _6924_ (.A1(_3598_),
    .A2(_3602_),
    .A3(_2982_),
    .B1(_2993_),
    .C1(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__and3_1 _6925_ (.A(_3611_),
    .B(_3615_),
    .C(_3606_),
    .X(_3026_));
 sky130_fd_sc_hd__a21oi_1 _6926_ (.A1(_3615_),
    .A2(_3610_),
    .B1(_3026_),
    .Y(_3027_));
 sky130_fd_sc_hd__nand2_1 _6927_ (.A(_3025_),
    .B(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__o21ai_0 _6928_ (.A1(_3614_),
    .A2(_3028_),
    .B1(_3619_),
    .Y(_3029_));
 sky130_fd_sc_hd__nand2b_1 _6929_ (.A_N(_3618_),
    .B(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__xnor2_1 _6930_ (.A(_3623_),
    .B(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__mux2i_1 _6931_ (.A0(_3023_),
    .A1(_3031_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[23] ));
 sky130_fd_sc_hd__nand4_1 _6932_ (.A(net107),
    .B(net115),
    .C(_2971_),
    .D(_3021_),
    .Y(_3032_));
 sky130_fd_sc_hd__xor2_1 _6933_ (.A(net116),
    .B(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__and3_1 _6934_ (.A(_3615_),
    .B(_3619_),
    .C(_3623_),
    .X(_3034_));
 sky130_fd_sc_hd__nand3_1 _6935_ (.A(_3015_),
    .B(_3018_),
    .C(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__and3_1 _6936_ (.A(_3619_),
    .B(_3623_),
    .C(_3614_),
    .X(_3036_));
 sky130_fd_sc_hd__a21oi_1 _6937_ (.A1(_3623_),
    .A2(_3618_),
    .B1(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__and2_1 _6938_ (.A(_3035_),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__nand2b_1 _6939_ (.A_N(_3622_),
    .B(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__xor2_1 _6940_ (.A(_3627_),
    .B(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__inv_1 _6941_ (.A(_3040_),
    .Y(_3041_));
 sky130_fd_sc_hd__mux2i_1 _6942_ (.A0(_3033_),
    .A1(_3041_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[24] ));
 sky130_fd_sc_hd__and3_1 _6943_ (.A(net115),
    .B(net116),
    .C(_3021_),
    .X(_3042_));
 sky130_fd_sc_hd__nand2_1 _6944_ (.A(_2977_),
    .B(_3042_),
    .Y(_3043_));
 sky130_fd_sc_hd__xor2_1 _6945_ (.A(net117),
    .B(_3043_),
    .X(_3044_));
 sky130_fd_sc_hd__nor3_1 _6946_ (.A(_3614_),
    .B(_3618_),
    .C(_3622_),
    .Y(_3045_));
 sky130_fd_sc_hd__or2_0 _6947_ (.A(_3619_),
    .B(_3618_),
    .X(_3046_));
 sky130_fd_sc_hd__a21oi_1 _6948_ (.A1(_3623_),
    .A2(_3046_),
    .B1(_3622_),
    .Y(_3047_));
 sky130_fd_sc_hd__a31oi_2 _6949_ (.A1(_3025_),
    .A2(_3027_),
    .A3(_3045_),
    .B1(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21oi_1 _6950_ (.A1(_3627_),
    .A2(_3048_),
    .B1(_3626_),
    .Y(_3049_));
 sky130_fd_sc_hd__xor2_1 _6951_ (.A(_3631_),
    .B(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__mux2i_1 _6952_ (.A0(_3044_),
    .A1(_3050_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[25] ));
 sky130_fd_sc_hd__nand2_1 _6953_ (.A(net117),
    .B(_3042_),
    .Y(_3051_));
 sky130_fd_sc_hd__nor2_1 _6954_ (.A(_2997_),
    .B(_3051_),
    .Y(_3052_));
 sky130_fd_sc_hd__xnor2_1 _6955_ (.A(net118),
    .B(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__nor3_1 _6956_ (.A(_3622_),
    .B(_3626_),
    .C(_3630_),
    .Y(_3054_));
 sky130_fd_sc_hd__or2_0 _6957_ (.A(_3627_),
    .B(_3626_),
    .X(_3055_));
 sky130_fd_sc_hd__a21oi_1 _6958_ (.A1(_3631_),
    .A2(_3055_),
    .B1(_3630_),
    .Y(_3056_));
 sky130_fd_sc_hd__a21oi_1 _6959_ (.A1(_3038_),
    .A2(_3054_),
    .B1(_3056_),
    .Y(_3057_));
 sky130_fd_sc_hd__xnor2_2 _6960_ (.A(_3635_),
    .B(_3057_),
    .Y(_3058_));
 sky130_fd_sc_hd__mux2i_1 _6961_ (.A0(_3053_),
    .A1(_3058_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[26] ));
 sky130_fd_sc_hd__and4_1 _6962_ (.A(net117),
    .B(net118),
    .C(_2977_),
    .D(_3042_),
    .X(_3059_));
 sky130_fd_sc_hd__xnor2_1 _6963_ (.A(net119),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__nand2_1 _6964_ (.A(_3635_),
    .B(_3630_),
    .Y(_3061_));
 sky130_fd_sc_hd__nand3_1 _6965_ (.A(_3631_),
    .B(_3635_),
    .C(_3626_),
    .Y(_3062_));
 sky130_fd_sc_hd__nand2_1 _6966_ (.A(_3061_),
    .B(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__a41oi_2 _6967_ (.A1(_3627_),
    .A2(_3631_),
    .A3(_3635_),
    .A4(_3048_),
    .B1(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__nor2b_1 _6968_ (.A(_3634_),
    .B_N(_3064_),
    .Y(_3065_));
 sky130_fd_sc_hd__xor2_1 _6969_ (.A(_3639_),
    .B(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__mux2i_1 _6970_ (.A0(_3060_),
    .A1(_3066_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[27] ));
 sky130_fd_sc_hd__nand3_1 _6971_ (.A(net118),
    .B(net119),
    .C(_3052_),
    .Y(_3067_));
 sky130_fd_sc_hd__xor2_2 _6972_ (.A(net120),
    .B(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__inv_1 _6973_ (.A(_3635_),
    .Y(_3069_));
 sky130_fd_sc_hd__a311oi_1 _6974_ (.A1(_3035_),
    .A2(_3037_),
    .A3(_3054_),
    .B1(_3056_),
    .C1(_3069_),
    .Y(_3070_));
 sky130_fd_sc_hd__o21ai_1 _6975_ (.A1(_3634_),
    .A2(_3070_),
    .B1(_3639_),
    .Y(_3071_));
 sky130_fd_sc_hd__nor2_1 _6976_ (.A(_3643_),
    .B(_3638_),
    .Y(_3072_));
 sky130_fd_sc_hd__inv_1 _6977_ (.A(_3638_),
    .Y(_3073_));
 sky130_fd_sc_hd__a21boi_1 _6978_ (.A1(_3073_),
    .A2(_3071_),
    .B1_N(_3643_),
    .Y(_3074_));
 sky130_fd_sc_hd__a21o_1 _6979_ (.A1(_3071_),
    .A2(_3072_),
    .B1(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__mux2i_1 _6980_ (.A0(_3068_),
    .A1(_3075_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[28] ));
 sky130_fd_sc_hd__nand3_1 _6981_ (.A(net119),
    .B(net120),
    .C(_3059_),
    .Y(_3076_));
 sky130_fd_sc_hd__xor2_1 _6982_ (.A(net121),
    .B(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__nor3_1 _6983_ (.A(_3634_),
    .B(_3638_),
    .C(_3642_),
    .Y(_3078_));
 sky130_fd_sc_hd__or2_0 _6984_ (.A(_3639_),
    .B(_3638_),
    .X(_3079_));
 sky130_fd_sc_hd__a21oi_1 _6985_ (.A1(_3643_),
    .A2(_3079_),
    .B1(_3642_),
    .Y(_3080_));
 sky130_fd_sc_hd__a21oi_1 _6986_ (.A1(_3064_),
    .A2(_3078_),
    .B1(_3080_),
    .Y(_3081_));
 sky130_fd_sc_hd__xnor2_1 _6987_ (.A(_3647_),
    .B(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__mux2i_1 _6989_ (.A0(_3077_),
    .A1(_3082_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[29] ));
 sky130_fd_sc_hd__xnor2_1 _6990_ (.A(_3273_),
    .B(_3537_),
    .Y(_3084_));
 sky130_fd_sc_hd__mux2i_1 _6991_ (.A0(net122),
    .A1(_3084_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[2] ));
 sky130_fd_sc_hd__and3_1 _6992_ (.A(net119),
    .B(net120),
    .C(net121),
    .X(_3085_));
 sky130_fd_sc_hd__nand3_1 _6993_ (.A(net118),
    .B(_3052_),
    .C(_3085_),
    .Y(_3086_));
 sky130_fd_sc_hd__xor2_2 _6994_ (.A(net123),
    .B(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__nor3b_1 _6995_ (.A(_3642_),
    .B(_3646_),
    .C_N(_3651_),
    .Y(_3088_));
 sky130_fd_sc_hd__nor2b_1 _6996_ (.A(_3651_),
    .B_N(_3647_),
    .Y(_3089_));
 sky130_fd_sc_hd__mux2_1 _6997_ (.A0(_3088_),
    .A1(_3089_),
    .S(_3074_),
    .X(_3090_));
 sky130_fd_sc_hd__inv_1 _6998_ (.A(_3646_),
    .Y(_3091_));
 sky130_fd_sc_hd__nor3b_1 _6999_ (.A(_3647_),
    .B(_3646_),
    .C_N(_3651_),
    .Y(_3092_));
 sky130_fd_sc_hd__a21oi_1 _7000_ (.A1(_3642_),
    .A2(_3089_),
    .B1(_3092_),
    .Y(_3093_));
 sky130_fd_sc_hd__o21ai_0 _7001_ (.A1(_3651_),
    .A2(_3091_),
    .B1(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__nor2_1 _7002_ (.A(_3090_),
    .B(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__mux2i_1 _7003_ (.A0(_3087_),
    .A1(_3095_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[30] ));
 sky130_fd_sc_hd__nand3_1 _7004_ (.A(net123),
    .B(_3059_),
    .C(_3085_),
    .Y(_3096_));
 sky130_fd_sc_hd__xor2_2 _7005_ (.A(net124),
    .B(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__nand2_1 _7006_ (.A(net124),
    .B(_2743_),
    .Y(_3098_));
 sky130_fd_sc_hd__o21ai_0 _7007_ (.A1(_0274_),
    .A2(_2743_),
    .B1(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__xnor2_1 _7008_ (.A(net25),
    .B(_3099_),
    .Y(_3100_));
 sky130_fd_sc_hd__a21o_1 _7009_ (.A1(_3647_),
    .A2(_3081_),
    .B1(_3646_),
    .X(_3101_));
 sky130_fd_sc_hd__a21oi_2 _7010_ (.A1(_3651_),
    .A2(_3101_),
    .B1(_3650_),
    .Y(_3102_));
 sky130_fd_sc_hd__xnor2_2 _7011_ (.A(_3102_),
    .B(_3100_),
    .Y(_3103_));
 sky130_fd_sc_hd__mux2i_1 _7012_ (.A0(_3097_),
    .A1(_3103_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[31] ));
 sky130_fd_sc_hd__xor2_1 _7013_ (.A(_3541_),
    .B(_2928_),
    .X(_3104_));
 sky130_fd_sc_hd__mux2_1 _7014_ (.A0(_3543_),
    .A1(_3104_),
    .S(_2902_),
    .X(\dp.ISRmux.d0[3] ));
 sky130_fd_sc_hd__xnor2_1 _7015_ (.A(net126),
    .B(_3542_),
    .Y(_3105_));
 sky130_fd_sc_hd__xnor2_1 _7016_ (.A(_2912_),
    .B(_2914_),
    .Y(_3106_));
 sky130_fd_sc_hd__mux2i_1 _7017_ (.A0(_3105_),
    .A1(_3106_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[4] ));
 sky130_fd_sc_hd__nand3_1 _7018_ (.A(net122),
    .B(net125),
    .C(net126),
    .Y(_3107_));
 sky130_fd_sc_hd__xor2_1 _7019_ (.A(net127),
    .B(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__nor2_1 _7020_ (.A(_3546_),
    .B(_2930_),
    .Y(_3109_));
 sky130_fd_sc_hd__xor2_1 _7021_ (.A(_3551_),
    .B(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__mux2i_1 _7022_ (.A0(_3108_),
    .A1(_3110_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[5] ));
 sky130_fd_sc_hd__nand3_1 _7023_ (.A(net126),
    .B(_3542_),
    .C(net127),
    .Y(_3111_));
 sky130_fd_sc_hd__xor2_1 _7024_ (.A(net128),
    .B(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__o21bai_1 _7025_ (.A1(_2912_),
    .A2(_2914_),
    .B1_N(_3546_),
    .Y(_3113_));
 sky130_fd_sc_hd__a21oi_1 _7026_ (.A1(_3551_),
    .A2(_3113_),
    .B1(_3550_),
    .Y(_3114_));
 sky130_fd_sc_hd__xor2_1 _7027_ (.A(_3555_),
    .B(_3114_),
    .X(_3115_));
 sky130_fd_sc_hd__mux2i_1 _7028_ (.A0(_3112_),
    .A1(_3115_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[6] ));
 sky130_fd_sc_hd__nor2_1 _7029_ (.A(_2906_),
    .B(_2923_),
    .Y(_3116_));
 sky130_fd_sc_hd__xnor2_2 _7030_ (.A(net129),
    .B(_3116_),
    .Y(_3117_));
 sky130_fd_sc_hd__nor2_1 _7031_ (.A(_3554_),
    .B(_2917_),
    .Y(_3118_));
 sky130_fd_sc_hd__nor2_1 _7032_ (.A(_3118_),
    .B(_2931_),
    .Y(_3119_));
 sky130_fd_sc_hd__xnor2_2 _7033_ (.A(_3559_),
    .B(_3119_),
    .Y(_3120_));
 sky130_fd_sc_hd__mux2i_1 _7034_ (.A0(_3117_),
    .A1(_3120_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[7] ));
 sky130_fd_sc_hd__xor2_1 _7035_ (.A(net130),
    .B(_2937_),
    .X(_3121_));
 sky130_fd_sc_hd__a21oi_1 _7036_ (.A1(_2916_),
    .A2(_2918_),
    .B1(_3558_),
    .Y(_3122_));
 sky130_fd_sc_hd__xor2_2 _7037_ (.A(_3563_),
    .B(_3122_),
    .X(_3123_));
 sky130_fd_sc_hd__mux2i_1 _7038_ (.A0(_3121_),
    .A1(_3123_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[8] ));
 sky130_fd_sc_hd__nand2_1 _7039_ (.A(net130),
    .B(_2924_),
    .Y(_3124_));
 sky130_fd_sc_hd__xor2_1 _7040_ (.A(net131),
    .B(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__a21o_1 _7041_ (.A1(_2918_),
    .A2(_2932_),
    .B1(_3558_),
    .X(_3126_));
 sky130_fd_sc_hd__a21oi_1 _7042_ (.A1(_3563_),
    .A2(_3126_),
    .B1(_3562_),
    .Y(_3127_));
 sky130_fd_sc_hd__xor2_2 _7043_ (.A(_3567_),
    .B(_3127_),
    .X(_3128_));
 sky130_fd_sc_hd__mux2i_1 _7044_ (.A0(_3125_),
    .A1(_3128_),
    .S(_2902_),
    .Y(\dp.ISRmux.d0[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__nand2_1 _7046_ (.A(net66),
    .B(_1960_),
    .Y(_3130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__nand2_8 _7048_ (.A(_2781_),
    .B(_2741_),
    .Y(_3132_));
 sky130_fd_sc_hd__a21oi_1 _7049_ (.A1(net33),
    .A2(net98),
    .B1(_3132_),
    .Y(_3133_));
 sky130_fd_sc_hd__o22ai_2 _7050_ (.A1(net100),
    .A2(_2781_),
    .B1(_2741_),
    .B2(_3531_),
    .Y(_3134_));
 sky130_fd_sc_hd__a21oi_4 _7051_ (.A1(_3130_),
    .A2(_3133_),
    .B1(_3134_),
    .Y(\dp.result2[0] ));
 sky130_fd_sc_hd__nor2_8 _7052_ (.A(net28),
    .B(_0119_),
    .Y(_3135_));
 sky130_fd_sc_hd__nor2_8 _7053_ (.A(_0128_),
    .B(_3135_),
    .Y(_3136_));
 sky130_fd_sc_hd__nand2_8 _7054_ (.A(_1960_),
    .B(_3136_),
    .Y(_3137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__nand3b_4 _7056_ (.A_N(net99),
    .B(_0109_),
    .C(_1805_),
    .Y(_3139_));
 sky130_fd_sc_hd__nor4_4 _7057_ (.A(net4),
    .B(net5),
    .C(net99),
    .D(_1797_),
    .Y(_3140_));
 sky130_fd_sc_hd__a31o_4 _7058_ (.A1(_1813_),
    .A2(net62),
    .A3(net273),
    .B1(_1960_),
    .X(_3141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__a21oi_2 _7060_ (.A1(net34),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3143_));
 sky130_fd_sc_hd__a221oi_4 _7061_ (.A1(net202),
    .A2(_2909_),
    .B1(_2922_),
    .B2(_3135_),
    .C1(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__o21a_4 _7062_ (.A1(net67),
    .A2(_3137_),
    .B1(_3144_),
    .X(\dp.result2[10] ));
 sky130_fd_sc_hd__a21oi_1 _7063_ (.A1(net35),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3145_));
 sky130_fd_sc_hd__a221oi_1 _7064_ (.A1(net202),
    .A2(_2926_),
    .B1(_2936_),
    .B2(_3135_),
    .C1(_3145_),
    .Y(_3146_));
 sky130_fd_sc_hd__o21a_4 _7065_ (.A1(net68),
    .A2(_3137_),
    .B1(_3146_),
    .X(\dp.result2[11] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__a21oi_1 _7068_ (.A1(net36),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3149_));
 sky130_fd_sc_hd__nor2_1 _7069_ (.A(_3132_),
    .B(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__o21ai_4 _7070_ (.A1(net98),
    .A2(net69),
    .B1(_3150_),
    .Y(_3151_));
 sky130_fd_sc_hd__o221ai_4 _7071_ (.A1(_2781_),
    .A2(_2940_),
    .B1(_2947_),
    .B2(_2741_),
    .C1(_3151_),
    .Y(\dp.result2[12] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__nand2_1 _7073_ (.A(_3135_),
    .B(_2956_),
    .Y(_3153_));
 sky130_fd_sc_hd__a21oi_1 _7074_ (.A1(net37),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3154_));
 sky130_fd_sc_hd__a21oi_1 _7075_ (.A1(net202),
    .A2(_2951_),
    .B1(_3154_),
    .Y(_3155_));
 sky130_fd_sc_hd__o211a_4 _7076_ (.A1(net70),
    .A2(_3137_),
    .B1(_3153_),
    .C1(_3155_),
    .X(\dp.result2[13] ));
 sky130_fd_sc_hd__a21oi_1 _7077_ (.A1(net38),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3156_));
 sky130_fd_sc_hd__nor2_1 _7078_ (.A(_3132_),
    .B(_3156_),
    .Y(_3157_));
 sky130_fd_sc_hd__o21ai_2 _7079_ (.A1(net98),
    .A2(net71),
    .B1(_3157_),
    .Y(_3158_));
 sky130_fd_sc_hd__o221ai_4 _7080_ (.A1(_2781_),
    .A2(_2958_),
    .B1(_2962_),
    .B2(_2741_),
    .C1(_3158_),
    .Y(\dp.result2[14] ));
 sky130_fd_sc_hd__a21oi_1 _7081_ (.A1(net39),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3159_));
 sky130_fd_sc_hd__a221oi_1 _7082_ (.A1(net202),
    .A2(_2964_),
    .B1(_2969_),
    .B2(_3135_),
    .C1(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__o21a_4 _7083_ (.A1(net72),
    .A2(_3137_),
    .B1(_3160_),
    .X(\dp.result2[15] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__nor2_1 _7085_ (.A(_1806_),
    .B(_1960_),
    .Y(_3162_));
 sky130_fd_sc_hd__nand3_4 _7086_ (.A(_1813_),
    .B(net39),
    .C(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__o21ai_0 _7089_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net40),
    .Y(_3166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__a21oi_1 _7091_ (.A1(_3163_),
    .A2(_3166_),
    .B1(net273),
    .Y(_3168_));
 sky130_fd_sc_hd__nand2_1 _7092_ (.A(net202),
    .B(_2972_),
    .Y(_3169_));
 sky130_fd_sc_hd__o21ai_1 _7093_ (.A1(_3141_),
    .A2(_3168_),
    .B1(_3169_),
    .Y(_3170_));
 sky130_fd_sc_hd__nor2_1 _7094_ (.A(net73),
    .B(_3137_),
    .Y(_3171_));
 sky130_fd_sc_hd__a211oi_4 _7095_ (.A1(_3135_),
    .A2(_2976_),
    .B1(_3170_),
    .C1(_3171_),
    .Y(\dp.result2[16] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__o21ai_0 _7097_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net41),
    .Y(_3173_));
 sky130_fd_sc_hd__a21oi_1 _7098_ (.A1(_3163_),
    .A2(_3173_),
    .B1(net273),
    .Y(_3174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__o221ai_4 _7100_ (.A1(net98),
    .A2(net74),
    .B1(_3141_),
    .B2(_3174_),
    .C1(_3136_),
    .Y(_3176_));
 sky130_fd_sc_hd__o221ai_4 _7101_ (.A1(_2781_),
    .A2(_2979_),
    .B1(_2983_),
    .B2(_2741_),
    .C1(_3176_),
    .Y(\dp.result2[17] ));
 sky130_fd_sc_hd__o21ai_0 _7102_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net42),
    .Y(_3177_));
 sky130_fd_sc_hd__a21oi_1 _7103_ (.A1(_3163_),
    .A2(_3177_),
    .B1(net273),
    .Y(_3178_));
 sky130_fd_sc_hd__o221ai_4 _7104_ (.A1(net98),
    .A2(net321),
    .B1(_3141_),
    .B2(_3178_),
    .C1(_3136_),
    .Y(_3179_));
 sky130_fd_sc_hd__o221ai_4 _7105_ (.A1(_2781_),
    .A2(_2985_),
    .B1(_2988_),
    .B2(_2741_),
    .C1(net663),
    .Y(\dp.result2[18] ));
 sky130_fd_sc_hd__o21ai_0 _7106_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net43),
    .Y(_3180_));
 sky130_fd_sc_hd__a21oi_1 _7107_ (.A1(_3163_),
    .A2(_3180_),
    .B1(net273),
    .Y(_3181_));
 sky130_fd_sc_hd__nor2_1 _7108_ (.A(_3141_),
    .B(_3181_),
    .Y(_3182_));
 sky130_fd_sc_hd__nor2_1 _7109_ (.A(_3132_),
    .B(_3182_),
    .Y(_3183_));
 sky130_fd_sc_hd__o21ai_1 _7110_ (.A1(_2464_),
    .A2(_2475_),
    .B1(_1960_),
    .Y(_3184_));
 sky130_fd_sc_hd__o22ai_1 _7111_ (.A1(_2781_),
    .A2(_2990_),
    .B1(_2995_),
    .B2(_2741_),
    .Y(_3185_));
 sky130_fd_sc_hd__a21o_4 _7112_ (.A1(_3183_),
    .A2(_3184_),
    .B1(_3185_),
    .X(\dp.result2[19] ));
 sky130_fd_sc_hd__nor2_1 _7113_ (.A(net98),
    .B(_3132_),
    .Y(_3186_));
 sky130_fd_sc_hd__o22ai_1 _7114_ (.A1(_2903_),
    .A2(_2781_),
    .B1(_2741_),
    .B2(_3274_),
    .Y(_3187_));
 sky130_fd_sc_hd__a221o_4 _7115_ (.A1(net44),
    .A2(net98),
    .B1(net77),
    .B2(_3186_),
    .C1(_3187_),
    .X(\dp.result2[1] ));
 sky130_fd_sc_hd__o21ai_0 _7116_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net45),
    .Y(_3188_));
 sky130_fd_sc_hd__a21oi_1 _7117_ (.A1(_3163_),
    .A2(_3188_),
    .B1(net273),
    .Y(_3189_));
 sky130_fd_sc_hd__o221ai_4 _7118_ (.A1(net78),
    .A2(net98),
    .B1(_3141_),
    .B2(_3189_),
    .C1(_3136_),
    .Y(_3190_));
 sky130_fd_sc_hd__o221ai_4 _7119_ (.A1(_2781_),
    .A2(_3000_),
    .B1(_3004_),
    .B2(_2741_),
    .C1(net851),
    .Y(\dp.result2[20] ));
 sky130_fd_sc_hd__o21ai_0 _7120_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net46),
    .Y(_3191_));
 sky130_fd_sc_hd__a21oi_1 _7121_ (.A1(_3163_),
    .A2(_3191_),
    .B1(net273),
    .Y(_3192_));
 sky130_fd_sc_hd__o221ai_4 _7122_ (.A1(net98),
    .A2(net609),
    .B1(_3141_),
    .B2(_3192_),
    .C1(_3136_),
    .Y(_3193_));
 sky130_fd_sc_hd__o221ai_4 _7123_ (.A1(_2781_),
    .A2(_3008_),
    .B1(_3011_),
    .B2(_2741_),
    .C1(net814),
    .Y(\dp.result2[21] ));
 sky130_fd_sc_hd__o21ai_0 _7124_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net47),
    .Y(_3194_));
 sky130_fd_sc_hd__a21oi_1 _7125_ (.A1(_3163_),
    .A2(_3194_),
    .B1(net273),
    .Y(_3195_));
 sky130_fd_sc_hd__o221ai_4 _7126_ (.A1(net80),
    .A2(net98),
    .B1(_3141_),
    .B2(_3195_),
    .C1(_3136_),
    .Y(_3196_));
 sky130_fd_sc_hd__o221ai_4 _7127_ (.A1(_2781_),
    .A2(_3013_),
    .B1(_3020_),
    .B2(_2741_),
    .C1(net660),
    .Y(\dp.result2[22] ));
 sky130_fd_sc_hd__o21ai_0 _7128_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net48),
    .Y(_3197_));
 sky130_fd_sc_hd__a21oi_1 _7129_ (.A1(_3163_),
    .A2(_3197_),
    .B1(net273),
    .Y(_3198_));
 sky130_fd_sc_hd__o22ai_4 _7130_ (.A1(net625),
    .A2(net98),
    .B1(_3141_),
    .B2(_3198_),
    .Y(_3199_));
 sky130_fd_sc_hd__a22oi_2 _7131_ (.A1(_0128_),
    .A2(_3023_),
    .B1(_3031_),
    .B2(_3135_),
    .Y(_3200_));
 sky130_fd_sc_hd__a21boi_4 _7132_ (.A1(_3136_),
    .A2(net711),
    .B1_N(_3200_),
    .Y(\dp.result2[23] ));
 sky130_fd_sc_hd__nor2_1 _7133_ (.A(_2781_),
    .B(_3033_),
    .Y(_3201_));
 sky130_fd_sc_hd__a21oi_4 _7134_ (.A1(_3040_),
    .A2(_3135_),
    .B1(_3201_),
    .Y(_3202_));
 sky130_fd_sc_hd__nand2_4 _7135_ (.A(_3202_),
    .B(_1960_),
    .Y(_3203_));
 sky130_fd_sc_hd__o21ai_0 _7136_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net49),
    .Y(_3204_));
 sky130_fd_sc_hd__a21oi_1 _7137_ (.A1(_3163_),
    .A2(_3204_),
    .B1(_3140_),
    .Y(_3205_));
 sky130_fd_sc_hd__o21ai_1 _7138_ (.A1(_3141_),
    .A2(_3205_),
    .B1(_3136_),
    .Y(_3206_));
 sky130_fd_sc_hd__a2bb2oi_4 _7139_ (.A1_N(net301),
    .A2_N(_3203_),
    .B1(_3206_),
    .B2(_3202_),
    .Y(\dp.result2[24] ));
 sky130_fd_sc_hd__o21ai_1 _7140_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net50),
    .Y(_3207_));
 sky130_fd_sc_hd__a21oi_4 _7141_ (.A1(_3163_),
    .A2(_3207_),
    .B1(net273),
    .Y(_3208_));
 sky130_fd_sc_hd__nor2_1 _7142_ (.A(_3141_),
    .B(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__a221oi_1 _7143_ (.A1(_0128_),
    .A2(_3044_),
    .B1(_3050_),
    .B2(_3135_),
    .C1(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__o21a_4 _7144_ (.A1(_3137_),
    .A2(net617),
    .B1(_3210_),
    .X(\dp.result2[25] ));
 sky130_fd_sc_hd__o21ai_4 _7145_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net51),
    .Y(_3211_));
 sky130_fd_sc_hd__a21oi_1 _7146_ (.A1(_3163_),
    .A2(_3211_),
    .B1(_3140_),
    .Y(_3212_));
 sky130_fd_sc_hd__nand2_1 _7147_ (.A(_0128_),
    .B(_3053_),
    .Y(_3213_));
 sky130_fd_sc_hd__o221ai_4 _7148_ (.A1(_3137_),
    .A2(net284),
    .B1(_3141_),
    .B2(_3212_),
    .C1(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__a21oi_4 _7149_ (.A1(_3135_),
    .A2(_3058_),
    .B1(net607),
    .Y(\dp.result2[26] ));
 sky130_fd_sc_hd__o22ai_2 _7150_ (.A1(_2781_),
    .A2(_3060_),
    .B1(_3066_),
    .B2(_2741_),
    .Y(_3215_));
 sky130_fd_sc_hd__o21ai_0 _7151_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net52),
    .Y(_3216_));
 sky130_fd_sc_hd__a21oi_1 _7152_ (.A1(_3163_),
    .A2(_3216_),
    .B1(_3140_),
    .Y(_3217_));
 sky130_fd_sc_hd__o21ai_0 _7153_ (.A1(_3141_),
    .A2(_3217_),
    .B1(_3136_),
    .Y(_3218_));
 sky130_fd_sc_hd__nand2b_1 _7154_ (.A_N(_3215_),
    .B(_3218_),
    .Y(_3219_));
 sky130_fd_sc_hd__o31a_4 _7155_ (.A1(net98),
    .A2(_3215_),
    .A3(net85),
    .B1(_3219_),
    .X(\dp.result2[27] ));
 sky130_fd_sc_hd__o21ai_0 _7156_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net53),
    .Y(_3220_));
 sky130_fd_sc_hd__a21oi_1 _7157_ (.A1(_3163_),
    .A2(_3220_),
    .B1(_3140_),
    .Y(_3221_));
 sky130_fd_sc_hd__o221ai_4 _7158_ (.A1(net98),
    .A2(net280),
    .B1(_3141_),
    .B2(_3221_),
    .C1(_3136_),
    .Y(_3222_));
 sky130_fd_sc_hd__o221ai_4 _7159_ (.A1(_2781_),
    .A2(_3068_),
    .B1(_3075_),
    .B2(_2741_),
    .C1(_3222_),
    .Y(\dp.result2[28] ));
 sky130_fd_sc_hd__o21ai_0 _7160_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net54),
    .Y(_3223_));
 sky130_fd_sc_hd__a21oi_1 _7161_ (.A1(_3163_),
    .A2(_3223_),
    .B1(_3140_),
    .Y(_3224_));
 sky130_fd_sc_hd__o21ai_2 _7162_ (.A1(_3141_),
    .A2(_3224_),
    .B1(_3136_),
    .Y(_3225_));
 sky130_fd_sc_hd__nor2_1 _7163_ (.A(_2741_),
    .B(_3082_),
    .Y(_3226_));
 sky130_fd_sc_hd__o22ai_1 _7164_ (.A1(_2781_),
    .A2(_3077_),
    .B1(_3225_),
    .B2(_1960_),
    .Y(_3227_));
 sky130_fd_sc_hd__nor2_4 _7165_ (.A(_3226_),
    .B(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hd__o21ai_4 _7166_ (.A1(net420),
    .A2(_3225_),
    .B1(_3228_),
    .Y(\dp.result2[29] ));
 sky130_fd_sc_hd__a22oi_1 _7167_ (.A1(net122),
    .A2(net202),
    .B1(_3135_),
    .B2(_3084_),
    .Y(_3229_));
 sky130_fd_sc_hd__o221a_4 _7168_ (.A1(net55),
    .A2(_1960_),
    .B1(net88),
    .B2(_3137_),
    .C1(_3229_),
    .X(\dp.result2[2] ));
 sky130_fd_sc_hd__o21ai_1 _7169_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net56),
    .Y(_3230_));
 sky130_fd_sc_hd__a21oi_4 _7170_ (.A1(_3163_),
    .A2(_3230_),
    .B1(net273),
    .Y(_3231_));
 sky130_fd_sc_hd__o21ai_2 _7171_ (.A1(_3141_),
    .A2(_3231_),
    .B1(_3136_),
    .Y(_3232_));
 sky130_fd_sc_hd__a21oi_4 _7172_ (.A1(net275),
    .A2(_2692_),
    .B1(net98),
    .Y(_3233_));
 sky130_fd_sc_hd__o21ai_4 _7173_ (.A1(_3090_),
    .A2(_3094_),
    .B1(_3135_),
    .Y(_3234_));
 sky130_fd_sc_hd__o221ai_4 _7174_ (.A1(_2781_),
    .A2(_3087_),
    .B1(_3232_),
    .B2(net530),
    .C1(_3234_),
    .Y(\dp.result2[30] ));
 sky130_fd_sc_hd__o21ai_0 _7175_ (.A1(_1806_),
    .A2(_1960_),
    .B1(net57),
    .Y(_3235_));
 sky130_fd_sc_hd__a21oi_1 _7176_ (.A1(_3163_),
    .A2(_3235_),
    .B1(net273),
    .Y(_3236_));
 sky130_fd_sc_hd__or2_2 _7177_ (.A(_3141_),
    .B(_3236_),
    .X(_3237_));
 sky130_fd_sc_hd__and3_1 _7178_ (.A(_1818_),
    .B(_2721_),
    .C(_3237_),
    .X(_3238_));
 sky130_fd_sc_hd__o31ai_1 _7179_ (.A1(_2701_),
    .A2(_2707_),
    .A3(_2709_),
    .B1(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__and3_1 _7180_ (.A(_2714_),
    .B(_2721_),
    .C(_3237_),
    .X(_3240_));
 sky130_fd_sc_hd__a21oi_1 _7181_ (.A1(net98),
    .A2(_3237_),
    .B1(_3240_),
    .Y(_3241_));
 sky130_fd_sc_hd__and3_4 _7182_ (.A(_3136_),
    .B(_3241_),
    .C(_3239_),
    .X(_3242_));
 sky130_fd_sc_hd__a221oi_4 _7183_ (.A1(_0128_),
    .A2(_3097_),
    .B1(_3103_),
    .B2(_3135_),
    .C1(_3242_),
    .Y(\dp.result2[31] ));
 sky130_fd_sc_hd__nand2_1 _7184_ (.A(_1960_),
    .B(net91),
    .Y(_3243_));
 sky130_fd_sc_hd__a21oi_1 _7185_ (.A1(net58),
    .A2(net98),
    .B1(_3132_),
    .Y(_3244_));
 sky130_fd_sc_hd__o22ai_2 _7186_ (.A1(_3543_),
    .A2(_2781_),
    .B1(_2741_),
    .B2(_3104_),
    .Y(_3245_));
 sky130_fd_sc_hd__a21oi_4 _7187_ (.A1(_3243_),
    .A2(_3244_),
    .B1(_3245_),
    .Y(\dp.result2[3] ));
 sky130_fd_sc_hd__mux2_1 _7188_ (.A0(net59),
    .A1(net92),
    .S(_1960_),
    .X(_3246_));
 sky130_fd_sc_hd__o22ai_2 _7189_ (.A1(_2781_),
    .A2(_3105_),
    .B1(_3106_),
    .B2(_2741_),
    .Y(_3247_));
 sky130_fd_sc_hd__a21o_4 _7190_ (.A1(_3136_),
    .A2(_3246_),
    .B1(_3247_),
    .X(\dp.result2[4] ));
 sky130_fd_sc_hd__a22oi_2 _7191_ (.A1(net202),
    .A2(_3108_),
    .B1(_3110_),
    .B2(_3135_),
    .Y(_3248_));
 sky130_fd_sc_hd__o221a_4 _7192_ (.A1(net60),
    .A2(_1960_),
    .B1(net93),
    .B2(_3137_),
    .C1(_3248_),
    .X(\dp.result2[5] ));
 sky130_fd_sc_hd__mux2i_4 _7193_ (.A0(net61),
    .A1(net613),
    .S(_1960_),
    .Y(_3249_));
 sky130_fd_sc_hd__a22oi_1 _7194_ (.A1(net202),
    .A2(_3112_),
    .B1(_3115_),
    .B2(_3135_),
    .Y(_3250_));
 sky130_fd_sc_hd__a21boi_4 _7195_ (.A1(_3249_),
    .A2(_3136_),
    .B1_N(_3250_),
    .Y(\dp.result2[6] ));
 sky130_fd_sc_hd__and2_0 _7196_ (.A(net62),
    .B(net98),
    .X(_3251_));
 sky130_fd_sc_hd__a211oi_4 _7197_ (.A1(_1960_),
    .A2(net493),
    .B1(_3132_),
    .C1(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__a221oi_4 _7198_ (.A1(net202),
    .A2(_3117_),
    .B1(_3120_),
    .B2(_3135_),
    .C1(_3252_),
    .Y(\dp.result2[7] ));
 sky130_fd_sc_hd__a21oi_1 _7199_ (.A1(net63),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3253_));
 sky130_fd_sc_hd__nor2_1 _7200_ (.A(_3132_),
    .B(_3253_),
    .Y(_3254_));
 sky130_fd_sc_hd__o21ai_2 _7201_ (.A1(net98),
    .A2(net96),
    .B1(_3254_),
    .Y(_3255_));
 sky130_fd_sc_hd__o221ai_4 _7202_ (.A1(_2781_),
    .A2(_3121_),
    .B1(_3123_),
    .B2(_2741_),
    .C1(_3255_),
    .Y(\dp.result2[8] ));
 sky130_fd_sc_hd__a21oi_1 _7203_ (.A1(net64),
    .A2(_3139_),
    .B1(_3141_),
    .Y(_3256_));
 sky130_fd_sc_hd__nor2_1 _7204_ (.A(_3132_),
    .B(_3256_),
    .Y(_3257_));
 sky130_fd_sc_hd__o21ai_2 _7205_ (.A1(net98),
    .A2(net97),
    .B1(_3257_),
    .Y(_3258_));
 sky130_fd_sc_hd__o221ai_4 _7206_ (.A1(_2781_),
    .A2(_3125_),
    .B1(_3128_),
    .B2(_2741_),
    .C1(_3258_),
    .Y(\dp.result2[9] ));
 sky130_fd_sc_hd__and4_1 _7207_ (.A(net27),
    .B(net28),
    .C(net29),
    .D(_0041_),
    .X(net132));
 sky130_fd_sc_hd__nand3_2 _7208_ (.A(net99),
    .B(_0109_),
    .C(_1805_),
    .Y(_3259_));
 sky130_fd_sc_hd__and2_0 _7209_ (.A(_1378_),
    .B(_3259_),
    .X(net134));
 sky130_fd_sc_hd__and3_2 _7210_ (.A(net99),
    .B(_0109_),
    .C(_1805_),
    .X(_3260_));
 sky130_fd_sc_hd__nor3_2 _7211_ (.A(_0401_),
    .B(_1340_),
    .C(_3260_),
    .Y(net135));
 sky130_fd_sc_hd__nor2_2 _7212_ (.A(_1299_),
    .B(_3260_),
    .Y(net136));
 sky130_fd_sc_hd__and2_0 _7213_ (.A(_1264_),
    .B(_3259_),
    .X(net137));
 sky130_fd_sc_hd__and2_0 _7214_ (.A(_1218_),
    .B(_3259_),
    .X(net138));
 sky130_fd_sc_hd__nor2_2 _7215_ (.A(_1174_),
    .B(_3260_),
    .Y(net139));
 sky130_fd_sc_hd__nor2b_4 _7216_ (.A(net5),
    .B_N(net99),
    .Y(_3261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__nor2_1 _7219_ (.A(_1127_),
    .B(_3261_),
    .Y(net140));
 sky130_fd_sc_hd__nor2_1 _7220_ (.A(_1060_),
    .B(_3261_),
    .Y(net141));
 sky130_fd_sc_hd__nor2_1 _7221_ (.A(_1002_),
    .B(_3261_),
    .Y(net142));
 sky130_fd_sc_hd__inv_1 _7222_ (.A(_0950_),
    .Y(_3264_));
 sky130_fd_sc_hd__nor2_1 _7223_ (.A(_3264_),
    .B(_3261_),
    .Y(net143));
 sky130_fd_sc_hd__nor2_2 _7224_ (.A(_0881_),
    .B(_3261_),
    .Y(net145));
 sky130_fd_sc_hd__nor2_2 _7225_ (.A(_0838_),
    .B(_3261_),
    .Y(net146));
 sky130_fd_sc_hd__nor2_2 _7226_ (.A(_0794_),
    .B(_3261_),
    .Y(net147));
 sky130_fd_sc_hd__nor3_2 _7227_ (.A(_0401_),
    .B(_0747_),
    .C(_3261_),
    .Y(net148));
 sky130_fd_sc_hd__nor2_2 _7228_ (.A(_0694_),
    .B(_3261_),
    .Y(net149));
 sky130_fd_sc_hd__nor2_2 _7229_ (.A(_0636_),
    .B(_3261_),
    .Y(net150));
 sky130_fd_sc_hd__nor2_2 _7230_ (.A(_0571_),
    .B(_3261_),
    .Y(net151));
 sky130_fd_sc_hd__nor2_2 _7231_ (.A(_0516_),
    .B(_3261_),
    .Y(net152));
 sky130_fd_sc_hd__nor2_2 _7232_ (.A(_0458_),
    .B(_3261_),
    .Y(net153));
 sky130_fd_sc_hd__nor3_2 _7233_ (.A(_0383_),
    .B(_0403_),
    .C(_3261_),
    .Y(net154));
 sky130_fd_sc_hd__nor2_1 _7234_ (.A(_0324_),
    .B(_3261_),
    .Y(net156));
 sky130_fd_sc_hd__nor2_2 _7235_ (.A(_0298_),
    .B(_3261_),
    .Y(net157));
 sky130_fd_sc_hd__nor2_1 _7236_ (.A(_1455_),
    .B(_3260_),
    .Y(net163));
 sky130_fd_sc_hd__nor2_1 _7237_ (.A(_1419_),
    .B(_3260_),
    .Y(net164));
 sky130_fd_sc_hd__fa_2 _7238_ (.A(_3266_),
    .B(_3265_),
    .CIN(_3267_),
    .COUT(_3268_),
    .SUM(_3269_));
 sky130_fd_sc_hd__fa_2 _7239_ (.A(_3270_),
    .B(_3271_),
    .CIN(_3272_),
    .COUT(_3273_),
    .SUM(_3274_));
 sky130_fd_sc_hd__ha_1 _7240_ (.A(_3275_),
    .B(_3276_),
    .COUT(_3277_),
    .SUM(_3278_));
 sky130_fd_sc_hd__ha_1 _7241_ (.A(net498),
    .B(_3280_),
    .COUT(_3281_),
    .SUM(_3282_));
 sky130_fd_sc_hd__ha_1 _7242_ (.A(_3283_),
    .B(_3284_),
    .COUT(_3285_),
    .SUM(_3286_));
 sky130_fd_sc_hd__ha_1 _7243_ (.A(_3287_),
    .B(_0274_),
    .COUT(_3289_),
    .SUM(_3290_));
 sky130_fd_sc_hd__ha_1 _7244_ (.A(_3291_),
    .B(_3292_),
    .COUT(_3293_),
    .SUM(_3294_));
 sky130_fd_sc_hd__ha_1 _7245_ (.A(_0371_),
    .B(_3296_),
    .COUT(_3297_),
    .SUM(_3298_));
 sky130_fd_sc_hd__ha_2 _7246_ (.A(_3299_),
    .B(_3300_),
    .COUT(_3301_),
    .SUM(_3302_));
 sky130_fd_sc_hd__ha_1 _7247_ (.A(_3303_),
    .B(_3304_),
    .COUT(_3305_),
    .SUM(_3306_));
 sky130_fd_sc_hd__ha_2 _7248_ (.A(_3307_),
    .B(_3308_),
    .COUT(_3309_),
    .SUM(_3310_));
 sky130_fd_sc_hd__ha_1 _7249_ (.A(_3311_),
    .B(_3312_),
    .COUT(_3313_),
    .SUM(_3314_));
 sky130_fd_sc_hd__ha_1 _7250_ (.A(_3315_),
    .B(_3316_),
    .COUT(_3317_),
    .SUM(_3318_));
 sky130_fd_sc_hd__ha_1 _7251_ (.A(_3319_),
    .B(_3320_),
    .COUT(_3321_),
    .SUM(_3322_));
 sky130_fd_sc_hd__ha_1 _7252_ (.A(_3323_),
    .B(_3324_),
    .COUT(_3325_),
    .SUM(_3326_));
 sky130_fd_sc_hd__ha_1 _7253_ (.A(_0621_),
    .B(_3328_),
    .COUT(_3329_),
    .SUM(_3330_));
 sky130_fd_sc_hd__ha_1 _7254_ (.A(_3331_),
    .B(_3332_),
    .COUT(_3333_),
    .SUM(_3334_));
 sky130_fd_sc_hd__ha_1 _7255_ (.A(_3335_),
    .B(_3336_),
    .COUT(_3337_),
    .SUM(_3338_));
 sky130_fd_sc_hd__ha_2 _7256_ (.A(_3339_),
    .B(_3340_),
    .COUT(_3341_),
    .SUM(_3342_));
 sky130_fd_sc_hd__ha_1 _7257_ (.A(_3343_),
    .B(_3344_),
    .COUT(_3345_),
    .SUM(_3346_));
 sky130_fd_sc_hd__ha_1 _7258_ (.A(_3347_),
    .B(_3348_),
    .COUT(_3349_),
    .SUM(_3350_));
 sky130_fd_sc_hd__ha_1 _7259_ (.A(_3351_),
    .B(_3352_),
    .COUT(_3353_),
    .SUM(_3354_));
 sky130_fd_sc_hd__ha_2 _7260_ (.A(_3355_),
    .B(_3356_),
    .COUT(_3357_),
    .SUM(_3358_));
 sky130_fd_sc_hd__ha_1 _7261_ (.A(_3359_),
    .B(_3360_),
    .COUT(_3361_),
    .SUM(_3362_));
 sky130_fd_sc_hd__ha_2 _7262_ (.A(_3363_),
    .B(_3364_),
    .COUT(_3365_),
    .SUM(_3366_));
 sky130_fd_sc_hd__ha_1 _7263_ (.A(_3367_),
    .B(_3368_),
    .COUT(_3369_),
    .SUM(_3370_));
 sky130_fd_sc_hd__ha_1 _7264_ (.A(_3371_),
    .B(_3372_),
    .COUT(_3373_),
    .SUM(_3374_));
 sky130_fd_sc_hd__ha_1 _7265_ (.A(_3375_),
    .B(_3376_),
    .COUT(_3377_),
    .SUM(_3378_));
 sky130_fd_sc_hd__ha_1 _7266_ (.A(_3379_),
    .B(_3380_),
    .COUT(_3381_),
    .SUM(_3382_));
 sky130_fd_sc_hd__ha_1 _7267_ (.A(_3383_),
    .B(_3384_),
    .COUT(_3385_),
    .SUM(_3386_));
 sky130_fd_sc_hd__ha_2 _7268_ (.A(_3387_),
    .B(_3388_),
    .COUT(_3389_),
    .SUM(_3390_));
 sky130_fd_sc_hd__ha_1 _7269_ (.A(_1031_),
    .B(_3392_),
    .COUT(_3393_),
    .SUM(_3394_));
 sky130_fd_sc_hd__ha_2 _7270_ (.A(_3395_),
    .B(_3396_),
    .COUT(_3397_),
    .SUM(_3398_));
 sky130_fd_sc_hd__ha_1 _7271_ (.A(_3399_),
    .B(_3400_),
    .COUT(_3401_),
    .SUM(_3402_));
 sky130_fd_sc_hd__ha_2 _7272_ (.A(_3403_),
    .B(_3404_),
    .COUT(_3405_),
    .SUM(_3406_));
 sky130_fd_sc_hd__ha_1 _7273_ (.A(_3407_),
    .B(_3408_),
    .COUT(_3409_),
    .SUM(_3410_));
 sky130_fd_sc_hd__ha_2 _7274_ (.A(_3411_),
    .B(_3412_),
    .COUT(_3413_),
    .SUM(_3414_));
 sky130_fd_sc_hd__ha_1 _7275_ (.A(_3415_),
    .B(_3416_),
    .COUT(_3417_),
    .SUM(_3418_));
 sky130_fd_sc_hd__ha_2 _7276_ (.A(_3419_),
    .B(_3420_),
    .COUT(_3421_),
    .SUM(_3422_));
 sky130_fd_sc_hd__ha_1 _7277_ (.A(_3423_),
    .B(_3424_),
    .COUT(_3425_),
    .SUM(_3426_));
 sky130_fd_sc_hd__ha_2 _7278_ (.A(_3427_),
    .B(_3428_),
    .COUT(_3429_),
    .SUM(_3430_));
 sky130_fd_sc_hd__ha_1 _7279_ (.A(_3431_),
    .B(_3432_),
    .COUT(_3433_),
    .SUM(_3434_));
 sky130_fd_sc_hd__ha_2 _7280_ (.A(_3435_),
    .B(_3436_),
    .COUT(_3437_),
    .SUM(_3438_));
 sky130_fd_sc_hd__ha_1 _7281_ (.A(_3439_),
    .B(_3440_),
    .COUT(_3441_),
    .SUM(_3442_));
 sky130_fd_sc_hd__ha_2 _7282_ (.A(_3443_),
    .B(_3444_),
    .COUT(_3445_),
    .SUM(_3446_));
 sky130_fd_sc_hd__ha_1 _7283_ (.A(_3447_),
    .B(_3448_),
    .COUT(_3449_),
    .SUM(_3450_));
 sky130_fd_sc_hd__ha_2 _7284_ (.A(_3451_),
    .B(_3452_),
    .COUT(_3453_),
    .SUM(_3454_));
 sky130_fd_sc_hd__ha_1 _7285_ (.A(_3455_),
    .B(_3456_),
    .COUT(_3457_),
    .SUM(_3458_));
 sky130_fd_sc_hd__ha_2 _7286_ (.A(_3459_),
    .B(_3460_),
    .COUT(_3461_),
    .SUM(_3462_));
 sky130_fd_sc_hd__ha_1 _7287_ (.A(net852),
    .B(_3464_),
    .COUT(_3465_),
    .SUM(_3466_));
 sky130_fd_sc_hd__ha_2 _7288_ (.A(_3467_),
    .B(_3468_),
    .COUT(_3469_),
    .SUM(_3470_));
 sky130_fd_sc_hd__ha_1 _7289_ (.A(_3471_),
    .B(_3472_),
    .COUT(_3473_),
    .SUM(_3474_));
 sky130_fd_sc_hd__ha_2 _7290_ (.A(_3475_),
    .B(_3476_),
    .COUT(_3477_),
    .SUM(_3478_));
 sky130_fd_sc_hd__ha_1 _7291_ (.A(_3479_),
    .B(_3480_),
    .COUT(_3481_),
    .SUM(_3482_));
 sky130_fd_sc_hd__ha_2 _7292_ (.A(_3483_),
    .B(_3484_),
    .COUT(_3485_),
    .SUM(_3486_));
 sky130_fd_sc_hd__ha_1 _7293_ (.A(net515),
    .B(_3488_),
    .COUT(_3489_),
    .SUM(_3490_));
 sky130_fd_sc_hd__ha_1 _7294_ (.A(_3491_),
    .B(_3492_),
    .COUT(_3493_),
    .SUM(_3494_));
 sky130_fd_sc_hd__ha_1 _7295_ (.A(_3495_),
    .B(_3496_),
    .COUT(_3497_),
    .SUM(_3498_));
 sky130_fd_sc_hd__ha_2 _7296_ (.A(_3499_),
    .B(_3500_),
    .COUT(_3501_),
    .SUM(_3502_));
 sky130_fd_sc_hd__ha_1 _7297_ (.A(_3503_),
    .B(_3504_),
    .COUT(_3505_),
    .SUM(_3506_));
 sky130_fd_sc_hd__ha_1 _7298_ (.A(_3508_),
    .B(_3507_),
    .COUT(_3509_),
    .SUM(_3510_));
 sky130_fd_sc_hd__ha_1 _7299_ (.A(_1689_),
    .B(_3512_),
    .COUT(_3513_),
    .SUM(_3514_));
 sky130_fd_sc_hd__ha_1 _7300_ (.A(_3516_),
    .B(_3515_),
    .COUT(_3517_),
    .SUM(_3518_));
 sky130_fd_sc_hd__ha_1 _7301_ (.A(_3519_),
    .B(_3520_),
    .COUT(_3521_),
    .SUM(_3522_));
 sky130_fd_sc_hd__ha_1 _7302_ (.A(_3266_),
    .B(_3267_),
    .COUT(_3523_),
    .SUM(_3524_));
 sky130_fd_sc_hd__ha_1 _7303_ (.A(_3525_),
    .B(_3526_),
    .COUT(_3527_),
    .SUM(_3528_));
 sky130_fd_sc_hd__ha_2 _7304_ (.A(_3529_),
    .B(_3530_),
    .COUT(_3270_),
    .SUM(_3531_));
 sky130_fd_sc_hd__ha_1 _7305_ (.A(_3271_),
    .B(_3272_),
    .COUT(_3532_),
    .SUM(_3533_));
 sky130_fd_sc_hd__ha_1 _7306_ (.A(_3534_),
    .B(_3535_),
    .COUT(_3536_),
    .SUM(_3537_));
 sky130_fd_sc_hd__ha_1 _7307_ (.A(_3538_),
    .B(_3539_),
    .COUT(_3540_),
    .SUM(_3541_));
 sky130_fd_sc_hd__ha_2 _7308_ (.A(net122),
    .B(net125),
    .COUT(_3542_),
    .SUM(_3543_));
 sky130_fd_sc_hd__ha_1 _7309_ (.A(_3544_),
    .B(_3545_),
    .COUT(_3546_),
    .SUM(_3547_));
 sky130_fd_sc_hd__ha_1 _7310_ (.A(_3548_),
    .B(_3549_),
    .COUT(_3550_),
    .SUM(_3551_));
 sky130_fd_sc_hd__ha_1 _7311_ (.A(_3552_),
    .B(_3553_),
    .COUT(_3554_),
    .SUM(_3555_));
 sky130_fd_sc_hd__ha_1 _7312_ (.A(_3556_),
    .B(_3557_),
    .COUT(_3558_),
    .SUM(_3559_));
 sky130_fd_sc_hd__ha_1 _7313_ (.A(_3560_),
    .B(_3561_),
    .COUT(_3562_),
    .SUM(_3563_));
 sky130_fd_sc_hd__ha_1 _7314_ (.A(_3564_),
    .B(_3565_),
    .COUT(_3566_),
    .SUM(_3567_));
 sky130_fd_sc_hd__ha_1 _7315_ (.A(_3568_),
    .B(_3569_),
    .COUT(_3570_),
    .SUM(_3571_));
 sky130_fd_sc_hd__ha_1 _7316_ (.A(_3572_),
    .B(_3573_),
    .COUT(_3574_),
    .SUM(_3575_));
 sky130_fd_sc_hd__ha_1 _7317_ (.A(_3576_),
    .B(_3577_),
    .COUT(_3578_),
    .SUM(_3579_));
 sky130_fd_sc_hd__ha_2 _7318_ (.A(_3580_),
    .B(_3581_),
    .COUT(_3582_),
    .SUM(_3583_));
 sky130_fd_sc_hd__ha_2 _7319_ (.A(_3584_),
    .B(_3585_),
    .COUT(_3586_),
    .SUM(_3587_));
 sky130_fd_sc_hd__ha_1 _7320_ (.A(_3588_),
    .B(_3589_),
    .COUT(_3590_),
    .SUM(_3591_));
 sky130_fd_sc_hd__ha_2 _7321_ (.A(_3592_),
    .B(_3593_),
    .COUT(_3594_),
    .SUM(_3595_));
 sky130_fd_sc_hd__ha_2 _7322_ (.A(_3596_),
    .B(_3597_),
    .COUT(_3598_),
    .SUM(_3599_));
 sky130_fd_sc_hd__ha_2 _7323_ (.A(_3600_),
    .B(_3601_),
    .COUT(_3602_),
    .SUM(_3603_));
 sky130_fd_sc_hd__ha_2 _7324_ (.A(_3604_),
    .B(_3605_),
    .COUT(_3606_),
    .SUM(_3607_));
 sky130_fd_sc_hd__ha_1 _7325_ (.A(_3608_),
    .B(_3609_),
    .COUT(_3610_),
    .SUM(_3611_));
 sky130_fd_sc_hd__ha_2 _7326_ (.A(_3612_),
    .B(_3613_),
    .COUT(_3614_),
    .SUM(_3615_));
 sky130_fd_sc_hd__ha_1 _7327_ (.A(_3616_),
    .B(_3617_),
    .COUT(_3618_),
    .SUM(_3619_));
 sky130_fd_sc_hd__ha_1 _7328_ (.A(_3620_),
    .B(_3621_),
    .COUT(_3622_),
    .SUM(_3623_));
 sky130_fd_sc_hd__ha_1 _7329_ (.A(_3624_),
    .B(_3625_),
    .COUT(_3626_),
    .SUM(_3627_));
 sky130_fd_sc_hd__ha_1 _7330_ (.A(_3628_),
    .B(_3629_),
    .COUT(_3630_),
    .SUM(_3631_));
 sky130_fd_sc_hd__ha_2 _7331_ (.A(_3632_),
    .B(_3633_),
    .COUT(_3634_),
    .SUM(_3635_));
 sky130_fd_sc_hd__ha_1 _7332_ (.A(_3636_),
    .B(_3637_),
    .COUT(_3638_),
    .SUM(_3639_));
 sky130_fd_sc_hd__ha_1 _7333_ (.A(_3640_),
    .B(_3641_),
    .COUT(_3642_),
    .SUM(_3643_));
 sky130_fd_sc_hd__ha_1 _7334_ (.A(_3644_),
    .B(_3645_),
    .COUT(_3646_),
    .SUM(_3647_));
 sky130_fd_sc_hd__ha_1 _7335_ (.A(_3648_),
    .B(_3649_),
    .COUT(_3650_),
    .SUM(_3651_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[0]$_DFFE_PP0P_  (.D(_0032_),
    .Q(net100),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[10]$_DFF_PP0_  (.D(\dp.ISRmux.d0[10] ),
    .Q(net101),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[11]$_DFF_PP0_  (.D(\dp.ISRmux.d0[11] ),
    .Q(net102),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[12]$_DFF_PP0_  (.D(\dp.ISRmux.d0[12] ),
    .Q(net103),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[13]$_DFF_PP0_  (.D(\dp.ISRmux.d0[13] ),
    .Q(net104),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[14]$_DFF_PP0_  (.D(\dp.ISRmux.d0[14] ),
    .Q(net105),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[15]$_DFF_PP0_  (.D(\dp.ISRmux.d0[15] ),
    .Q(net106),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[16]$_DFF_PP0_  (.D(\dp.ISRmux.d0[16] ),
    .Q(net107),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[17]$_DFF_PP0_  (.D(\dp.ISRmux.d0[17] ),
    .Q(net108),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[18]$_DFF_PP0_  (.D(\dp.ISRmux.d0[18] ),
    .Q(net109),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[19]$_DFF_PP0_  (.D(\dp.ISRmux.d0[19] ),
    .Q(net110),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \dp.pcreg.q[1]$_DFFE_PP0P_  (.D(_0033_),
    .Q(net111),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[20]$_DFF_PP0_  (.D(\dp.ISRmux.d0[20] ),
    .Q(net112),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[21]$_DFF_PP0_  (.D(\dp.ISRmux.d0[21] ),
    .Q(net113),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[22]$_DFF_PP0_  (.D(\dp.ISRmux.d0[22] ),
    .Q(net114),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[23]$_DFF_PP0_  (.D(\dp.ISRmux.d0[23] ),
    .Q(net115),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[24]$_DFF_PP0_  (.D(\dp.ISRmux.d0[24] ),
    .Q(net116),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[25]$_DFF_PP0_  (.D(\dp.ISRmux.d0[25] ),
    .Q(net117),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[26]$_DFF_PP0_  (.D(\dp.ISRmux.d0[26] ),
    .Q(net118),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[27]$_DFF_PP0_  (.D(\dp.ISRmux.d0[27] ),
    .Q(net119),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[28]$_DFF_PP0_  (.D(\dp.ISRmux.d0[28] ),
    .Q(net120),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[29]$_DFF_PP0_  (.D(\dp.ISRmux.d0[29] ),
    .Q(net121),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[2]$_DFF_PP0_  (.D(\dp.ISRmux.d0[2] ),
    .Q(net122),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[30]$_DFF_PP0_  (.D(\dp.ISRmux.d0[30] ),
    .Q(net123),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[31]$_DFF_PP0_  (.D(\dp.ISRmux.d0[31] ),
    .Q(net124),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[3]$_DFF_PP0_  (.D(\dp.ISRmux.d0[3] ),
    .Q(net125),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[4]$_DFF_PP0_  (.D(\dp.ISRmux.d0[4] ),
    .Q(net126),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_2 \dp.pcreg.q[5]$_DFF_PP0_  (.D(\dp.ISRmux.d0[5] ),
    .Q(net127),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \dp.pcreg.q[6]$_DFF_PP0_  (.D(\dp.ISRmux.d0[6] ),
    .Q(net128),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[7]$_DFF_PP0_  (.D(\dp.ISRmux.d0[7] ),
    .Q(net129),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[8]$_DFF_PP0_  (.D(\dp.ISRmux.d0[8] ),
    .Q(net130),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[9]$_DFF_PP0_  (.D(\dp.ISRmux.d0[9] ),
    .Q(net131),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][0]$_DFFE_PP_  (.D(net309),
    .DE(net216),
    .Q(\dp.rf.rf[0][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net217),
    .Q(\dp.rf.rf[0][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(net218),
    .Q(\dp.rf.rf[0][11] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][12]$_DFFE_PP_  (.D(net638),
    .DE(net219),
    .Q(\dp.rf.rf[0][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net220),
    .Q(\dp.rf.rf[0][13] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net221),
    .Q(\dp.rf.rf[0][14] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net222),
    .Q(\dp.rf.rf[0][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][18]$_DFFE_PP_  (.D(net661),
    .DE(net223),
    .Q(\dp.rf.rf[0][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(net224),
    .Q(\dp.rf.rf[0][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net225),
    .Q(\dp.rf.rf[0][1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][20]$_DFFE_PP_  (.D(net850),
    .DE(net226),
    .Q(\dp.rf.rf[0][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][21]$_DFFE_PP_  (.D(net742),
    .DE(net227),
    .Q(\dp.rf.rf[0][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][22]$_DFFE_PP_  (.D(net649),
    .DE(net228),
    .Q(\dp.rf.rf[0][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][23]$_DFFE_PP_  (.D(net614),
    .DE(net229),
    .Q(\dp.rf.rf[0][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][24]$_DFFE_PP_  (.D(net678),
    .DE(net230),
    .Q(\dp.rf.rf[0][24] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][25]$_DFFE_PP_  (.D(net931),
    .DE(net231),
    .Q(\dp.rf.rf[0][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][26]$_DFFE_PP_  (.D(net608),
    .DE(net232),
    .Q(\dp.rf.rf[0][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(net233),
    .Q(\dp.rf.rf[0][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net234),
    .Q(\dp.rf.rf[0][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][29]$_DFFE_PP_  (.D(net734),
    .DE(net235),
    .Q(\dp.rf.rf[0][29] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net236),
    .Q(\dp.rf.rf[0][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][30]$_DFFE_PP_  (.D(net474),
    .DE(net237),
    .Q(\dp.rf.rf[0][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][31]$_DFFE_PP_  (.D(net524),
    .DE(net238),
    .Q(\dp.rf.rf[0][31] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net239),
    .Q(\dp.rf.rf[0][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net240),
    .Q(\dp.rf.rf[0][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net241),
    .Q(\dp.rf.rf[0][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(net242),
    .Q(\dp.rf.rf[0][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][7]$_DFFE_PP_  (.D(net272),
    .DE(net243),
    .Q(\dp.rf.rf[0][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net244),
    .Q(\dp.rf.rf[0][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net245),
    .Q(\dp.rf.rf[0][9] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][13] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][16]$_DFFE_PP_  (.D(net933),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][17]$_DFFE_PP_  (.D(net934),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][18]$_DFFE_PP_  (.D(net736),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][19] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][20] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][22]$_DFFE_PP_  (.D(net650),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][23]$_DFFE_PP_  (.D(net614),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][23] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][24]$_DFFE_PP_  (.D(net735),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][24] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][25] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][28]$_DFFE_PP_  (.D(net635),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][29]$_DFFE_PP_  (.D(net734),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][29] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][30]$_DFFE_PP_  (.D(net475),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][31]$_DFFE_PP_  (.D(net688),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][3] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][7]$_DFFE_PP_  (.D(net272),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][8] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][13] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][16]$_DFFE_PP_  (.D(net933),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][17]$_DFFE_PP_  (.D(net934),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][18]$_DFFE_PP_  (.D(net736),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][20] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][22] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][23]$_DFFE_PP_  (.D(net614),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][23] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][24]$_DFFE_PP_  (.D(net733),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][25] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][28]$_DFFE_PP_  (.D(net635),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][29]$_DFFE_PP_  (.D(net712),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][30]$_DFFE_PP_  (.D(net475),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][31]$_DFFE_PP_  (.D(net688),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][7]$_DFFE_PP_  (.D(net272),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][0]$_DFFE_PP_  (.D(net358),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][0] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][12]$_DFFE_PP_  (.D(net638),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][12] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][15] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][16]$_DFFE_PP_  (.D(net849),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][16] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][18]$_DFFE_PP_  (.D(net661),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][18] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][19] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][20] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][21]$_DFFE_PP_  (.D(net737),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][21] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][22]$_DFFE_PP_  (.D(net658),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][23]$_DFFE_PP_  (.D(net614),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][24]$_DFFE_PP_  (.D(net733),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][25]$_DFFE_PP_  (.D(net931),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][26]$_DFFE_PP_  (.D(net588),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][29]$_DFFE_PP_  (.D(net712),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][30]$_DFFE_PP_  (.D(net531),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][31]$_DFFE_PP_  (.D(net514),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][7]$_DFFE_PP_  (.D(net272),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][0]$_DFFE_PP_  (.D(net358),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][0] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][12]$_DFFE_PP_  (.D(net648),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][12] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][15] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][16]$_DFFE_PP_  (.D(net849),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][16] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][17]$_DFFE_PP_  (.D(net934),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][18]$_DFFE_PP_  (.D(net661),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][19] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][20] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][22]$_DFFE_PP_  (.D(net658),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][23]$_DFFE_PP_  (.D(net614),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][24]$_DFFE_PP_  (.D(net733),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][25]$_DFFE_PP_  (.D(net931),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][26]$_DFFE_PP_  (.D(net588),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][29]$_DFFE_PP_  (.D(net734),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][30]$_DFFE_PP_  (.D(net475),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][31]$_DFFE_PP_  (.D(net688),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][7]$_DFFE_PP_  (.D(net272),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][0]$_DFFE_PP_  (.D(net308),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][12]$_DFFE_PP_  (.D(net639),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][12] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][16]$_DFFE_PP_  (.D(net933),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][17]$_DFFE_PP_  (.D(net934),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][20] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][22]$_DFFE_PP_  (.D(net649),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][23]$_DFFE_PP_  (.D(net614),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][23] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][24]$_DFFE_PP_  (.D(net733),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][26]$_DFFE_PP_  (.D(net588),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][28]$_DFFE_PP_  (.D(net635),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][29]$_DFFE_PP_  (.D(net712),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][30]$_DFFE_PP_  (.D(net475),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][31]$_DFFE_PP_  (.D(net688),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][7]$_DFFE_PP_  (.D(net272),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][0]$_DFFE_PP_  (.D(net309),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][12]$_DFFE_PP_  (.D(net648),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][12] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][16]$_DFFE_PP_  (.D(net933),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][17]$_DFFE_PP_  (.D(net934),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][18]$_DFFE_PP_  (.D(net736),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][19] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][20] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][22]$_DFFE_PP_  (.D(net649),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][23]$_DFFE_PP_  (.D(net614),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][23] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][24]$_DFFE_PP_  (.D(net733),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][25]$_DFFE_PP_  (.D(net931),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][28]$_DFFE_PP_  (.D(net635),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][29]$_DFFE_PP_  (.D(net712),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][30]$_DFFE_PP_  (.D(net475),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][31]$_DFFE_PP_  (.D(net688),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][7]$_DFFE_PP_  (.D(net272),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][0]$_DFFE_PP_  (.D(net358),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][0] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][12]$_DFFE_PP_  (.D(net639),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][15] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][16]$_DFFE_PP_  (.D(net933),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][18] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][19] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][20]$_DFFE_PP_  (.D(net850),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][21]$_DFFE_PP_  (.D(net737),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][22]$_DFFE_PP_  (.D(net658),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][23]$_DFFE_PP_  (.D(net906),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][24]$_DFFE_PP_  (.D(net735),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][24] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][25]$_DFFE_PP_  (.D(net931),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][26]$_DFFE_PP_  (.D(net608),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][29]$_DFFE_PP_  (.D(net712),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][2] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][30]$_DFFE_PP_  (.D(net474),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][31]$_DFFE_PP_  (.D(net687),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][7]$_DFFE_PP_  (.D(net272),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][9] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][0]$_DFFE_PP_  (.D(net358),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][0] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][11] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][12]$_DFFE_PP_  (.D(net639),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][12] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][16]$_DFFE_PP_  (.D(net848),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][18]$_DFFE_PP_  (.D(net661),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][19] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][20]$_DFFE_PP_  (.D(net850),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][21]$_DFFE_PP_  (.D(net737),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][22]$_DFFE_PP_  (.D(net649),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][23]$_DFFE_PP_  (.D(net906),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][24]$_DFFE_PP_  (.D(net733),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][25]$_DFFE_PP_  (.D(net931),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][26]$_DFFE_PP_  (.D(net608),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][28]$_DFFE_PP_  (.D(net634),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][29]$_DFFE_PP_  (.D(net712),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][2] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][31]$_DFFE_PP_  (.D(net687),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][6]$_DFFE_PP_  (.D(net936),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][7]$_DFFE_PP_  (.D(net272),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][8] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][9] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][0]$_DFFE_PP_  (.D(net358),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][0] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][12]$_DFFE_PP_  (.D(net639),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][16]$_DFFE_PP_  (.D(net848),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][17] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][18]$_DFFE_PP_  (.D(net662),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][18] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][19] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][20]$_DFFE_PP_  (.D(net850),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][21]$_DFFE_PP_  (.D(net737),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][22]$_DFFE_PP_  (.D(net658),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][22] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][23]$_DFFE_PP_  (.D(net906),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][24]$_DFFE_PP_  (.D(net678),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][24] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][25]$_DFFE_PP_  (.D(net931),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][26]$_DFFE_PP_  (.D(net587),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][28]$_DFFE_PP_  (.D(net634),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][29]$_DFFE_PP_  (.D(net712),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][31]$_DFFE_PP_  (.D(net687),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][7]$_DFFE_PP_  (.D(net272),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][9] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][0]$_DFFE_PP_  (.D(net358),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][0] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][10] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][11] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][12]$_DFFE_PP_  (.D(net639),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][12] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][16]$_DFFE_PP_  (.D(net849),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][17] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][18]$_DFFE_PP_  (.D(net662),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][20] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][21]$_DFFE_PP_  (.D(net737),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][22]$_DFFE_PP_  (.D(net658),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][23]$_DFFE_PP_  (.D(net906),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][24]$_DFFE_PP_  (.D(net678),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][25]$_DFFE_PP_  (.D(net931),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][26]$_DFFE_PP_  (.D(net587),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][28]$_DFFE_PP_  (.D(net634),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][29]$_DFFE_PP_  (.D(net712),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][2] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][30]$_DFFE_PP_  (.D(net474),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][31]$_DFFE_PP_  (.D(net687),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][7]$_DFFE_PP_  (.D(net272),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][9] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][0]$_DFFE_PP_  (.D(net309),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][11] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][12]$_DFFE_PP_  (.D(net638),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][13] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][15] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][16]$_DFFE_PP_  (.D(net849),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][17] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][18]$_DFFE_PP_  (.D(net661),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][18] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][1] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][21]$_DFFE_PP_  (.D(net742),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][22]$_DFFE_PP_  (.D(net649),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][23]$_DFFE_PP_  (.D(net614),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][24]$_DFFE_PP_  (.D(net733),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][25]$_DFFE_PP_  (.D(net931),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][26]$_DFFE_PP_  (.D(net608),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][28]$_DFFE_PP_  (.D(net635),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][29]$_DFFE_PP_  (.D(net734),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][29] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][30]$_DFFE_PP_  (.D(net474),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][31]$_DFFE_PP_  (.D(net688),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][6]$_DFFE_PP_  (.D(net936),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][7]$_DFFE_PP_  (.D(net272),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][9] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][10] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][12]$_DFFE_PP_  (.D(net648),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][15] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][16]$_DFFE_PP_  (.D(net933),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][18] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][19] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][20]$_DFFE_PP_  (.D(net850),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][21]$_DFFE_PP_  (.D(net737),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][22]$_DFFE_PP_  (.D(net650),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][23]$_DFFE_PP_  (.D(net906),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][24]$_DFFE_PP_  (.D(net733),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][25]$_DFFE_PP_  (.D(net931),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][26]$_DFFE_PP_  (.D(net587),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][29]$_DFFE_PP_  (.D(net712),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][2] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][30]$_DFFE_PP_  (.D(net474),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][31]$_DFFE_PP_  (.D(net687),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][4] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][6]$_DFFE_PP_  (.D(net936),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][7]$_DFFE_PP_  (.D(net272),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][9] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][0]$_DFFE_PP_  (.D(net308),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][10] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][12]$_DFFE_PP_  (.D(net648),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][15] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][16]$_DFFE_PP_  (.D(net848),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][16] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][18]$_DFFE_PP_  (.D(net662),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][19] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][1] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][20]$_DFFE_PP_  (.D(net850),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][21]$_DFFE_PP_  (.D(net737),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][22]$_DFFE_PP_  (.D(net650),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][23]$_DFFE_PP_  (.D(net906),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][24]$_DFFE_PP_  (.D(net733),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][25]$_DFFE_PP_  (.D(net931),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][26]$_DFFE_PP_  (.D(net587),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][28]$_DFFE_PP_  (.D(net634),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][29]$_DFFE_PP_  (.D(net712),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][2] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][31]$_DFFE_PP_  (.D(net687),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][31] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][3] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][4] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][6]$_DFFE_PP_  (.D(net936),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][6] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][7]$_DFFE_PP_  (.D(net272),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][0]$_DFFE_PP_  (.D(net309),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][12]$_DFFE_PP_  (.D(net648),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][13] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][15] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][16]$_DFFE_PP_  (.D(net848),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][17]$_DFFE_PP_  (.D(net935),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][18]$_DFFE_PP_  (.D(net662),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][19] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][20]$_DFFE_PP_  (.D(net850),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][21]$_DFFE_PP_  (.D(net737),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][22]$_DFFE_PP_  (.D(net650),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][23]$_DFFE_PP_  (.D(net906),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][24]$_DFFE_PP_  (.D(net678),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][25]$_DFFE_PP_  (.D(net931),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][26]$_DFFE_PP_  (.D(net587),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][28]$_DFFE_PP_  (.D(net634),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][29]$_DFFE_PP_  (.D(net712),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][2] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][31]$_DFFE_PP_  (.D(net687),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][31] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][3] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][6]$_DFFE_PP_  (.D(net936),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][7]$_DFFE_PP_  (.D(net272),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][9] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][0]$_DFFE_PP_  (.D(net309),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][12]$_DFFE_PP_  (.D(net648),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][15] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][16]$_DFFE_PP_  (.D(net933),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][17] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][18]$_DFFE_PP_  (.D(net662),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][19] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][20]$_DFFE_PP_  (.D(net850),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][21]$_DFFE_PP_  (.D(net737),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][22]$_DFFE_PP_  (.D(net650),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][23]$_DFFE_PP_  (.D(net906),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][23] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][24]$_DFFE_PP_  (.D(net678),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][24] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][25]$_DFFE_PP_  (.D(net931),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][28]$_DFFE_PP_  (.D(net637),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][29]$_DFFE_PP_  (.D(net712),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][2] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][31]$_DFFE_PP_  (.D(net687),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][31] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][3] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][6]$_DFFE_PP_  (.D(net936),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][7]$_DFFE_PP_  (.D(net272),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][0]$_DFFE_PP_  (.D(net309),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][10] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][11] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][12]$_DFFE_PP_  (.D(net638),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][12] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][13] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][16]$_DFFE_PP_  (.D(net933),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][17]$_DFFE_PP_  (.D(net935),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][18]$_DFFE_PP_  (.D(net661),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][19] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][20]$_DFFE_PP_  (.D(net850),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][21]$_DFFE_PP_  (.D(net737),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][22] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][23]$_DFFE_PP_  (.D(net710),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][23] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][24]$_DFFE_PP_  (.D(net733),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][24] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][26]$_DFFE_PP_  (.D(net587),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][29]$_DFFE_PP_  (.D(net712),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][2] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][30]$_DFFE_PP_  (.D(net531),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][31]$_DFFE_PP_  (.D(net526),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][3] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][6]$_DFFE_PP_  (.D(net936),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][7]$_DFFE_PP_  (.D(net272),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][10] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][12]$_DFFE_PP_  (.D(net648),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][12] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][13] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][16]$_DFFE_PP_  (.D(net640),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][17]$_DFFE_PP_  (.D(net935),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][18]$_DFFE_PP_  (.D(net736),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][19] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][20]$_DFFE_PP_  (.D(net850),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][21]$_DFFE_PP_  (.D(net737),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][22]$_DFFE_PP_  (.D(net650),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][23]$_DFFE_PP_  (.D(net710),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][24]$_DFFE_PP_  (.D(net735),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][26]$_DFFE_PP_  (.D(net587),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][28]$_DFFE_PP_  (.D(net637),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][28] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][29]$_DFFE_PP_  (.D(net712),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][30]$_DFFE_PP_  (.D(net531),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][31]$_DFFE_PP_  (.D(net526),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][6]$_DFFE_PP_  (.D(net936),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][6] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][7]$_DFFE_PP_  (.D(net272),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][7] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][9] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][0]$_DFFE_PP_  (.D(net308),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][15] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][16]$_DFFE_PP_  (.D(net933),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][17]$_DFFE_PP_  (.D(net934),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][18]$_DFFE_PP_  (.D(net662),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][18] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][19] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][20]$_DFFE_PP_  (.D(net850),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][21]$_DFFE_PP_  (.D(net737),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][23]$_DFFE_PP_  (.D(net710),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][24]$_DFFE_PP_  (.D(net735),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][26]$_DFFE_PP_  (.D(net587),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][27] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][28]$_DFFE_PP_  (.D(net637),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][29]$_DFFE_PP_  (.D(net734),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][30]$_DFFE_PP_  (.D(net531),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][31]$_DFFE_PP_  (.D(net525),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][3] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][6]$_DFFE_PP_  (.D(net936),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][7]$_DFFE_PP_  (.D(net272),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][0]$_DFFE_PP_  (.D(net308),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][16]$_DFFE_PP_  (.D(net933),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][17]$_DFFE_PP_  (.D(net935),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][17] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][18]$_DFFE_PP_  (.D(net662),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][19] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][20]$_DFFE_PP_  (.D(net850),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][21]$_DFFE_PP_  (.D(net742),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][23]$_DFFE_PP_  (.D(net710),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][24]$_DFFE_PP_  (.D(net735),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][26]$_DFFE_PP_  (.D(net608),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][27] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][28]$_DFFE_PP_  (.D(net637),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][29]$_DFFE_PP_  (.D(net712),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][31]$_DFFE_PP_  (.D(net525),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][5] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][6]$_DFFE_PP_  (.D(net936),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][7]$_DFFE_PP_  (.D(net272),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][0]$_DFFE_PP_  (.D(net308),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][10] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][12]$_DFFE_PP_  (.D(net639),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][16]$_DFFE_PP_  (.D(net933),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][17]$_DFFE_PP_  (.D(net934),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][18] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][19] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][20]$_DFFE_PP_  (.D(net850),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][21]$_DFFE_PP_  (.D(net737),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][22] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][23]$_DFFE_PP_  (.D(net710),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][24]$_DFFE_PP_  (.D(net735),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][25] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][26]$_DFFE_PP_  (.D(net608),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][26] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][28]$_DFFE_PP_  (.D(net637),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][28] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][29]$_DFFE_PP_  (.D(net734),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][2] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][30]$_DFFE_PP_  (.D(net531),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][31]$_DFFE_PP_  (.D(net514),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][6]$_DFFE_PP_  (.D(net936),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][7]$_DFFE_PP_  (.D(net272),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][9] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][0]$_DFFE_PP_  (.D(net358),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][0] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][12]$_DFFE_PP_  (.D(net639),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][13] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][14] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][16]$_DFFE_PP_  (.D(net933),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][17]$_DFFE_PP_  (.D(net934),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][17] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][18] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][19] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][20]$_DFFE_PP_  (.D(net850),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][21]$_DFFE_PP_  (.D(net742),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][22] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][23]$_DFFE_PP_  (.D(net710),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][24]$_DFFE_PP_  (.D(net735),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][28] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][29]$_DFFE_PP_  (.D(net734),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][30]$_DFFE_PP_  (.D(net531),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][31]$_DFFE_PP_  (.D(net514),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][7]$_DFFE_PP_  (.D(net272),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][12]$_DFFE_PP_  (.D(net638),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][13] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][16]$_DFFE_PP_  (.D(net849),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][16] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][17] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][18]$_DFFE_PP_  (.D(net736),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][20] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][21]$_DFFE_PP_  (.D(net742),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][22]$_DFFE_PP_  (.D(net649),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][23]$_DFFE_PP_  (.D(net614),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][24]$_DFFE_PP_  (.D(net733),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][26]$_DFFE_PP_  (.D(net608),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][28]$_DFFE_PP_  (.D(net634),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][29]$_DFFE_PP_  (.D(net734),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][31]$_DFFE_PP_  (.D(net514),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][7]$_DFFE_PP_  (.D(net272),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][9] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][0]$_DFFE_PP_  (.D(net308),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][12]$_DFFE_PP_  (.D(net638),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][16]$_DFFE_PP_  (.D(net933),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][17]$_DFFE_PP_  (.D(net935),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][18] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][20]$_DFFE_PP_  (.D(net850),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][21]$_DFFE_PP_  (.D(net742),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][23]$_DFFE_PP_  (.D(net710),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][24]$_DFFE_PP_  (.D(net735),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][24] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][28]$_DFFE_PP_  (.D(net637),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][29]$_DFFE_PP_  (.D(net734),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][2] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][30]$_DFFE_PP_  (.D(net531),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][31]$_DFFE_PP_  (.D(net514),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][3] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][5] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][6]$_DFFE_PP_  (.D(net936),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][7]$_DFFE_PP_  (.D(net272),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][7] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][0]$_DFFE_PP_  (.D(net308),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][0] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][10] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][11] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][13] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][14] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][16]$_DFFE_PP_  (.D(net933),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][16] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][17]$_DFFE_PP_  (.D(net935),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][17] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][18]$_DFFE_PP_  (.D(net662),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][18] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][20]$_DFFE_PP_  (.D(net850),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][20] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][21]$_DFFE_PP_  (.D(net742),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][23]$_DFFE_PP_  (.D(net710),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][24]$_DFFE_PP_  (.D(net678),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][24] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][25] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][28]$_DFFE_PP_  (.D(net637),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][28] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][29]$_DFFE_PP_  (.D(net734),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][30]$_DFFE_PP_  (.D(\dp.result2[30] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][31]$_DFFE_PP_  (.D(net514),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][5] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][6]$_DFFE_PP_  (.D(net936),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][7]$_DFFE_PP_  (.D(net272),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][7] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][12]$_DFFE_PP_  (.D(net638),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][13] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][16]$_DFFE_PP_  (.D(net849),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][17] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][18]$_DFFE_PP_  (.D(net736),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][1] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][20] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][22]$_DFFE_PP_  (.D(net649),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][23]$_DFFE_PP_  (.D(net614),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][24]$_DFFE_PP_  (.D(net678),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][24] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][26]$_DFFE_PP_  (.D(net608),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][28]$_DFFE_PP_  (.D(net634),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][29]$_DFFE_PP_  (.D(net734),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][30]$_DFFE_PP_  (.D(net531),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][30] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][31]$_DFFE_PP_  (.D(net524),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][7]$_DFFE_PP_  (.D(net272),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][7] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][0]$_DFFE_PP_  (.D(net309),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][15] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][16]$_DFFE_PP_  (.D(net849),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][17]$_DFFE_PP_  (.D(net935),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][17] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][18]$_DFFE_PP_  (.D(net736),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][21]$_DFFE_PP_  (.D(net737),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][22]$_DFFE_PP_  (.D(net650),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][23]$_DFFE_PP_  (.D(net614),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][24]$_DFFE_PP_  (.D(net733),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][25]$_DFFE_PP_  (.D(net931),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][26]$_DFFE_PP_  (.D(net588),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][28]$_DFFE_PP_  (.D(net635),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][29]$_DFFE_PP_  (.D(net734),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][30]$_DFFE_PP_  (.D(net474),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][31]$_DFFE_PP_  (.D(net688),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][3] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][6]$_DFFE_PP_  (.D(net936),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][7]$_DFFE_PP_  (.D(net272),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][8] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][0]$_DFFE_PP_  (.D(net309),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][0] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][12]$_DFFE_PP_  (.D(net639),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][16]$_DFFE_PP_  (.D(net849),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][17] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][18] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][21]$_DFFE_PP_  (.D(net737),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][22]$_DFFE_PP_  (.D(net658),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][23]$_DFFE_PP_  (.D(net614),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][24]$_DFFE_PP_  (.D(net733),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][26]$_DFFE_PP_  (.D(net588),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][28]$_DFFE_PP_  (.D(net634),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][29]$_DFFE_PP_  (.D(net734),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][30]$_DFFE_PP_  (.D(net474),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][31]$_DFFE_PP_  (.D(net524),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][6]$_DFFE_PP_  (.D(net936),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][7]$_DFFE_PP_  (.D(net272),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][14] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][16]$_DFFE_PP_  (.D(net849),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][17] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][18] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][20] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][22]$_DFFE_PP_  (.D(net658),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][23]$_DFFE_PP_  (.D(net614),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][24]$_DFFE_PP_  (.D(net733),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][25]$_DFFE_PP_  (.D(net931),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][26]$_DFFE_PP_  (.D(net588),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][28]$_DFFE_PP_  (.D(net635),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][29]$_DFFE_PP_  (.D(net734),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][30]$_DFFE_PP_  (.D(net475),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][31]$_DFFE_PP_  (.D(net524),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][7]$_DFFE_PP_  (.D(net272),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][7] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][8] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][10] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][11] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][12] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][16]$_DFFE_PP_  (.D(net849),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][17] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][18]$_DFFE_PP_  (.D(net736),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][20] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][21]$_DFFE_PP_  (.D(net737),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][22]$_DFFE_PP_  (.D(net649),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][23]$_DFFE_PP_  (.D(net614),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][24]$_DFFE_PP_  (.D(net733),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][26]$_DFFE_PP_  (.D(net588),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][28]$_DFFE_PP_  (.D(net635),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][29]$_DFFE_PP_  (.D(net734),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][30]$_DFFE_PP_  (.D(net475),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][31]$_DFFE_PP_  (.D(net524),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][31] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][4] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][5] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][7]$_DFFE_PP_  (.D(net272),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][0]$_DFFE_PP_  (.D(net308),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][0] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][10] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][12]$_DFFE_PP_  (.D(net638),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][12] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][13] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][15] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][16]$_DFFE_PP_  (.D(net849),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][18]$_DFFE_PP_  (.D(net661),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][18] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][19] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][1] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][20] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][21]$_DFFE_PP_  (.D(net742),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][22]$_DFFE_PP_  (.D(net650),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][22] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][23]$_DFFE_PP_  (.D(net614),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][23] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][24]$_DFFE_PP_  (.D(net678),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][24] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][26]$_DFFE_PP_  (.D(\dp.result2[26] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][28]$_DFFE_PP_  (.D(net637),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][28] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][29]$_DFFE_PP_  (.D(net712),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][30]$_DFFE_PP_  (.D(net475),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][31]$_DFFE_PP_  (.D(net524),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][31] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][6]$_DFFE_PP_  (.D(net936),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][6] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][7]$_DFFE_PP_  (.D(net272),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][8] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][9] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][0]$_DFFE_PP_  (.D(net358),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][0] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][10] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][11] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][12]$_DFFE_PP_  (.D(net648),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][12] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][13] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][14] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][15] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][16]$_DFFE_PP_  (.D(net849),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][16] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][17]$_DFFE_PP_  (.D(\dp.result2[17] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][17] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][18]$_DFFE_PP_  (.D(net661),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][18] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][19]$_DFFE_PP_  (.D(\dp.result2[19] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][1] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][20] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][21] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][22]$_DFFE_PP_  (.D(net658),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][23]$_DFFE_PP_  (.D(net614),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][23] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][24]$_DFFE_PP_  (.D(net733),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][24] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][25]$_DFFE_PP_  (.D(net931),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][26]$_DFFE_PP_  (.D(net588),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][27]$_DFFE_PP_  (.D(\dp.result2[27] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][27] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][29]$_DFFE_PP_  (.D(net734),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][30]$_DFFE_PP_  (.D(net474),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][31]$_DFFE_PP_  (.D(net688),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][3] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][6] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][7]$_DFFE_PP_  (.D(net272),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][7] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][8] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][9] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1780 ();
 sky130_fd_sc_hd__buf_6 input1 (.A(instr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(instr[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(instr[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(instr[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_16 input5 (.A(instr[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_8 input6 (.A(instr[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_16 input7 (.A(instr[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_16 input8 (.A(instr[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(instr[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_16 input10 (.A(instr[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_16 input11 (.A(instr[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(instr[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_16 input13 (.A(instr[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_16 input14 (.A(instr[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_16 input15 (.A(instr[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_16 input16 (.A(instr[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_16 input17 (.A(instr[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(instr[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(instr[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(instr[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(instr[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(instr[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(instr[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_8 input24 (.A(instr[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(instr[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(instr[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(instr[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(instr[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(instr[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(instr[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(instr[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(instr[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(readdata[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(readdata[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(readdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(readdata[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(readdata[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(readdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(readdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(readdata[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(readdata[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(readdata[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(readdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(readdata[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(readdata[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(readdata[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(readdata[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(readdata[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(readdata[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(readdata[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(readdata[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(readdata[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(readdata[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(readdata[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(readdata[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(readdata[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(readdata[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(readdata[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(readdata[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(readdata[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(readdata[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(readdata[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(readdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(readdata[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_6 input65 (.A(reset),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(aluout[0]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(aluout[10]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(aluout[11]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(aluout[12]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(aluout[13]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(aluout[14]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(aluout[15]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(aluout[16]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(aluout[17]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(aluout[18]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(aluout[19]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(aluout[1]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(aluout[20]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(aluout[21]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(aluout[22]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(aluout[23]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(aluout[24]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(aluout[25]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(aluout[26]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(aluout[27]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(aluout[28]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(aluout[29]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(aluout[2]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(aluout[30]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(aluout[31]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(aluout[3]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(aluout[4]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(aluout[5]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(aluout[6]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(aluout[7]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(aluout[8]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(aluout[9]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(memread));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net99),
    .X(memwrite));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net100),
    .X(pc[0]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net101),
    .X(pc[10]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net102),
    .X(pc[11]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net103),
    .X(pc[12]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net104),
    .X(pc[13]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(pc[14]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(pc[15]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(pc[16]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net108),
    .X(pc[17]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(pc[18]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net110),
    .X(pc[19]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(pc[1]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(pc[20]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(pc[21]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(pc[22]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net115),
    .X(pc[23]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net116),
    .X(pc[24]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net117),
    .X(pc[25]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net118),
    .X(pc[26]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net119),
    .X(pc[27]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net120),
    .X(pc[28]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net121),
    .X(pc[29]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net122),
    .X(pc[2]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net123),
    .X(pc[30]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net124),
    .X(pc[31]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net125),
    .X(pc[3]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net126),
    .X(pc[4]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net127),
    .X(pc[5]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net128),
    .X(pc[6]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(pc[7]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(pc[8]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net131),
    .X(pc[9]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net132),
    .X(suspend));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net133),
    .X(writedata[0]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(writedata[10]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net135),
    .X(writedata[11]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net136),
    .X(writedata[12]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net137),
    .X(writedata[13]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(writedata[14]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net139),
    .X(writedata[15]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net140),
    .X(writedata[16]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net141),
    .X(writedata[17]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(writedata[18]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(writedata[19]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net413),
    .X(writedata[1]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net145),
    .X(writedata[20]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(writedata[21]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(writedata[22]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net148),
    .X(writedata[23]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net149),
    .X(writedata[24]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(writedata[25]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net151),
    .X(writedata[26]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(writedata[27]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net153),
    .X(writedata[28]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net154),
    .X(writedata[29]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(writedata[2]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net156),
    .X(writedata[30]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net157),
    .X(writedata[31]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(writedata[3]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net159),
    .X(writedata[4]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net160),
    .X(writedata[5]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(writedata[6]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net162),
    .X(writedata[7]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(writedata[8]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(writedata[9]));
 sky130_fd_sc_hd__buf_12 load_slew165 (.A(_1921_),
    .X(net165));
 sky130_fd_sc_hd__buf_16 load_slew166 (.A(_1921_),
    .X(net166));
 sky130_fd_sc_hd__buf_12 load_slew167 (.A(net707),
    .X(net167));
 sky130_fd_sc_hd__buf_16 load_slew168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_16 load_slew169 (.A(net246),
    .X(net169));
 sky130_fd_sc_hd__buf_16 load_slew170 (.A(_1890_),
    .X(net170));
 sky130_fd_sc_hd__buf_16 load_slew171 (.A(_1890_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 load_slew172 (.A(net175),
    .X(net172));
 sky130_fd_sc_hd__buf_6 load_slew173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_6 load_slew174 (.A(_1803_),
    .X(net174));
 sky130_fd_sc_hd__buf_6 load_slew175 (.A(_1803_),
    .X(net175));
 sky130_fd_sc_hd__buf_8 max_cap176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_8 max_cap177 (.A(_1809_),
    .X(net177));
 sky130_fd_sc_hd__buf_8 load_slew178 (.A(_0132_),
    .X(net178));
 sky130_fd_sc_hd__buf_16 load_slew179 (.A(_0132_),
    .X(net179));
 sky130_fd_sc_hd__buf_16 load_slew180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_16 load_slew181 (.A(_0348_),
    .X(net181));
 sky130_fd_sc_hd__buf_12 wire182 (.A(_0337_),
    .X(net182));
 sky130_fd_sc_hd__buf_16 load_slew183 (.A(_0337_),
    .X(net183));
 sky130_fd_sc_hd__buf_12 wire184 (.A(_0290_),
    .X(net184));
 sky130_fd_sc_hd__buf_12 wire185 (.A(_0256_),
    .X(net185));
 sky130_fd_sc_hd__buf_16 load_slew186 (.A(_0256_),
    .X(net186));
 sky130_fd_sc_hd__buf_16 load_slew187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_16 load_slew188 (.A(_0232_),
    .X(net188));
 sky130_fd_sc_hd__buf_16 load_slew189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__buf_12 wire190 (.A(_0221_),
    .X(net190));
 sky130_fd_sc_hd__buf_16 load_slew191 (.A(_0221_),
    .X(net191));
 sky130_fd_sc_hd__buf_16 load_slew192 (.A(_0212_),
    .X(net192));
 sky130_fd_sc_hd__buf_8 load_slew193 (.A(_0209_),
    .X(net193));
 sky130_fd_sc_hd__buf_8 load_slew194 (.A(_0209_),
    .X(net194));
 sky130_fd_sc_hd__buf_16 load_slew195 (.A(_0202_),
    .X(net195));
 sky130_fd_sc_hd__buf_16 max_cap196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_16 load_slew197 (.A(_0202_),
    .X(net197));
 sky130_fd_sc_hd__buf_16 load_slew198 (.A(_0192_),
    .X(net198));
 sky130_fd_sc_hd__buf_16 load_slew199 (.A(_0192_),
    .X(net199));
 sky130_fd_sc_hd__buf_16 load_slew200 (.A(_0176_),
    .X(net200));
 sky130_fd_sc_hd__buf_12 wire201 (.A(_0176_),
    .X(net201));
 sky130_fd_sc_hd__buf_16 load_slew202 (.A(_0128_),
    .X(net202));
 sky130_fd_sc_hd__buf_12 load_slew203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_12 wire204 (.A(_0263_),
    .X(net204));
 sky130_fd_sc_hd__buf_16 load_slew205 (.A(_0224_),
    .X(net205));
 sky130_fd_sc_hd__buf_16 load_slew206 (.A(net208),
    .X(net206));
 sky130_fd_sc_hd__buf_16 load_slew207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_16 load_slew208 (.A(net9),
    .X(net208));
 sky130_fd_sc_hd__buf_16 load_slew209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_16 load_slew210 (.A(net7),
    .X(net210));
 sky130_fd_sc_hd__buf_16 load_slew211 (.A(net7),
    .X(net211));
 sky130_fd_sc_hd__buf_16 load_slew212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_16 load_slew213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_16 load_slew214 (.A(net13),
    .X(net214));
 sky130_fd_sc_hd__buf_16 load_slew215 (.A(net13),
    .X(net215));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][0]$_DFFE_PP__216  (.LO(net216));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][10]$_DFFE_PP__217  (.LO(net217));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][11]$_DFFE_PP__218  (.LO(net218));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][12]$_DFFE_PP__219  (.LO(net219));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][13]$_DFFE_PP__220  (.LO(net220));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][14]$_DFFE_PP__221  (.LO(net221));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][15]$_DFFE_PP__222  (.LO(net222));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][18]$_DFFE_PP__223  (.LO(net223));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][19]$_DFFE_PP__224  (.LO(net224));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][1]$_DFFE_PP__225  (.LO(net225));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][20]$_DFFE_PP__226  (.LO(net226));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][21]$_DFFE_PP__227  (.LO(net227));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][22]$_DFFE_PP__228  (.LO(net228));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][23]$_DFFE_PP__229  (.LO(net229));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][24]$_DFFE_PP__230  (.LO(net230));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][25]$_DFFE_PP__231  (.LO(net231));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][26]$_DFFE_PP__232  (.LO(net232));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][27]$_DFFE_PP__233  (.LO(net233));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][28]$_DFFE_PP__234  (.LO(net234));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][29]$_DFFE_PP__235  (.LO(net235));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][2]$_DFFE_PP__236  (.LO(net236));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][30]$_DFFE_PP__237  (.LO(net237));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][31]$_DFFE_PP__238  (.LO(net238));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][3]$_DFFE_PP__239  (.LO(net239));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][4]$_DFFE_PP__240  (.LO(net240));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][5]$_DFFE_PP__241  (.LO(net241));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][6]$_DFFE_PP__242  (.LO(net242));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][7]$_DFFE_PP__243  (.LO(net243));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][8]$_DFFE_PP__244  (.LO(net244));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][9]$_DFFE_PP__245  (.LO(net245));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload1 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload3 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload4 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkinv_1 clkload10 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinv_1 clkload11 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_1 clkload12 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkinv_1 clkload13 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinv_2 clkload15 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__bufinv_16 clkload16 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload17 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_1 clkload18 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_1 clkload19 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkinv_4 clkload21 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload22 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload24 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__bufinv_16 clkload26 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__bufinv_16 clkload27 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__bufinv_16 clkload28 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_4 clkload29 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkinv_1 clkload30 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkinv_2 clkload31 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkinv_4 clkload32 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_1 clkload33 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload35 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_1 clkload36 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_2 clkload37 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload38 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_1 clkload39 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_1 clkload40 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkinv_1 clkload41 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinv_1 clkload43 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinv_2 clkload44 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__bufinv_16 clkload45 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload46 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload47 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload48 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinv_1 clkload49 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinv_1 clkload51 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkinv_2 clkload52 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_1 clkload53 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_1 clkload54 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload55 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_1 clkload56 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_2 clkload57 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinv_1 clkload58 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_2 clkload59 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__bufinv_16 clkload60 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_2 clkload61 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_1 clkload62 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkinv_2 clkload63 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkinv_2 clkload64 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload65 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload66 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_2 clkload67 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload68 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_2 clkload69 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_1 clkload70 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__bufinv_16 clkload71 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload72 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkinv_2 clkload73 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_1 clkload75 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload76 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_2 clkload77 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload78 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__bufinv_16 clkload80 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload81 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_6 clkload82 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__inv_6 clkload83 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload84 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkinv_1 clkload85 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkinv_2 clkload87 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_2 clkload88 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_1 clkload89 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload90 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload91 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_2 clkload92 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_1 clkload93 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__bufinv_16 clkload94 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkinv_1 clkload95 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__buf_8 rebuffer1 (.A(_1893_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net246),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net246),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net263),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net263),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(net246),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net246),
    .X(net252));
 sky130_fd_sc_hd__buf_4 rebuffer8 (.A(net252),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net253),
    .X(net254));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer10 (.A(net253),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_1893_),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_16 clone12 (.A(net260),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net169),
    .X(net258));
 sky130_fd_sc_hd__buf_2 rebuffer14 (.A(net258),
    .X(net259));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer15 (.A(net258),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_16 clone16 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(net246),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_16 clone18 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(_1893_),
    .X(net264));
 sky130_fd_sc_hd__o21a_2 clone20 (.A1(net408),
    .A2(_0138_),
    .B1(_1753_),
    .X(net265));
 sky130_fd_sc_hd__mux2i_2 clone21 (.A0(_1605_),
    .A1(net430),
    .S(net178),
    .Y(net266));
 sky130_fd_sc_hd__o21a_2 clone22 (.A1(net178),
    .A2(_3535_),
    .B1(net433),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer23 (.A(\dp.rf.rf[11][0] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(\dp.rf.rf[10][0] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 rebuffer25 (.A(_3518_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer26 (.A(net270),
    .X(net271));
 sky130_fd_sc_hd__buf_2 rebuffer30 (.A(_2697_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_16 clone31 (.A(net169),
    .X(net276));
 sky130_fd_sc_hd__buf_6 rebuffer35 (.A(net86),
    .X(net280));
 sky130_fd_sc_hd__buf_6 rebuffer39 (.A(net84),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(_1845_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 rebuffer56 (.A(net82),
    .X(net301));
 sky130_fd_sc_hd__a21oi_4 clone63 (.A1(_3130_),
    .A2(_3133_),
    .B1(_3134_),
    .Y(net308));
 sky130_fd_sc_hd__a21oi_4 clone64 (.A1(_3133_),
    .A2(_3130_),
    .B1(_3134_),
    .Y(net309));
 sky130_fd_sc_hd__a21oi_4 clone113 (.A1(_3130_),
    .A2(_3133_),
    .B1(_3134_),
    .Y(net358));
 sky130_fd_sc_hd__o21ai_4 clone162 (.A1(net410),
    .A2(_0138_),
    .B1(_1753_),
    .Y(net407));
 sky130_fd_sc_hd__buf_6 rebuffer163 (.A(net144),
    .X(net408));
 sky130_fd_sc_hd__buf_6 rebuffer164 (.A(net408),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer165 (.A(net409),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer166 (.A(net409),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer167 (.A(net409),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer168 (.A(net408),
    .X(net413));
 sky130_fd_sc_hd__buf_6 rebuffer175 (.A(_2680_),
    .X(net420));
 sky130_fd_sc_hd__buf_2 rebuffer176 (.A(_1702_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer177 (.A(net421),
    .X(net422));
 sky130_fd_sc_hd__buf_2 rebuffer178 (.A(net421),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer179 (.A(net423),
    .X(net424));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer180 (.A(net423),
    .X(net425));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer181 (.A(net421),
    .X(net426));
 sky130_fd_sc_hd__buf_2 rebuffer182 (.A(net426),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer183 (.A(_1618_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer184 (.A(_1618_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer185 (.A(net429),
    .X(net430));
 sky130_fd_sc_hd__mux2_4 clone186 (.A0(_3539_),
    .A1(net158),
    .S(net178),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer187 (.A(_1701_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer188 (.A(net432),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer189 (.A(\dp.rf.rf[21][2] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer190 (.A(_3510_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer191 (.A(\dp.rf.rf[20][2] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer192 (.A(_1619_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer193 (.A(net437),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer194 (.A(net437),
    .X(net439));
 sky130_fd_sc_hd__buf_6 rebuffer195 (.A(net437),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer196 (.A(net440),
    .X(net441));
 sky130_fd_sc_hd__buf_2 rebuffer197 (.A(net441),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer198 (.A(net440),
    .X(net443));
 sky130_fd_sc_hd__mux2_4 clone220 (.A0(_3539_),
    .A1(net158),
    .S(net178),
    .X(net465));
 sky130_fd_sc_hd__o21a_2 clone221 (.A1(net409),
    .A2(_0138_),
    .B1(_1753_),
    .X(net466));
 sky130_fd_sc_hd__o221ai_4 clone229 (.A1(_2781_),
    .A2(_3087_),
    .B1(_3232_),
    .B2(net530),
    .C1(_3234_),
    .Y(net474));
 sky130_fd_sc_hd__o221ai_4 clone230 (.A1(_2781_),
    .A2(_3087_),
    .B1(_3232_),
    .B2(net530),
    .C1(_3234_),
    .Y(net475));
 sky130_fd_sc_hd__buf_8 rebuffer252 (.A(_3279_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer253 (.A(net497),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer254 (.A(net497),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer255 (.A(net499),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer256 (.A(net497),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer257 (.A(net497),
    .X(net502));
 sky130_fd_sc_hd__buf_12 rebuffer285 (.A(_3233_),
    .X(net530));
 sky130_fd_sc_hd__o221ai_4 clone286 (.A1(_2781_),
    .A2(_3087_),
    .B1(_3232_),
    .B2(net530),
    .C1(_3234_),
    .Y(net531));
 sky130_fd_sc_hd__a21oi_4 clone342 (.A1(_3135_),
    .A2(_3058_),
    .B1(net607),
    .Y(net587));
 sky130_fd_sc_hd__a21oi_4 clone343 (.A1(_3135_),
    .A2(_3058_),
    .B1(net607),
    .Y(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer46 (.A(_2336_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer360 (.A(_3268_),
    .X(net605));
 sky130_fd_sc_hd__buf_6 rebuffer361 (.A(_0139_),
    .X(net606));
 sky130_fd_sc_hd__buf_12 rebuffer362 (.A(_3214_),
    .X(net607));
 sky130_fd_sc_hd__a21oi_4 clone363 (.A1(_3135_),
    .A2(_3058_),
    .B1(net607),
    .Y(net608));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer364 (.A(net79),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_2 rebuffer372 (.A(net83),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer380 (.A(net81),
    .X(net625));
 sky130_fd_sc_hd__o221ai_4 clone389 (.A1(_2781_),
    .A2(_3068_),
    .B1(_3075_),
    .B2(_2741_),
    .C1(_3222_),
    .Y(net634));
 sky130_fd_sc_hd__o221ai_4 clone390 (.A1(_2781_),
    .A2(_3068_),
    .B1(_3075_),
    .B2(_2741_),
    .C1(net636),
    .Y(net635));
 sky130_fd_sc_hd__buf_6 rebuffer391 (.A(_3222_),
    .X(net636));
 sky130_fd_sc_hd__o221ai_4 clone392 (.A1(_2781_),
    .A2(_3068_),
    .B1(_3075_),
    .B2(_2741_),
    .C1(_3222_),
    .Y(net637));
 sky130_fd_sc_hd__o221ai_4 clone393 (.A1(_2781_),
    .A2(_2940_),
    .B1(_2947_),
    .B2(_2741_),
    .C1(net492),
    .Y(net638));
 sky130_fd_sc_hd__o221ai_4 clone394 (.A1(_2781_),
    .A2(_2940_),
    .B1(_2947_),
    .B2(_2741_),
    .C1(net492),
    .Y(net639));
 sky130_fd_sc_hd__a211oi_4 clone395 (.A1(_3135_),
    .A2(_2976_),
    .B1(_3170_),
    .C1(_3171_),
    .Y(net640));
 sky130_fd_sc_hd__o221ai_4 clone403 (.A1(_2781_),
    .A2(_2940_),
    .B1(_2947_),
    .B2(_2741_),
    .C1(net492),
    .Y(net648));
 sky130_fd_sc_hd__o221ai_4 clone404 (.A1(_2781_),
    .A2(_3013_),
    .B1(_3020_),
    .B2(_2741_),
    .C1(net659),
    .Y(net649));
 sky130_fd_sc_hd__o221ai_4 clone405 (.A1(_2781_),
    .A2(_3013_),
    .B1(_3020_),
    .B2(_2741_),
    .C1(net659),
    .Y(net650));
 sky130_fd_sc_hd__o221ai_4 clone413 (.A1(_2781_),
    .A2(_3013_),
    .B1(_3020_),
    .B2(_2741_),
    .C1(net659),
    .Y(net658));
 sky130_fd_sc_hd__buf_12 rebuffer414 (.A(_3196_),
    .X(net659));
 sky130_fd_sc_hd__buf_6 rebuffer415 (.A(net659),
    .X(net660));
 sky130_fd_sc_hd__o221ai_4 clone416 (.A1(_2781_),
    .A2(_2985_),
    .B1(_2988_),
    .B2(_2741_),
    .C1(net663),
    .Y(net661));
 sky130_fd_sc_hd__o221ai_4 clone417 (.A1(_2781_),
    .A2(_2985_),
    .B1(_2988_),
    .B2(_2741_),
    .C1(net663),
    .Y(net662));
 sky130_fd_sc_hd__buf_12 rebuffer418 (.A(_3179_),
    .X(net663));
 sky130_fd_sc_hd__a2bb2oi_4 clone433 (.A1_N(net301),
    .A2_N(_3203_),
    .B1(_3206_),
    .B2(_3202_),
    .Y(net678));
 sky130_fd_sc_hd__a221oi_4 clone441 (.A1(_0128_),
    .A2(_3097_),
    .B1(net523),
    .B2(_3135_),
    .C1(net527),
    .Y(net686));
 sky130_fd_sc_hd__buf_6 rebuffer442 (.A(net686),
    .X(net687));
 sky130_fd_sc_hd__buf_6 rebuffer443 (.A(net686),
    .X(net688));
 sky130_fd_sc_hd__buf_6 rebuffer462 (.A(_1896_),
    .X(net707));
 sky130_fd_sc_hd__buf_2 rebuffer463 (.A(_1896_),
    .X(net708));
 sky130_fd_sc_hd__buf_6 rebuffer464 (.A(net708),
    .X(net709));
 sky130_fd_sc_hd__a21boi_4 clone465 (.A1(_3136_),
    .A2(net711),
    .B1_N(_3200_),
    .Y(net710));
 sky130_fd_sc_hd__buf_12 rebuffer466 (.A(_3199_),
    .X(net711));
 sky130_fd_sc_hd__o21ai_4 clone467 (.A1(_3225_),
    .A2(net420),
    .B1(_3228_),
    .Y(net712));
 sky130_fd_sc_hd__buf_16 wire1 (.A(\dp.result2[7] ),
    .X(net272));
 sky130_fd_sc_hd__buf_8 load_slew2 (.A(_3140_),
    .X(net273));
 sky130_fd_sc_hd__buf_16 load_slew3 (.A(net14),
    .X(net274));
 sky130_fd_sc_hd__buf_16 load_slew4 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_16 load_slew5 (.A(net14),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(_1844_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(_2268_),
    .X(net305));
 sky130_fd_sc_hd__buf_6 rebuffer62 (.A(net75),
    .X(net321));
 sky130_fd_sc_hd__buf_12 rebuffer226 (.A(_3151_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer227 (.A(net95),
    .X(net493));
 sky130_fd_sc_hd__buf_6 rebuffer242 (.A(net525),
    .X(net514));
 sky130_fd_sc_hd__buf_12 rebuffer243 (.A(_3487_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer244 (.A(net515),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer245 (.A(net515),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer246 (.A(net517),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer247 (.A(_3495_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer248 (.A(net519),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer249 (.A(_3495_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer250 (.A(net521),
    .X(net522));
 sky130_fd_sc_hd__buf_2 rebuffer251 (.A(_3103_),
    .X(net523));
 sky130_fd_sc_hd__buf_2 clone252 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_6 rebuffer258 (.A(\dp.result2[31] ),
    .X(net525));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer259 (.A(net525),
    .X(net526));
 sky130_fd_sc_hd__buf_12 rebuffer260 (.A(_3242_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer338 (.A(net94),
    .X(net613));
 sky130_fd_sc_hd__buf_12 rebuffer339 (.A(\dp.result2[23] ),
    .X(net614));
 sky130_fd_sc_hd__buf_12 rebuffer440 (.A(\dp.result2[24] ),
    .X(net733));
 sky130_fd_sc_hd__buf_12 rebuffer441 (.A(\dp.result2[29] ),
    .X(net734));
 sky130_fd_sc_hd__a2bb2oi_4 clone442 (.A1_N(net301),
    .A2_N(_3203_),
    .B1(_3206_),
    .B2(_3202_),
    .Y(net735));
 sky130_fd_sc_hd__o221ai_4 clone443 (.A1(_2781_),
    .A2(_2985_),
    .B1(_2988_),
    .B2(_2741_),
    .C1(net663),
    .Y(net736));
 sky130_fd_sc_hd__o221ai_4 clone444 (.A1(_2781_),
    .A2(_3008_),
    .B1(_3011_),
    .B2(_2741_),
    .C1(net814),
    .Y(net737));
 sky130_fd_sc_hd__o221ai_4 clone449 (.A1(_2781_),
    .A2(_3008_),
    .B1(_3011_),
    .B2(_2741_),
    .C1(net815),
    .Y(net742));
 sky130_fd_sc_hd__buf_12 rebuffer525 (.A(_3193_),
    .X(net814));
 sky130_fd_sc_hd__buf_4 rebuffer526 (.A(net814),
    .X(net815));
 sky130_fd_sc_hd__buf_6 rebuffer559 (.A(\dp.result2[16] ),
    .X(net848));
 sky130_fd_sc_hd__buf_6 rebuffer560 (.A(net848),
    .X(net849));
 sky130_fd_sc_hd__o221ai_4 clone561 (.A1(_2781_),
    .A2(_3000_),
    .B1(_3004_),
    .B2(_2741_),
    .C1(net851),
    .Y(net850));
 sky130_fd_sc_hd__buf_12 rebuffer562 (.A(_3190_),
    .X(net851));
 sky130_fd_sc_hd__buf_8 rebuffer563 (.A(_3463_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer564 (.A(net852),
    .X(net853));
 sky130_fd_sc_hd__buf_1 rebuffer565 (.A(net853),
    .X(net854));
 sky130_fd_sc_hd__buf_4 rebuffer566 (.A(net853),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer567 (.A(net855),
    .X(net856));
 sky130_fd_sc_hd__a21boi_4 clone617 (.A1(_3136_),
    .A2(net711),
    .B1_N(_3200_),
    .Y(net906));
 sky130_fd_sc_hd__o21a_2 clone642 (.A1(_3137_),
    .A2(net617),
    .B1(_3210_),
    .X(net931));
 sky130_fd_sc_hd__o21ai_2 clone643 (.A1(net178),
    .A2(_3535_),
    .B1(net432),
    .Y(net932));
 sky130_fd_sc_hd__buf_6 rebuffer644 (.A(net640),
    .X(net933));
 sky130_fd_sc_hd__o221ai_4 clone645 (.A1(_2781_),
    .A2(_2979_),
    .B1(_2983_),
    .B2(_2741_),
    .C1(_3176_),
    .Y(net934));
 sky130_fd_sc_hd__o221ai_4 clone646 (.A1(_2781_),
    .A2(_2979_),
    .B1(_2983_),
    .B2(_2741_),
    .C1(_3176_),
    .Y(net935));
 sky130_fd_sc_hd__a21boi_4 clone647 (.A1(_3249_),
    .A2(_3136_),
    .B1_N(_3250_),
    .Y(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\dp.result2[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\dp.result2[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_2833_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_752 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_801 ();
endmodule
