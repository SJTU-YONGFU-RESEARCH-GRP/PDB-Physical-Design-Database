module parameterized_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \clk_divider[0] ;
 wire \clk_divider[1] ;
 wire \clk_divider[2] ;
 wire \rx_shift[0] ;
 wire \rx_shift[1] ;
 wire \rx_shift[2] ;
 wire \rx_shift[3] ;
 wire \rx_shift[4] ;
 wire \rx_shift[5] ;
 wire \rx_shift[6] ;
 wire \rx_shift[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \tx_shift[0] ;
 wire \tx_shift[1] ;
 wire \tx_shift[2] ;
 wire \tx_shift[3] ;
 wire \tx_shift[4] ;
 wire \tx_shift[5] ;
 wire \tx_shift[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 INV_X2 _220_ (.A(net1),
    .ZN(_039_));
 BUF_X2 _221_ (.A(\state[0] ),
    .Z(_040_));
 BUF_X2 _222_ (.A(_195_),
    .Z(_041_));
 INV_X1 _223_ (.A(\clk_divider[2] ),
    .ZN(_042_));
 BUF_X2 _224_ (.A(_003_),
    .Z(_043_));
 INV_X1 _225_ (.A(net21),
    .ZN(_044_));
 NAND2_X1 _226_ (.A1(\bit_count[3] ),
    .A2(_199_),
    .ZN(_045_));
 CLKBUF_X2 _227_ (.A(\bit_count[2] ),
    .Z(_046_));
 OAI21_X1 _228_ (.A(_044_),
    .B1(_045_),
    .B2(_046_),
    .ZN(_047_));
 NAND4_X1 _229_ (.A1(_041_),
    .A2(_042_),
    .A3(_043_),
    .A4(_047_),
    .ZN(_048_));
 BUF_X4 _230_ (.A(\state[2] ),
    .Z(_049_));
 CLKBUF_X3 _231_ (.A(_049_),
    .Z(_050_));
 AOI22_X1 _232_ (.A1(net11),
    .A2(_040_),
    .B1(_048_),
    .B2(_050_),
    .ZN(_051_));
 NOR2_X1 _233_ (.A1(_039_),
    .A2(_051_),
    .ZN(_002_));
 INV_X1 _234_ (.A(_046_),
    .ZN(_052_));
 CLKBUF_X2 _235_ (.A(_201_),
    .Z(_053_));
 INV_X1 _236_ (.A(_053_),
    .ZN(_054_));
 NOR3_X4 _237_ (.A1(_052_),
    .A2(\bit_count[3] ),
    .A3(_054_),
    .ZN(_214_));
 CLKBUF_X3 _238_ (.A(\state[1] ),
    .Z(_055_));
 BUF_X2 _239_ (.A(net1),
    .Z(_056_));
 INV_X1 _240_ (.A(_040_),
    .ZN(_057_));
 OAI21_X1 _241_ (.A(_056_),
    .B1(_057_),
    .B2(net11),
    .ZN(_058_));
 OR2_X1 _242_ (.A1(_055_),
    .A2(_058_),
    .ZN(_001_));
 INV_X2 _243_ (.A(\state[2] ),
    .ZN(_059_));
 NAND2_X1 _244_ (.A1(_041_),
    .A2(_042_),
    .ZN(_060_));
 OR4_X1 _245_ (.A1(_046_),
    .A2(net21),
    .A3(_039_),
    .A4(_045_),
    .ZN(_061_));
 NOR3_X1 _246_ (.A1(_059_),
    .A2(_060_),
    .A3(_061_),
    .ZN(_000_));
 BUF_X1 _247_ (.A(\bit_count[0] ),
    .Z(_062_));
 NAND3_X1 _248_ (.A1(_046_),
    .A2(_062_),
    .A3(\bit_count[1] ),
    .ZN(_204_));
 INV_X1 _249_ (.A(_214_),
    .ZN(_207_));
 OR2_X1 _250_ (.A1(\bit_count[3] ),
    .A2(_204_),
    .ZN(_217_));
 NOR2_X2 _251_ (.A1(_049_),
    .A2(_040_),
    .ZN(_063_));
 INV_X1 _252_ (.A(net11),
    .ZN(_064_));
 AOI21_X2 _253_ (.A(_063_),
    .B1(_040_),
    .B2(_064_),
    .ZN(_065_));
 INV_X1 _254_ (.A(_041_),
    .ZN(_066_));
 NOR3_X2 _255_ (.A1(_066_),
    .A2(\clk_divider[2] ),
    .A3(_043_),
    .ZN(_067_));
 OAI21_X2 _256_ (.A(_065_),
    .B1(_067_),
    .B2(_059_),
    .ZN(_068_));
 OR4_X2 _257_ (.A1(_066_),
    .A2(\clk_divider[2] ),
    .A3(_059_),
    .A4(_210_),
    .ZN(_069_));
 NOR3_X4 _258_ (.A1(_043_),
    .A2(_214_),
    .A3(_069_),
    .ZN(_070_));
 OR4_X1 _259_ (.A1(_059_),
    .A2(_062_),
    .A3(_068_),
    .A4(_070_),
    .ZN(_071_));
 OAI21_X1 _260_ (.A(_062_),
    .B1(_068_),
    .B2(_070_),
    .ZN(_072_));
 AOI21_X1 _261_ (.A(_039_),
    .B1(_071_),
    .B2(_072_),
    .ZN(_004_));
 OAI21_X1 _262_ (.A(\bit_count[1] ),
    .B1(_068_),
    .B2(_070_),
    .ZN(_073_));
 BUF_X1 _263_ (.A(_200_),
    .Z(_074_));
 OR2_X1 _264_ (.A1(_049_),
    .A2(_040_),
    .ZN(_075_));
 OAI21_X1 _265_ (.A(_075_),
    .B1(_057_),
    .B2(net11),
    .ZN(_076_));
 OR3_X1 _266_ (.A1(_066_),
    .A2(\clk_divider[2] ),
    .A3(_043_),
    .ZN(_077_));
 AOI21_X2 _267_ (.A(_076_),
    .B1(_077_),
    .B2(_050_),
    .ZN(_078_));
 OR3_X1 _268_ (.A1(_043_),
    .A2(_214_),
    .A3(_069_),
    .ZN(_079_));
 NAND4_X1 _269_ (.A1(_050_),
    .A2(_074_),
    .A3(_078_),
    .A4(_079_),
    .ZN(_080_));
 AOI21_X1 _270_ (.A(_039_),
    .B1(_073_),
    .B2(_080_),
    .ZN(_005_));
 NOR2_X1 _271_ (.A1(_059_),
    .A2(_053_),
    .ZN(_081_));
 NOR3_X1 _272_ (.A1(_068_),
    .A2(_070_),
    .A3(_081_),
    .ZN(_082_));
 BUF_X2 _273_ (.A(_056_),
    .Z(_083_));
 NAND4_X1 _274_ (.A1(_052_),
    .A2(_083_),
    .A3(_050_),
    .A4(_053_),
    .ZN(_084_));
 OAI33_X1 _275_ (.A1(_052_),
    .A2(_039_),
    .A3(_082_),
    .B1(_084_),
    .B2(_068_),
    .B3(_070_),
    .ZN(_006_));
 OAI21_X1 _276_ (.A(\bit_count[3] ),
    .B1(_068_),
    .B2(_070_),
    .ZN(_085_));
 NAND4_X1 _277_ (.A1(_050_),
    .A2(_206_),
    .A3(_078_),
    .A4(_079_),
    .ZN(_086_));
 AOI21_X1 _278_ (.A(_039_),
    .B1(_085_),
    .B2(_086_),
    .ZN(_007_));
 MUX2_X1 _279_ (.A(_059_),
    .B(_075_),
    .S(\clk_divider[0] ),
    .Z(_087_));
 NOR2_X1 _280_ (.A1(_039_),
    .A2(_087_),
    .ZN(_008_));
 NAND3_X1 _281_ (.A1(_050_),
    .A2(_196_),
    .A3(_060_),
    .ZN(_088_));
 NAND2_X1 _282_ (.A1(\clk_divider[1] ),
    .A2(_063_),
    .ZN(_089_));
 AOI21_X1 _283_ (.A(_039_),
    .B1(_088_),
    .B2(_089_),
    .ZN(_009_));
 AOI21_X1 _284_ (.A(_063_),
    .B1(_050_),
    .B2(_066_),
    .ZN(_090_));
 NOR3_X1 _285_ (.A1(_042_),
    .A2(_039_),
    .A3(_090_),
    .ZN(_010_));
 BUF_X2 _286_ (.A(_083_),
    .Z(_091_));
 MUX2_X1 _287_ (.A(net12),
    .B(\rx_shift[0] ),
    .S(_055_),
    .Z(_092_));
 AND2_X1 _288_ (.A1(_091_),
    .A2(_092_),
    .ZN(_011_));
 MUX2_X1 _289_ (.A(net13),
    .B(\rx_shift[1] ),
    .S(_055_),
    .Z(_093_));
 AND2_X1 _290_ (.A1(_091_),
    .A2(_093_),
    .ZN(_012_));
 MUX2_X1 _291_ (.A(net14),
    .B(\rx_shift[2] ),
    .S(_055_),
    .Z(_094_));
 AND2_X1 _292_ (.A1(_091_),
    .A2(_094_),
    .ZN(_013_));
 MUX2_X1 _293_ (.A(net15),
    .B(\rx_shift[3] ),
    .S(_055_),
    .Z(_095_));
 AND2_X1 _294_ (.A1(_091_),
    .A2(_095_),
    .ZN(_014_));
 MUX2_X1 _295_ (.A(net16),
    .B(\rx_shift[4] ),
    .S(_055_),
    .Z(_096_));
 AND2_X1 _296_ (.A1(_091_),
    .A2(_096_),
    .ZN(_015_));
 MUX2_X1 _297_ (.A(net17),
    .B(\rx_shift[5] ),
    .S(_055_),
    .Z(_097_));
 AND2_X1 _298_ (.A1(_091_),
    .A2(_097_),
    .ZN(_016_));
 MUX2_X1 _299_ (.A(net18),
    .B(\rx_shift[6] ),
    .S(_055_),
    .Z(_098_));
 AND2_X1 _300_ (.A1(_091_),
    .A2(_098_),
    .ZN(_017_));
 MUX2_X1 _301_ (.A(net19),
    .B(\rx_shift[7] ),
    .S(_055_),
    .Z(_099_));
 AND2_X1 _302_ (.A1(_091_),
    .A2(_099_),
    .ZN(_018_));
 AND2_X1 _303_ (.A1(_056_),
    .A2(net2),
    .ZN(_100_));
 AND2_X1 _304_ (.A1(_083_),
    .A2(\rx_shift[0] ),
    .ZN(_101_));
 NOR4_X1 _305_ (.A1(_215_),
    .A2(_212_),
    .A3(_197_),
    .A4(_074_),
    .ZN(_102_));
 XNOR2_X2 _306_ (.A(_046_),
    .B(_053_),
    .ZN(_103_));
 AND2_X1 _307_ (.A1(_049_),
    .A2(_043_),
    .ZN(_104_));
 NAND4_X1 _308_ (.A1(_041_),
    .A2(_042_),
    .A3(_103_),
    .A4(_104_),
    .ZN(_105_));
 NOR2_X1 _309_ (.A1(_205_),
    .A2(_218_),
    .ZN(_106_));
 NAND3_X1 _310_ (.A1(_209_),
    .A2(_219_),
    .A3(_106_),
    .ZN(_107_));
 NOR2_X1 _311_ (.A1(_209_),
    .A2(_219_),
    .ZN(_108_));
 NAND3_X1 _312_ (.A1(_205_),
    .A2(_218_),
    .A3(_108_),
    .ZN(_109_));
 AOI21_X1 _313_ (.A(_105_),
    .B1(_107_),
    .B2(_109_),
    .ZN(_110_));
 NAND4_X1 _314_ (.A1(_209_),
    .A2(_206_),
    .A3(_102_),
    .A4(_110_),
    .ZN(_111_));
 MUX2_X1 _315_ (.A(_100_),
    .B(_101_),
    .S(_111_),
    .Z(_019_));
 AND2_X1 _316_ (.A1(_056_),
    .A2(\rx_shift[1] ),
    .ZN(_112_));
 NAND3_X1 _317_ (.A1(_041_),
    .A2(_042_),
    .A3(_104_),
    .ZN(_113_));
 NOR3_X2 _318_ (.A1(_206_),
    .A2(_103_),
    .A3(_113_),
    .ZN(_114_));
 INV_X1 _319_ (.A(_074_),
    .ZN(_115_));
 NOR2_X1 _320_ (.A1(_215_),
    .A2(_212_),
    .ZN(_116_));
 NAND4_X2 _321_ (.A1(_205_),
    .A2(_218_),
    .A3(_116_),
    .A4(_108_),
    .ZN(_117_));
 NOR3_X1 _322_ (.A1(_062_),
    .A2(_115_),
    .A3(_117_),
    .ZN(_118_));
 NAND2_X1 _323_ (.A1(_114_),
    .A2(_118_),
    .ZN(_119_));
 MUX2_X1 _324_ (.A(_100_),
    .B(_112_),
    .S(_119_),
    .Z(_020_));
 AND2_X1 _325_ (.A1(_056_),
    .A2(\rx_shift[2] ),
    .ZN(_120_));
 NOR3_X1 _326_ (.A1(_197_),
    .A2(_115_),
    .A3(_117_),
    .ZN(_121_));
 NAND2_X1 _327_ (.A1(_114_),
    .A2(_121_),
    .ZN(_122_));
 MUX2_X1 _328_ (.A(_100_),
    .B(_120_),
    .S(_122_),
    .Z(_021_));
 AND2_X1 _329_ (.A1(_056_),
    .A2(\rx_shift[3] ),
    .ZN(_123_));
 NOR3_X1 _330_ (.A1(_062_),
    .A2(_074_),
    .A3(_117_),
    .ZN(_124_));
 NAND2_X1 _331_ (.A1(_114_),
    .A2(_124_),
    .ZN(_125_));
 MUX2_X1 _332_ (.A(_100_),
    .B(_123_),
    .S(_125_),
    .Z(_022_));
 AND2_X1 _333_ (.A1(_056_),
    .A2(\rx_shift[4] ),
    .ZN(_126_));
 NOR3_X1 _334_ (.A1(_197_),
    .A2(_074_),
    .A3(_117_),
    .ZN(_127_));
 NAND2_X1 _335_ (.A1(_114_),
    .A2(_127_),
    .ZN(_128_));
 MUX2_X1 _336_ (.A(_100_),
    .B(_126_),
    .S(_128_),
    .Z(_023_));
 AND2_X1 _337_ (.A1(_056_),
    .A2(\rx_shift[5] ),
    .ZN(_129_));
 NOR2_X1 _338_ (.A1(_206_),
    .A2(_105_),
    .ZN(_130_));
 NAND2_X1 _339_ (.A1(_118_),
    .A2(_130_),
    .ZN(_131_));
 MUX2_X1 _340_ (.A(_100_),
    .B(_129_),
    .S(_131_),
    .Z(_024_));
 AND2_X1 _341_ (.A1(_056_),
    .A2(\rx_shift[6] ),
    .ZN(_132_));
 NAND2_X1 _342_ (.A1(_121_),
    .A2(_130_),
    .ZN(_133_));
 MUX2_X1 _343_ (.A(_100_),
    .B(_132_),
    .S(_133_),
    .Z(_025_));
 AND2_X1 _344_ (.A1(_056_),
    .A2(\rx_shift[7] ),
    .ZN(_134_));
 NAND2_X1 _345_ (.A1(_124_),
    .A2(_130_),
    .ZN(_135_));
 MUX2_X1 _346_ (.A(_100_),
    .B(_134_),
    .S(_135_),
    .Z(_026_));
 AND2_X1 _347_ (.A1(_091_),
    .A2(_055_),
    .ZN(_027_));
 OR3_X1 _348_ (.A1(_040_),
    .A2(\state[1] ),
    .A3(_113_),
    .ZN(_136_));
 NOR3_X1 _349_ (.A1(_050_),
    .A2(_040_),
    .A3(\state[1] ),
    .ZN(_137_));
 AOI21_X1 _350_ (.A(_137_),
    .B1(_060_),
    .B2(_050_),
    .ZN(_138_));
 OAI21_X1 _351_ (.A(_136_),
    .B1(_138_),
    .B2(_044_),
    .ZN(_139_));
 AND2_X1 _352_ (.A1(_091_),
    .A2(_139_),
    .ZN(_028_));
 AND2_X1 _353_ (.A1(_057_),
    .A2(net22),
    .ZN(_140_));
 OR2_X1 _354_ (.A1(_001_),
    .A2(_140_),
    .ZN(_029_));
 MUX2_X1 _355_ (.A(net10),
    .B(\tx_shift[6] ),
    .S(_050_),
    .Z(_141_));
 OAI221_X2 _356_ (.A(_065_),
    .B1(_069_),
    .B2(_044_),
    .C1(_059_),
    .C2(_067_),
    .ZN(_142_));
 BUF_X4 _357_ (.A(_142_),
    .Z(_143_));
 MUX2_X1 _358_ (.A(_141_),
    .B(net23),
    .S(_143_),
    .Z(_144_));
 AND2_X1 _359_ (.A1(_083_),
    .A2(_144_),
    .ZN(_030_));
 INV_X1 _360_ (.A(_058_),
    .ZN(_145_));
 INV_X1 _361_ (.A(net24),
    .ZN(_146_));
 OAI21_X1 _362_ (.A(_145_),
    .B1(_146_),
    .B2(_040_),
    .ZN(_031_));
 NAND2_X1 _363_ (.A1(\tx_shift[0] ),
    .A2(_143_),
    .ZN(_147_));
 NAND3_X1 _364_ (.A1(_059_),
    .A2(net3),
    .A3(_078_),
    .ZN(_148_));
 AOI21_X1 _365_ (.A(_039_),
    .B1(_147_),
    .B2(_148_),
    .ZN(_032_));
 MUX2_X1 _366_ (.A(net4),
    .B(\tx_shift[0] ),
    .S(_049_),
    .Z(_149_));
 MUX2_X1 _367_ (.A(_149_),
    .B(\tx_shift[1] ),
    .S(_143_),
    .Z(_150_));
 AND2_X1 _368_ (.A1(_083_),
    .A2(_150_),
    .ZN(_033_));
 MUX2_X1 _369_ (.A(net5),
    .B(\tx_shift[1] ),
    .S(_049_),
    .Z(_151_));
 MUX2_X1 _370_ (.A(_151_),
    .B(\tx_shift[2] ),
    .S(_143_),
    .Z(_152_));
 AND2_X1 _371_ (.A1(_083_),
    .A2(_152_),
    .ZN(_034_));
 MUX2_X1 _372_ (.A(net6),
    .B(\tx_shift[2] ),
    .S(_049_),
    .Z(_153_));
 MUX2_X1 _373_ (.A(_153_),
    .B(\tx_shift[3] ),
    .S(_143_),
    .Z(_154_));
 AND2_X1 _374_ (.A1(_083_),
    .A2(_154_),
    .ZN(_035_));
 MUX2_X1 _375_ (.A(net7),
    .B(\tx_shift[3] ),
    .S(_049_),
    .Z(_155_));
 MUX2_X1 _376_ (.A(_155_),
    .B(\tx_shift[4] ),
    .S(_143_),
    .Z(_156_));
 AND2_X1 _377_ (.A1(_083_),
    .A2(_156_),
    .ZN(_036_));
 MUX2_X1 _378_ (.A(net8),
    .B(\tx_shift[4] ),
    .S(_049_),
    .Z(_157_));
 MUX2_X1 _379_ (.A(_157_),
    .B(\tx_shift[5] ),
    .S(_143_),
    .Z(_158_));
 AND2_X1 _380_ (.A1(_083_),
    .A2(_158_),
    .ZN(_037_));
 MUX2_X1 _381_ (.A(net9),
    .B(\tx_shift[5] ),
    .S(_049_),
    .Z(_159_));
 MUX2_X1 _382_ (.A(_159_),
    .B(\tx_shift[6] ),
    .S(_143_),
    .Z(_160_));
 AND2_X1 _383_ (.A1(_083_),
    .A2(_160_),
    .ZN(_038_));
 HA_X1 _384_ (.A(\clk_divider[0] ),
    .B(\clk_divider[1] ),
    .CO(_195_),
    .S(_196_));
 HA_X1 _385_ (.A(_197_),
    .B(_198_),
    .CO(_199_),
    .S(_200_));
 HA_X1 _386_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_201_),
    .S(_202_));
 HA_X1 _387_ (.A(_203_),
    .B(_204_),
    .CO(_205_),
    .S(_206_));
 HA_X1 _388_ (.A(_203_),
    .B(_207_),
    .CO(_208_),
    .S(_209_));
 HA_X1 _389_ (.A(_203_),
    .B(_207_),
    .CO(_210_),
    .S(_211_));
 HA_X1 _390_ (.A(\bit_count[3] ),
    .B(_207_),
    .CO(_212_),
    .S(_213_));
 HA_X1 _391_ (.A(\bit_count[3] ),
    .B(_214_),
    .CO(_215_),
    .S(_216_));
 HA_X1 _392_ (.A(_203_),
    .B(_217_),
    .CO(_218_),
    .S(_219_));
 DFF_X2 \bit_count[0]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[0] ),
    .QN(_197_));
 DFF_X1 \bit_count[1]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[1] ),
    .QN(_198_));
 DFF_X1 \bit_count[2]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[2] ),
    .QN(_191_));
 DFF_X2 \bit_count[3]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[3] ),
    .QN(_203_));
 DFF_X1 \clk_divider[0]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\clk_divider[0] ),
    .QN(_190_));
 DFF_X1 \clk_divider[1]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\clk_divider[1] ),
    .QN(_189_));
 DFF_X2 \clk_divider[2]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\clk_divider[2] ),
    .QN(_188_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net12),
    .QN(_187_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_186_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net14),
    .QN(_185_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_184_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net16),
    .QN(_183_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net17),
    .QN(_182_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net18),
    .QN(_181_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net19),
    .QN(_180_));
 DFF_X1 \rx_shift[0]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[0] ),
    .QN(_179_));
 DFF_X1 \rx_shift[1]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[1] ),
    .QN(_178_));
 DFF_X1 \rx_shift[2]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[2] ),
    .QN(_177_));
 DFF_X1 \rx_shift[3]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[3] ),
    .QN(_176_));
 DFF_X1 \rx_shift[4]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[4] ),
    .QN(_175_));
 DFF_X1 \rx_shift[5]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift[5] ),
    .QN(_174_));
 DFF_X1 \rx_shift[6]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[6] ),
    .QN(_173_));
 DFF_X1 \rx_shift[7]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift[7] ),
    .QN(_172_));
 DFF_X1 \rx_valid$_SDFF_PN0_  (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net20),
    .QN(_171_));
 DFF_X1 \spi_clk$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net21),
    .QN(_003_));
 DFF_X1 \spi_cs_n$_SDFFE_PN1P_  (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net22),
    .QN(_170_));
 DFF_X1 \spi_mosi$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net23),
    .QN(_192_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[0] ),
    .QN(_193_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[1] ),
    .QN(_194_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[2] ),
    .QN(_169_));
 DFF_X1 \tx_ready$_SDFFE_PN1P_  (.D(_031_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net24),
    .QN(_168_));
 DFF_X1 \tx_shift[0]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[0] ),
    .QN(_167_));
 DFF_X1 \tx_shift[1]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[1] ),
    .QN(_166_));
 DFF_X1 \tx_shift[2]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[2] ),
    .QN(_165_));
 DFF_X1 \tx_shift[3]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[3] ),
    .QN(_164_));
 DFF_X1 \tx_shift[4]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[4] ),
    .QN(_163_));
 DFF_X1 \tx_shift[5]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift[5] ),
    .QN(_162_));
 DFF_X1 \tx_shift[6]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift[6] ),
    .QN(_161_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_89 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 input2 (.A(spi_miso),
    .Z(net2));
 BUF_X1 input3 (.A(tx_data[0]),
    .Z(net3));
 BUF_X1 input4 (.A(tx_data[1]),
    .Z(net4));
 BUF_X1 input5 (.A(tx_data[2]),
    .Z(net5));
 BUF_X1 input6 (.A(tx_data[3]),
    .Z(net6));
 BUF_X1 input7 (.A(tx_data[4]),
    .Z(net7));
 BUF_X1 input8 (.A(tx_data[5]),
    .Z(net8));
 BUF_X1 input9 (.A(tx_data[6]),
    .Z(net9));
 BUF_X1 input10 (.A(tx_data[7]),
    .Z(net10));
 CLKBUF_X2 input11 (.A(tx_valid),
    .Z(net11));
 BUF_X1 output12 (.A(net12),
    .Z(rx_data[0]));
 BUF_X1 output13 (.A(net13),
    .Z(rx_data[1]));
 BUF_X1 output14 (.A(net14),
    .Z(rx_data[2]));
 BUF_X1 output15 (.A(net15),
    .Z(rx_data[3]));
 BUF_X1 output16 (.A(net16),
    .Z(rx_data[4]));
 BUF_X1 output17 (.A(net17),
    .Z(rx_data[5]));
 BUF_X1 output18 (.A(net18),
    .Z(rx_data[6]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_data[7]));
 BUF_X1 output20 (.A(net20),
    .Z(rx_valid));
 BUF_X1 output21 (.A(net21),
    .Z(spi_clk));
 BUF_X1 output22 (.A(net22),
    .Z(spi_cs_n));
 BUF_X1 output23 (.A(net23),
    .Z(spi_mosi));
 BUF_X1 output24 (.A(net24),
    .Z(tx_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X4 clkload1 (.A(clknet_2_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_2_2__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_113 ();
 FILLCELL_X4 FILLER_0_120 ();
 FILLCELL_X2 FILLER_0_127 ();
 FILLCELL_X1 FILLER_0_129 ();
 FILLCELL_X4 FILLER_0_133 ();
 FILLCELL_X1 FILLER_0_137 ();
 FILLCELL_X8 FILLER_0_141 ();
 FILLCELL_X1 FILLER_0_149 ();
 FILLCELL_X8 FILLER_0_153 ();
 FILLCELL_X4 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_165 ();
 FILLCELL_X8 FILLER_0_174 ();
 FILLCELL_X2 FILLER_0_182 ();
 FILLCELL_X32 FILLER_0_190 ();
 FILLCELL_X32 FILLER_0_222 ();
 FILLCELL_X32 FILLER_0_254 ();
 FILLCELL_X32 FILLER_0_286 ();
 FILLCELL_X8 FILLER_0_318 ();
 FILLCELL_X4 FILLER_0_326 ();
 FILLCELL_X2 FILLER_0_330 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X1 FILLER_1_129 ();
 FILLCELL_X8 FILLER_1_137 ();
 FILLCELL_X4 FILLER_1_145 ();
 FILLCELL_X1 FILLER_1_149 ();
 FILLCELL_X16 FILLER_1_157 ();
 FILLCELL_X2 FILLER_1_173 ();
 FILLCELL_X1 FILLER_1_175 ();
 FILLCELL_X16 FILLER_1_179 ();
 FILLCELL_X2 FILLER_1_195 ();
 FILLCELL_X32 FILLER_1_214 ();
 FILLCELL_X32 FILLER_1_246 ();
 FILLCELL_X32 FILLER_1_278 ();
 FILLCELL_X16 FILLER_1_310 ();
 FILLCELL_X4 FILLER_1_326 ();
 FILLCELL_X2 FILLER_1_330 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X2 FILLER_2_136 ();
 FILLCELL_X8 FILLER_2_145 ();
 FILLCELL_X1 FILLER_2_153 ();
 FILLCELL_X2 FILLER_2_161 ();
 FILLCELL_X1 FILLER_2_163 ();
 FILLCELL_X16 FILLER_2_168 ();
 FILLCELL_X8 FILLER_2_184 ();
 FILLCELL_X32 FILLER_2_203 ();
 FILLCELL_X32 FILLER_2_235 ();
 FILLCELL_X32 FILLER_2_267 ();
 FILLCELL_X32 FILLER_2_299 ();
 FILLCELL_X1 FILLER_2_331 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X16 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_113 ();
 FILLCELL_X2 FILLER_3_117 ();
 FILLCELL_X1 FILLER_3_119 ();
 FILLCELL_X2 FILLER_3_141 ();
 FILLCELL_X1 FILLER_3_143 ();
 FILLCELL_X4 FILLER_3_148 ();
 FILLCELL_X1 FILLER_3_152 ();
 FILLCELL_X8 FILLER_3_177 ();
 FILLCELL_X2 FILLER_3_185 ();
 FILLCELL_X1 FILLER_3_187 ();
 FILLCELL_X2 FILLER_3_195 ();
 FILLCELL_X1 FILLER_3_197 ();
 FILLCELL_X32 FILLER_3_215 ();
 FILLCELL_X32 FILLER_3_247 ();
 FILLCELL_X32 FILLER_3_279 ();
 FILLCELL_X16 FILLER_3_311 ();
 FILLCELL_X4 FILLER_3_327 ();
 FILLCELL_X1 FILLER_3_331 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X16 FILLER_4_97 ();
 FILLCELL_X8 FILLER_4_113 ();
 FILLCELL_X4 FILLER_4_121 ();
 FILLCELL_X8 FILLER_4_132 ();
 FILLCELL_X8 FILLER_4_157 ();
 FILLCELL_X4 FILLER_4_165 ();
 FILLCELL_X2 FILLER_4_169 ();
 FILLCELL_X1 FILLER_4_171 ();
 FILLCELL_X4 FILLER_4_186 ();
 FILLCELL_X32 FILLER_4_201 ();
 FILLCELL_X32 FILLER_4_233 ();
 FILLCELL_X32 FILLER_4_265 ();
 FILLCELL_X32 FILLER_4_297 ();
 FILLCELL_X2 FILLER_4_329 ();
 FILLCELL_X1 FILLER_4_331 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_161 ();
 FILLCELL_X4 FILLER_5_169 ();
 FILLCELL_X1 FILLER_5_173 ();
 FILLCELL_X32 FILLER_5_178 ();
 FILLCELL_X32 FILLER_5_210 ();
 FILLCELL_X32 FILLER_5_242 ();
 FILLCELL_X32 FILLER_5_274 ();
 FILLCELL_X16 FILLER_5_306 ();
 FILLCELL_X8 FILLER_5_322 ();
 FILLCELL_X2 FILLER_5_330 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X16 FILLER_6_97 ();
 FILLCELL_X4 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_117 ();
 FILLCELL_X16 FILLER_6_149 ();
 FILLCELL_X4 FILLER_6_165 ();
 FILLCELL_X2 FILLER_6_169 ();
 FILLCELL_X32 FILLER_6_188 ();
 FILLCELL_X32 FILLER_6_220 ();
 FILLCELL_X32 FILLER_6_252 ();
 FILLCELL_X32 FILLER_6_284 ();
 FILLCELL_X16 FILLER_6_316 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X4 FILLER_7_129 ();
 FILLCELL_X1 FILLER_7_133 ();
 FILLCELL_X32 FILLER_7_138 ();
 FILLCELL_X32 FILLER_7_170 ();
 FILLCELL_X32 FILLER_7_202 ();
 FILLCELL_X32 FILLER_7_234 ();
 FILLCELL_X32 FILLER_7_266 ();
 FILLCELL_X32 FILLER_7_298 ();
 FILLCELL_X2 FILLER_7_330 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X16 FILLER_8_129 ();
 FILLCELL_X2 FILLER_8_145 ();
 FILLCELL_X1 FILLER_8_147 ();
 FILLCELL_X32 FILLER_8_151 ();
 FILLCELL_X8 FILLER_8_183 ();
 FILLCELL_X4 FILLER_8_191 ();
 FILLCELL_X2 FILLER_8_195 ();
 FILLCELL_X2 FILLER_8_202 ();
 FILLCELL_X1 FILLER_8_204 ();
 FILLCELL_X32 FILLER_8_222 ();
 FILLCELL_X32 FILLER_8_254 ();
 FILLCELL_X32 FILLER_8_286 ();
 FILLCELL_X8 FILLER_8_318 ();
 FILLCELL_X4 FILLER_8_326 ();
 FILLCELL_X2 FILLER_8_330 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X4 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_154 ();
 FILLCELL_X16 FILLER_9_186 ();
 FILLCELL_X1 FILLER_9_202 ();
 FILLCELL_X32 FILLER_9_220 ();
 FILLCELL_X32 FILLER_9_252 ();
 FILLCELL_X32 FILLER_9_284 ();
 FILLCELL_X16 FILLER_9_316 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X16 FILLER_10_129 ();
 FILLCELL_X2 FILLER_10_145 ();
 FILLCELL_X16 FILLER_10_151 ();
 FILLCELL_X2 FILLER_10_167 ();
 FILLCELL_X1 FILLER_10_169 ();
 FILLCELL_X1 FILLER_10_173 ();
 FILLCELL_X8 FILLER_10_188 ();
 FILLCELL_X4 FILLER_10_196 ();
 FILLCELL_X1 FILLER_10_207 ();
 FILLCELL_X2 FILLER_10_212 ();
 FILLCELL_X32 FILLER_10_224 ();
 FILLCELL_X32 FILLER_10_256 ();
 FILLCELL_X32 FILLER_10_288 ();
 FILLCELL_X8 FILLER_10_320 ();
 FILLCELL_X4 FILLER_10_328 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X16 FILLER_11_129 ();
 FILLCELL_X8 FILLER_11_145 ();
 FILLCELL_X4 FILLER_11_153 ();
 FILLCELL_X2 FILLER_11_157 ();
 FILLCELL_X16 FILLER_11_176 ();
 FILLCELL_X4 FILLER_11_192 ();
 FILLCELL_X2 FILLER_11_196 ();
 FILLCELL_X4 FILLER_11_205 ();
 FILLCELL_X32 FILLER_11_212 ();
 FILLCELL_X32 FILLER_11_244 ();
 FILLCELL_X32 FILLER_11_276 ();
 FILLCELL_X16 FILLER_11_308 ();
 FILLCELL_X8 FILLER_11_324 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X4 FILLER_12_161 ();
 FILLCELL_X2 FILLER_12_165 ();
 FILLCELL_X4 FILLER_12_170 ();
 FILLCELL_X4 FILLER_12_179 ();
 FILLCELL_X2 FILLER_12_183 ();
 FILLCELL_X2 FILLER_12_187 ();
 FILLCELL_X1 FILLER_12_197 ();
 FILLCELL_X16 FILLER_12_202 ();
 FILLCELL_X2 FILLER_12_218 ();
 FILLCELL_X1 FILLER_12_220 ();
 FILLCELL_X32 FILLER_12_231 ();
 FILLCELL_X32 FILLER_12_263 ();
 FILLCELL_X32 FILLER_12_295 ();
 FILLCELL_X4 FILLER_12_327 ();
 FILLCELL_X1 FILLER_12_331 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X16 FILLER_13_161 ();
 FILLCELL_X1 FILLER_13_177 ();
 FILLCELL_X2 FILLER_13_189 ();
 FILLCELL_X8 FILLER_13_207 ();
 FILLCELL_X2 FILLER_13_215 ();
 FILLCELL_X1 FILLER_13_217 ();
 FILLCELL_X16 FILLER_13_222 ();
 FILLCELL_X8 FILLER_13_238 ();
 FILLCELL_X4 FILLER_13_246 ();
 FILLCELL_X2 FILLER_13_250 ();
 FILLCELL_X32 FILLER_13_254 ();
 FILLCELL_X32 FILLER_13_286 ();
 FILLCELL_X8 FILLER_13_318 ();
 FILLCELL_X4 FILLER_13_326 ();
 FILLCELL_X2 FILLER_13_330 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X16 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_145 ();
 FILLCELL_X4 FILLER_14_153 ();
 FILLCELL_X4 FILLER_14_182 ();
 FILLCELL_X1 FILLER_14_193 ();
 FILLCELL_X4 FILLER_14_198 ();
 FILLCELL_X8 FILLER_14_205 ();
 FILLCELL_X2 FILLER_14_213 ();
 FILLCELL_X1 FILLER_14_215 ();
 FILLCELL_X32 FILLER_14_220 ();
 FILLCELL_X32 FILLER_14_252 ();
 FILLCELL_X32 FILLER_14_284 ();
 FILLCELL_X16 FILLER_14_316 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_169 ();
 FILLCELL_X1 FILLER_15_185 ();
 FILLCELL_X32 FILLER_15_220 ();
 FILLCELL_X32 FILLER_15_273 ();
 FILLCELL_X16 FILLER_15_305 ();
 FILLCELL_X8 FILLER_15_321 ();
 FILLCELL_X2 FILLER_15_329 ();
 FILLCELL_X1 FILLER_15_331 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X1 FILLER_16_169 ();
 FILLCELL_X1 FILLER_16_176 ();
 FILLCELL_X8 FILLER_16_195 ();
 FILLCELL_X4 FILLER_16_203 ();
 FILLCELL_X2 FILLER_16_207 ();
 FILLCELL_X1 FILLER_16_209 ();
 FILLCELL_X4 FILLER_16_224 ();
 FILLCELL_X2 FILLER_16_228 ();
 FILLCELL_X16 FILLER_16_234 ();
 FILLCELL_X4 FILLER_16_250 ();
 FILLCELL_X1 FILLER_16_254 ();
 FILLCELL_X4 FILLER_16_267 ();
 FILLCELL_X1 FILLER_16_271 ();
 FILLCELL_X1 FILLER_16_278 ();
 FILLCELL_X2 FILLER_16_298 ();
 FILLCELL_X16 FILLER_16_303 ();
 FILLCELL_X8 FILLER_16_319 ();
 FILLCELL_X4 FILLER_16_327 ();
 FILLCELL_X1 FILLER_16_331 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X4 FILLER_17_161 ();
 FILLCELL_X2 FILLER_17_165 ();
 FILLCELL_X1 FILLER_17_167 ();
 FILLCELL_X16 FILLER_17_181 ();
 FILLCELL_X8 FILLER_17_197 ();
 FILLCELL_X4 FILLER_17_205 ();
 FILLCELL_X1 FILLER_17_209 ();
 FILLCELL_X32 FILLER_17_214 ();
 FILLCELL_X8 FILLER_17_246 ();
 FILLCELL_X2 FILLER_17_254 ();
 FILLCELL_X32 FILLER_17_273 ();
 FILLCELL_X16 FILLER_17_305 ();
 FILLCELL_X8 FILLER_17_321 ();
 FILLCELL_X2 FILLER_17_329 ();
 FILLCELL_X1 FILLER_17_331 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X16 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_145 ();
 FILLCELL_X2 FILLER_18_153 ();
 FILLCELL_X1 FILLER_18_155 ();
 FILLCELL_X32 FILLER_18_177 ();
 FILLCELL_X8 FILLER_18_209 ();
 FILLCELL_X4 FILLER_18_217 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X4 FILLER_18_289 ();
 FILLCELL_X1 FILLER_18_293 ();
 FILLCELL_X32 FILLER_18_297 ();
 FILLCELL_X2 FILLER_18_329 ();
 FILLCELL_X1 FILLER_18_331 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X16 FILLER_19_129 ();
 FILLCELL_X4 FILLER_19_145 ();
 FILLCELL_X1 FILLER_19_149 ();
 FILLCELL_X16 FILLER_19_195 ();
 FILLCELL_X8 FILLER_19_211 ();
 FILLCELL_X4 FILLER_19_219 ();
 FILLCELL_X1 FILLER_19_223 ();
 FILLCELL_X32 FILLER_19_233 ();
 FILLCELL_X32 FILLER_19_265 ();
 FILLCELL_X32 FILLER_19_297 ();
 FILLCELL_X2 FILLER_19_329 ();
 FILLCELL_X1 FILLER_19_331 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X4 FILLER_20_129 ();
 FILLCELL_X2 FILLER_20_133 ();
 FILLCELL_X1 FILLER_20_135 ();
 FILLCELL_X8 FILLER_20_160 ();
 FILLCELL_X2 FILLER_20_168 ();
 FILLCELL_X1 FILLER_20_170 ();
 FILLCELL_X16 FILLER_20_173 ();
 FILLCELL_X4 FILLER_20_189 ();
 FILLCELL_X8 FILLER_20_205 ();
 FILLCELL_X2 FILLER_20_213 ();
 FILLCELL_X32 FILLER_20_222 ();
 FILLCELL_X32 FILLER_20_254 ();
 FILLCELL_X2 FILLER_20_286 ();
 FILLCELL_X1 FILLER_20_288 ();
 FILLCELL_X8 FILLER_20_293 ();
 FILLCELL_X4 FILLER_20_305 ();
 FILLCELL_X1 FILLER_20_309 ();
 FILLCELL_X4 FILLER_20_327 ();
 FILLCELL_X1 FILLER_20_331 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X16 FILLER_21_185 ();
 FILLCELL_X2 FILLER_21_201 ();
 FILLCELL_X16 FILLER_21_223 ();
 FILLCELL_X8 FILLER_21_239 ();
 FILLCELL_X1 FILLER_21_247 ();
 FILLCELL_X8 FILLER_21_273 ();
 FILLCELL_X1 FILLER_21_281 ();
 FILLCELL_X2 FILLER_21_289 ();
 FILLCELL_X1 FILLER_21_291 ();
 FILLCELL_X16 FILLER_21_309 ();
 FILLCELL_X1 FILLER_21_331 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X2 FILLER_22_21 ();
 FILLCELL_X32 FILLER_22_26 ();
 FILLCELL_X32 FILLER_22_58 ();
 FILLCELL_X32 FILLER_22_90 ();
 FILLCELL_X32 FILLER_22_122 ();
 FILLCELL_X4 FILLER_22_154 ();
 FILLCELL_X32 FILLER_22_162 ();
 FILLCELL_X4 FILLER_22_194 ();
 FILLCELL_X2 FILLER_22_198 ();
 FILLCELL_X1 FILLER_22_200 ();
 FILLCELL_X32 FILLER_22_211 ();
 FILLCELL_X2 FILLER_22_243 ();
 FILLCELL_X4 FILLER_22_255 ();
 FILLCELL_X1 FILLER_22_259 ();
 FILLCELL_X32 FILLER_22_284 ();
 FILLCELL_X16 FILLER_22_316 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X16 FILLER_23_129 ();
 FILLCELL_X2 FILLER_23_145 ();
 FILLCELL_X2 FILLER_23_157 ();
 FILLCELL_X8 FILLER_23_163 ();
 FILLCELL_X2 FILLER_23_171 ();
 FILLCELL_X2 FILLER_23_186 ();
 FILLCELL_X16 FILLER_23_193 ();
 FILLCELL_X4 FILLER_23_209 ();
 FILLCELL_X4 FILLER_23_221 ();
 FILLCELL_X1 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_231 ();
 FILLCELL_X32 FILLER_23_239 ();
 FILLCELL_X16 FILLER_23_271 ();
 FILLCELL_X8 FILLER_23_287 ();
 FILLCELL_X1 FILLER_23_295 ();
 FILLCELL_X8 FILLER_23_324 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X16 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_163 ();
 FILLCELL_X4 FILLER_24_179 ();
 FILLCELL_X2 FILLER_24_183 ();
 FILLCELL_X8 FILLER_24_189 ();
 FILLCELL_X4 FILLER_24_197 ();
 FILLCELL_X2 FILLER_24_211 ();
 FILLCELL_X1 FILLER_24_213 ();
 FILLCELL_X1 FILLER_24_231 ();
 FILLCELL_X16 FILLER_24_235 ();
 FILLCELL_X4 FILLER_24_251 ();
 FILLCELL_X2 FILLER_24_255 ();
 FILLCELL_X1 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_263 ();
 FILLCELL_X8 FILLER_24_295 ();
 FILLCELL_X16 FILLER_24_307 ();
 FILLCELL_X1 FILLER_24_323 ();
 FILLCELL_X4 FILLER_24_327 ();
 FILLCELL_X1 FILLER_24_331 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X4 FILLER_25_129 ();
 FILLCELL_X2 FILLER_25_133 ();
 FILLCELL_X1 FILLER_25_135 ();
 FILLCELL_X1 FILLER_25_155 ();
 FILLCELL_X4 FILLER_25_173 ();
 FILLCELL_X2 FILLER_25_180 ();
 FILLCELL_X2 FILLER_25_201 ();
 FILLCELL_X2 FILLER_25_207 ();
 FILLCELL_X1 FILLER_25_209 ();
 FILLCELL_X8 FILLER_25_237 ();
 FILLCELL_X1 FILLER_25_245 ();
 FILLCELL_X8 FILLER_25_249 ();
 FILLCELL_X2 FILLER_25_257 ();
 FILLCELL_X1 FILLER_25_259 ();
 FILLCELL_X2 FILLER_25_267 ();
 FILLCELL_X1 FILLER_25_269 ();
 FILLCELL_X16 FILLER_25_274 ();
 FILLCELL_X4 FILLER_25_290 ();
 FILLCELL_X2 FILLER_25_294 ();
 FILLCELL_X1 FILLER_25_296 ();
 FILLCELL_X8 FILLER_25_321 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X16 FILLER_26_129 ();
 FILLCELL_X4 FILLER_26_145 ();
 FILLCELL_X2 FILLER_26_149 ();
 FILLCELL_X16 FILLER_26_154 ();
 FILLCELL_X32 FILLER_26_183 ();
 FILLCELL_X4 FILLER_26_215 ();
 FILLCELL_X1 FILLER_26_219 ();
 FILLCELL_X8 FILLER_26_223 ();
 FILLCELL_X16 FILLER_26_243 ();
 FILLCELL_X2 FILLER_26_259 ();
 FILLCELL_X1 FILLER_26_261 ();
 FILLCELL_X32 FILLER_26_279 ();
 FILLCELL_X16 FILLER_26_311 ();
 FILLCELL_X4 FILLER_26_327 ();
 FILLCELL_X1 FILLER_26_331 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X4 FILLER_27_225 ();
 FILLCELL_X1 FILLER_27_229 ();
 FILLCELL_X1 FILLER_27_233 ();
 FILLCELL_X2 FILLER_27_237 ();
 FILLCELL_X1 FILLER_27_239 ();
 FILLCELL_X8 FILLER_27_249 ();
 FILLCELL_X4 FILLER_27_257 ();
 FILLCELL_X2 FILLER_27_268 ();
 FILLCELL_X1 FILLER_27_270 ();
 FILLCELL_X16 FILLER_27_275 ();
 FILLCELL_X8 FILLER_27_291 ();
 FILLCELL_X4 FILLER_27_299 ();
 FILLCELL_X1 FILLER_27_303 ();
 FILLCELL_X16 FILLER_27_308 ();
 FILLCELL_X8 FILLER_27_324 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X16 FILLER_28_161 ();
 FILLCELL_X8 FILLER_28_177 ();
 FILLCELL_X4 FILLER_28_185 ();
 FILLCELL_X2 FILLER_28_189 ();
 FILLCELL_X1 FILLER_28_191 ();
 FILLCELL_X32 FILLER_28_195 ();
 FILLCELL_X32 FILLER_28_227 ();
 FILLCELL_X4 FILLER_28_259 ();
 FILLCELL_X2 FILLER_28_263 ();
 FILLCELL_X1 FILLER_28_265 ();
 FILLCELL_X8 FILLER_28_283 ();
 FILLCELL_X4 FILLER_28_291 ();
 FILLCELL_X2 FILLER_28_295 ();
 FILLCELL_X1 FILLER_28_297 ();
 FILLCELL_X1 FILLER_28_322 ();
 FILLCELL_X4 FILLER_28_326 ();
 FILLCELL_X2 FILLER_28_330 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X2 FILLER_29_193 ();
 FILLCELL_X8 FILLER_29_199 ();
 FILLCELL_X4 FILLER_29_207 ();
 FILLCELL_X2 FILLER_29_211 ();
 FILLCELL_X32 FILLER_29_220 ();
 FILLCELL_X8 FILLER_29_252 ();
 FILLCELL_X2 FILLER_29_260 ();
 FILLCELL_X1 FILLER_29_262 ();
 FILLCELL_X2 FILLER_29_270 ();
 FILLCELL_X32 FILLER_29_276 ();
 FILLCELL_X16 FILLER_29_308 ();
 FILLCELL_X8 FILLER_29_324 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X4 FILLER_30_193 ();
 FILLCELL_X2 FILLER_30_214 ();
 FILLCELL_X4 FILLER_30_220 ();
 FILLCELL_X4 FILLER_30_235 ();
 FILLCELL_X1 FILLER_30_239 ();
 FILLCELL_X8 FILLER_30_247 ();
 FILLCELL_X1 FILLER_30_255 ();
 FILLCELL_X4 FILLER_30_260 ();
 FILLCELL_X8 FILLER_30_281 ();
 FILLCELL_X1 FILLER_30_289 ();
 FILLCELL_X16 FILLER_30_301 ();
 FILLCELL_X8 FILLER_30_317 ();
 FILLCELL_X4 FILLER_30_325 ();
 FILLCELL_X2 FILLER_30_329 ();
 FILLCELL_X1 FILLER_30_331 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X8 FILLER_31_193 ();
 FILLCELL_X2 FILLER_31_201 ();
 FILLCELL_X8 FILLER_31_207 ();
 FILLCELL_X2 FILLER_31_215 ();
 FILLCELL_X1 FILLER_31_217 ();
 FILLCELL_X8 FILLER_31_235 ();
 FILLCELL_X1 FILLER_31_243 ();
 FILLCELL_X32 FILLER_31_261 ();
 FILLCELL_X2 FILLER_31_293 ();
 FILLCELL_X1 FILLER_31_295 ();
 FILLCELL_X2 FILLER_31_313 ();
 FILLCELL_X8 FILLER_31_318 ();
 FILLCELL_X4 FILLER_31_326 ();
 FILLCELL_X2 FILLER_31_330 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X8 FILLER_32_321 ();
 FILLCELL_X2 FILLER_32_329 ();
 FILLCELL_X1 FILLER_32_331 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_193 ();
 FILLCELL_X4 FILLER_33_201 ();
 FILLCELL_X2 FILLER_33_205 ();
 FILLCELL_X8 FILLER_33_214 ();
 FILLCELL_X1 FILLER_33_222 ();
 FILLCELL_X16 FILLER_33_230 ();
 FILLCELL_X8 FILLER_33_246 ();
 FILLCELL_X32 FILLER_33_261 ();
 FILLCELL_X32 FILLER_33_293 ();
 FILLCELL_X4 FILLER_33_325 ();
 FILLCELL_X2 FILLER_33_329 ();
 FILLCELL_X1 FILLER_33_331 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X4 FILLER_34_214 ();
 FILLCELL_X16 FILLER_34_222 ();
 FILLCELL_X8 FILLER_34_238 ();
 FILLCELL_X4 FILLER_34_246 ();
 FILLCELL_X1 FILLER_34_250 ();
 FILLCELL_X32 FILLER_34_255 ();
 FILLCELL_X32 FILLER_34_287 ();
 FILLCELL_X8 FILLER_34_319 ();
 FILLCELL_X4 FILLER_34_327 ();
 FILLCELL_X1 FILLER_34_331 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X16 FILLER_35_193 ();
 FILLCELL_X4 FILLER_35_209 ();
 FILLCELL_X1 FILLER_35_213 ();
 FILLCELL_X16 FILLER_35_231 ();
 FILLCELL_X1 FILLER_35_247 ();
 FILLCELL_X32 FILLER_35_265 ();
 FILLCELL_X32 FILLER_35_297 ();
 FILLCELL_X2 FILLER_35_329 ();
 FILLCELL_X1 FILLER_35_331 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X8 FILLER_36_321 ();
 FILLCELL_X2 FILLER_36_329 ();
 FILLCELL_X1 FILLER_36_331 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X8 FILLER_37_321 ();
 FILLCELL_X2 FILLER_37_329 ();
 FILLCELL_X1 FILLER_37_331 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X8 FILLER_38_321 ();
 FILLCELL_X2 FILLER_38_329 ();
 FILLCELL_X1 FILLER_38_331 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X8 FILLER_39_321 ();
 FILLCELL_X2 FILLER_39_329 ();
 FILLCELL_X1 FILLER_39_331 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X8 FILLER_40_321 ();
 FILLCELL_X2 FILLER_40_329 ();
 FILLCELL_X1 FILLER_40_331 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X8 FILLER_41_321 ();
 FILLCELL_X2 FILLER_41_329 ();
 FILLCELL_X1 FILLER_41_331 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X8 FILLER_42_321 ();
 FILLCELL_X2 FILLER_42_329 ();
 FILLCELL_X1 FILLER_42_331 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X8 FILLER_43_321 ();
 FILLCELL_X2 FILLER_43_329 ();
 FILLCELL_X1 FILLER_43_331 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X16 FILLER_44_161 ();
 FILLCELL_X8 FILLER_44_177 ();
 FILLCELL_X2 FILLER_44_185 ();
 FILLCELL_X8 FILLER_44_190 ();
 FILLCELL_X1 FILLER_44_198 ();
 FILLCELL_X2 FILLER_44_202 ();
 FILLCELL_X8 FILLER_44_207 ();
 FILLCELL_X4 FILLER_44_215 ();
 FILLCELL_X32 FILLER_44_222 ();
 FILLCELL_X2 FILLER_44_254 ();
 FILLCELL_X1 FILLER_44_256 ();
 FILLCELL_X32 FILLER_44_260 ();
 FILLCELL_X32 FILLER_44_292 ();
 FILLCELL_X8 FILLER_44_324 ();
endmodule
