module uart (clk,
    m_axis_tready,
    m_axis_tvalid,
    rst,
    rx_busy,
    rx_frame_error,
    rx_overrun_error,
    rxd,
    s_axis_tready,
    s_axis_tvalid,
    tx_busy,
    txd,
    m_axis_tdata,
    prescale,
    s_axis_tdata);
 input clk;
 input m_axis_tready;
 output m_axis_tvalid;
 input rst;
 output rx_busy;
 output rx_frame_error;
 output rx_overrun_error;
 input rxd;
 output s_axis_tready;
 input s_axis_tvalid;
 output tx_busy;
 output txd;
 output [7:0] m_axis_tdata;
 input [15:0] prescale;
 input [7:0] s_axis_tdata;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire net41;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire \uart_rx_inst.bit_cnt[0] ;
 wire \uart_rx_inst.bit_cnt[1] ;
 wire \uart_rx_inst.bit_cnt[2] ;
 wire \uart_rx_inst.bit_cnt[3] ;
 wire \uart_rx_inst.data_reg[0] ;
 wire \uart_rx_inst.data_reg[1] ;
 wire \uart_rx_inst.data_reg[2] ;
 wire \uart_rx_inst.data_reg[3] ;
 wire \uart_rx_inst.data_reg[4] ;
 wire \uart_rx_inst.data_reg[5] ;
 wire \uart_rx_inst.data_reg[6] ;
 wire \uart_rx_inst.data_reg[7] ;
 wire \uart_rx_inst.prescale_reg[0] ;
 wire \uart_rx_inst.prescale_reg[10] ;
 wire \uart_rx_inst.prescale_reg[11] ;
 wire \uart_rx_inst.prescale_reg[12] ;
 wire \uart_rx_inst.prescale_reg[13] ;
 wire \uart_rx_inst.prescale_reg[14] ;
 wire \uart_rx_inst.prescale_reg[15] ;
 wire \uart_rx_inst.prescale_reg[16] ;
 wire \uart_rx_inst.prescale_reg[17] ;
 wire \uart_rx_inst.prescale_reg[18] ;
 wire \uart_rx_inst.prescale_reg[1] ;
 wire \uart_rx_inst.prescale_reg[2] ;
 wire \uart_rx_inst.prescale_reg[3] ;
 wire \uart_rx_inst.prescale_reg[4] ;
 wire \uart_rx_inst.prescale_reg[5] ;
 wire \uart_rx_inst.prescale_reg[6] ;
 wire \uart_rx_inst.prescale_reg[7] ;
 wire \uart_rx_inst.prescale_reg[8] ;
 wire \uart_rx_inst.prescale_reg[9] ;
 wire \uart_rx_inst.rxd_reg ;
 wire \uart_tx_inst.bit_cnt[0] ;
 wire \uart_tx_inst.bit_cnt[1] ;
 wire \uart_tx_inst.bit_cnt[2] ;
 wire \uart_tx_inst.bit_cnt[3] ;
 wire \uart_tx_inst.data_reg[0] ;
 wire \uart_tx_inst.data_reg[1] ;
 wire \uart_tx_inst.data_reg[2] ;
 wire \uart_tx_inst.data_reg[3] ;
 wire \uart_tx_inst.data_reg[4] ;
 wire \uart_tx_inst.data_reg[5] ;
 wire \uart_tx_inst.data_reg[6] ;
 wire \uart_tx_inst.data_reg[7] ;
 wire \uart_tx_inst.data_reg[8] ;
 wire \uart_tx_inst.prescale_reg[0] ;
 wire \uart_tx_inst.prescale_reg[10] ;
 wire \uart_tx_inst.prescale_reg[11] ;
 wire \uart_tx_inst.prescale_reg[12] ;
 wire \uart_tx_inst.prescale_reg[13] ;
 wire \uart_tx_inst.prescale_reg[14] ;
 wire \uart_tx_inst.prescale_reg[15] ;
 wire \uart_tx_inst.prescale_reg[16] ;
 wire \uart_tx_inst.prescale_reg[17] ;
 wire \uart_tx_inst.prescale_reg[18] ;
 wire \uart_tx_inst.prescale_reg[1] ;
 wire \uart_tx_inst.prescale_reg[2] ;
 wire \uart_tx_inst.prescale_reg[3] ;
 wire \uart_tx_inst.prescale_reg[4] ;
 wire \uart_tx_inst.prescale_reg[5] ;
 wire \uart_tx_inst.prescale_reg[6] ;
 wire \uart_tx_inst.prescale_reg[7] ;
 wire \uart_tx_inst.prescale_reg[8] ;
 wire \uart_tx_inst.prescale_reg[9] ;
 wire net2;
 wire net1;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net40;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;

 sky130_fd_sc_hd__buf_2 _431_ (.A(\uart_tx_inst.bit_cnt[0] ),
    .X(_081_));
 sky130_fd_sc_hd__nor4_4 _432_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .B(\uart_tx_inst.bit_cnt[3] ),
    .C(\uart_tx_inst.bit_cnt[1] ),
    .D(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__clkbuf_4 _433_ (.A(_082_),
    .X(_002_));
 sky130_fd_sc_hd__clkbuf_4 _434_ (.A(\uart_rx_inst.bit_cnt[3] ),
    .X(_083_));
 sky130_fd_sc_hd__buf_2 _435_ (.A(\uart_rx_inst.bit_cnt[2] ),
    .X(_084_));
 sky130_fd_sc_hd__nor2_1 _436_ (.A(\uart_rx_inst.bit_cnt[1] ),
    .B(_421_),
    .Y(_085_));
 sky130_fd_sc_hd__a21oi_1 _437_ (.A1(\uart_rx_inst.rxd_reg ),
    .A2(_421_),
    .B1(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__nor3_4 _438_ (.A(_083_),
    .B(_084_),
    .C(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__or4_4 _439_ (.A(\uart_rx_inst.prescale_reg[11] ),
    .B(\uart_rx_inst.prescale_reg[13] ),
    .C(\uart_rx_inst.prescale_reg[12] ),
    .D(\uart_rx_inst.prescale_reg[10] ),
    .X(_088_));
 sky130_fd_sc_hd__or3_4 _440_ (.A(\uart_rx_inst.prescale_reg[15] ),
    .B(\uart_rx_inst.prescale_reg[14] ),
    .C(_088_),
    .X(_089_));
 sky130_fd_sc_hd__or3_1 _441_ (.A(\uart_rx_inst.prescale_reg[17] ),
    .B(\uart_rx_inst.prescale_reg[18] ),
    .C(\uart_rx_inst.prescale_reg[16] ),
    .X(_090_));
 sky130_fd_sc_hd__nor3_2 _442_ (.A(\uart_rx_inst.prescale_reg[4] ),
    .B(\uart_rx_inst.prescale_reg[3] ),
    .C(\uart_rx_inst.prescale_reg[2] ),
    .Y(_091_));
 sky130_fd_sc_hd__nor3_1 _443_ (.A(\uart_rx_inst.prescale_reg[5] ),
    .B(\uart_rx_inst.prescale_reg[1] ),
    .C(\uart_rx_inst.prescale_reg[0] ),
    .Y(_092_));
 sky130_fd_sc_hd__nor4_2 _444_ (.A(\uart_rx_inst.prescale_reg[9] ),
    .B(\uart_rx_inst.prescale_reg[7] ),
    .C(\uart_rx_inst.prescale_reg[8] ),
    .D(\uart_rx_inst.prescale_reg[6] ),
    .Y(_093_));
 sky130_fd_sc_hd__nand3_2 _445_ (.A(_091_),
    .B(_092_),
    .C(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__or3_4 _446_ (.A(_090_),
    .B(_094_),
    .C(_089_),
    .X(_095_));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(_095_),
    .X(net41));
 sky130_fd_sc_hd__o21bai_2 _448_ (.A1(_423_),
    .A2(_425_),
    .B1_N(_084_),
    .Y(_097_));
 sky130_fd_sc_hd__and2_0 _449_ (.A(_083_),
    .B(_097_),
    .X(_098_));
 sky130_fd_sc_hd__or3_4 _450_ (.A(_095_),
    .B(_098_),
    .C(net14),
    .X(_099_));
 sky130_fd_sc_hd__nor2_8 _451_ (.A(_087_),
    .B(_099_),
    .Y(_001_));
 sky130_fd_sc_hd__clkbuf_4 _452_ (.A(net14),
    .X(_100_));
 sky130_fd_sc_hd__clkbuf_4 _453_ (.A(_100_),
    .X(_101_));
 sky130_fd_sc_hd__nand2b_1 _454_ (.A_N(net24),
    .B(_082_),
    .Y(_102_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(\uart_tx_inst.prescale_reg[5] ),
    .B(\uart_tx_inst.prescale_reg[4] ),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _456_ (.A(\uart_tx_inst.prescale_reg[1] ),
    .B(\uart_tx_inst.prescale_reg[0] ),
    .Y(_104_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(\uart_tx_inst.prescale_reg[3] ),
    .B(\uart_tx_inst.prescale_reg[2] ),
    .Y(_105_));
 sky130_fd_sc_hd__nor3_2 _458_ (.A(\uart_tx_inst.prescale_reg[8] ),
    .B(\uart_tx_inst.prescale_reg[7] ),
    .C(\uart_tx_inst.prescale_reg[6] ),
    .Y(_106_));
 sky130_fd_sc_hd__nand4_2 _459_ (.A(_103_),
    .B(_104_),
    .C(_105_),
    .D(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__nor4_2 _460_ (.A(\uart_tx_inst.prescale_reg[17] ),
    .B(\uart_tx_inst.prescale_reg[15] ),
    .C(\uart_tx_inst.prescale_reg[16] ),
    .D(\uart_tx_inst.prescale_reg[14] ),
    .Y(_108_));
 sky130_fd_sc_hd__nor3_1 _461_ (.A(\uart_tx_inst.prescale_reg[11] ),
    .B(\uart_tx_inst.prescale_reg[10] ),
    .C(\uart_tx_inst.prescale_reg[9] ),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _462_ (.A(\uart_tx_inst.prescale_reg[13] ),
    .B(\uart_tx_inst.prescale_reg[12] ),
    .Y(_110_));
 sky130_fd_sc_hd__nand4b_1 _463_ (.A_N(\uart_tx_inst.prescale_reg[18] ),
    .B(_108_),
    .C(_109_),
    .D(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__nor2_1 _464_ (.A(_107_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__buf_2 _465_ (.A(_112_),
    .X(_113_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(_102_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__nor4b_2 _467_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .B(\uart_tx_inst.bit_cnt[3] ),
    .C(\uart_tx_inst.bit_cnt[1] ),
    .D_N(_081_),
    .Y(_115_));
 sky130_fd_sc_hd__clkbuf_4 _468_ (.A(_115_),
    .X(_116_));
 sky130_fd_sc_hd__nor3_4 _469_ (.A(_101_),
    .B(_116_),
    .C(_114_),
    .Y(_000_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(\uart_tx_inst.data_reg[1] ),
    .A1(net16),
    .S(_002_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(\uart_tx_inst.data_reg[2] ),
    .A1(net17),
    .S(_002_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\uart_tx_inst.data_reg[3] ),
    .A1(net18),
    .S(_002_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(\uart_tx_inst.data_reg[4] ),
    .A1(net19),
    .S(_002_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(\uart_tx_inst.data_reg[5] ),
    .A1(net20),
    .S(_002_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(\uart_tx_inst.data_reg[6] ),
    .A1(net21),
    .S(_002_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(\uart_tx_inst.data_reg[7] ),
    .A1(net22),
    .S(_082_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(\uart_tx_inst.data_reg[8] ),
    .A1(net23),
    .S(_082_),
    .X(_010_));
 sky130_fd_sc_hd__inv_1 _478_ (.A(\uart_rx_inst.prescale_reg[0] ),
    .Y(_411_));
 sky130_fd_sc_hd__inv_1 _479_ (.A(net3),
    .Y(_415_));
 sky130_fd_sc_hd__inv_1 _480_ (.A(\uart_tx_inst.prescale_reg[0] ),
    .Y(_427_));
 sky130_fd_sc_hd__inv_1 _481_ (.A(\uart_rx_inst.bit_cnt[0] ),
    .Y(_419_));
 sky130_fd_sc_hd__inv_1 _482_ (.A(\uart_rx_inst.prescale_reg[1] ),
    .Y(_412_));
 sky130_fd_sc_hd__inv_1 _483_ (.A(net9),
    .Y(_416_));
 sky130_fd_sc_hd__inv_1 _484_ (.A(\uart_rx_inst.bit_cnt[1] ),
    .Y(_420_));
 sky130_fd_sc_hd__inv_1 _485_ (.A(\uart_tx_inst.prescale_reg[1] ),
    .Y(_428_));
 sky130_fd_sc_hd__clkbuf_4 _486_ (.A(_100_),
    .X(_117_));
 sky130_fd_sc_hd__clkbuf_4 _487_ (.A(\uart_rx_inst.rxd_reg ),
    .X(_118_));
 sky130_fd_sc_hd__nor3b_4 _488_ (.A(_083_),
    .B(_084_),
    .C_N(_421_),
    .Y(_119_));
 sky130_fd_sc_hd__a31o_2 _489_ (.A1(_118_),
    .A2(_083_),
    .A3(_097_),
    .B1(_119_),
    .X(_120_));
 sky130_fd_sc_hd__clkbuf_4 _490_ (.A(_120_),
    .X(_121_));
 sky130_fd_sc_hd__nor2_1 _491_ (.A(\uart_rx_inst.bit_cnt[0] ),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__nor2_1 _492_ (.A(_083_),
    .B(_084_),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _493_ (.A(_118_),
    .B(_421_),
    .Y(_124_));
 sky130_fd_sc_hd__o31ai_1 _494_ (.A1(\uart_rx_inst.bit_cnt[1] ),
    .A2(_421_),
    .A3(_425_),
    .B1(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a21oi_4 _495_ (.A1(_123_),
    .A2(_125_),
    .B1(net41),
    .Y(_126_));
 sky130_fd_sc_hd__mux2i_1 _496_ (.A0(\uart_rx_inst.bit_cnt[0] ),
    .A1(_122_),
    .S(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _497_ (.A(_117_),
    .B(_127_),
    .Y(_011_));
 sky130_fd_sc_hd__and3_1 _498_ (.A(_118_),
    .B(_083_),
    .C(_097_),
    .X(_128_));
 sky130_fd_sc_hd__or3b_1 _499_ (.A(_083_),
    .B(_084_),
    .C_N(_421_),
    .X(_129_));
 sky130_fd_sc_hd__buf_2 _500_ (.A(_129_),
    .X(_130_));
 sky130_fd_sc_hd__buf_2 _501_ (.A(_130_),
    .X(_131_));
 sky130_fd_sc_hd__o21ai_0 _502_ (.A1(_422_),
    .A2(_128_),
    .B1(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__mux2i_1 _503_ (.A0(\uart_rx_inst.bit_cnt[1] ),
    .A1(_132_),
    .S(_126_),
    .Y(_133_));
 sky130_fd_sc_hd__nor2_1 _504_ (.A(_117_),
    .B(_133_),
    .Y(_012_));
 sky130_fd_sc_hd__nor3_4 _505_ (.A(_094_),
    .B(_090_),
    .C(net40),
    .Y(_134_));
 sky130_fd_sc_hd__buf_6 _506_ (.A(_134_),
    .X(_135_));
 sky130_fd_sc_hd__o21ai_0 _507_ (.A1(_423_),
    .A2(_128_),
    .B1(net46),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(_084_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__buf_2 _509_ (.A(_130_),
    .X(_138_));
 sky130_fd_sc_hd__nand4b_1 _510_ (.A_N(_084_),
    .B(_423_),
    .C(_126_),
    .D(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__clkbuf_4 _511_ (.A(_100_),
    .X(_140_));
 sky130_fd_sc_hd__a21oi_1 _512_ (.A1(_137_),
    .A2(_139_),
    .B1(_140_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _513_ (.A(_118_),
    .B(_098_),
    .Y(_141_));
 sky130_fd_sc_hd__o31ai_1 _514_ (.A1(_084_),
    .A2(\uart_rx_inst.bit_cnt[1] ),
    .A3(\uart_rx_inst.bit_cnt[0] ),
    .B1(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__a21oi_1 _515_ (.A1(_420_),
    .A2(_419_),
    .B1(_421_),
    .Y(_143_));
 sky130_fd_sc_hd__nor2_1 _516_ (.A(_084_),
    .B(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__a21oi_1 _517_ (.A1(_126_),
    .A2(_144_),
    .B1(_083_),
    .Y(_145_));
 sky130_fd_sc_hd__a311oi_1 _518_ (.A1(_083_),
    .A2(net46),
    .A3(_142_),
    .B1(_145_),
    .C1(_100_),
    .Y(_014_));
 sky130_fd_sc_hd__or3_1 _519_ (.A(_118_),
    .B(_095_),
    .C(_130_),
    .X(_146_));
 sky130_fd_sc_hd__buf_6 _520_ (.A(_095_),
    .X(_147_));
 sky130_fd_sc_hd__o21ai_0 _521_ (.A1(_147_),
    .A2(_138_),
    .B1(net34),
    .Y(_148_));
 sky130_fd_sc_hd__a21oi_1 _522_ (.A1(_146_),
    .A2(_148_),
    .B1(_140_),
    .Y(_015_));
 sky130_fd_sc_hd__and2_0 _523_ (.A(\uart_rx_inst.data_reg[1] ),
    .B(_138_),
    .X(_016_));
 sky130_fd_sc_hd__and2_0 _524_ (.A(\uart_rx_inst.data_reg[2] ),
    .B(_138_),
    .X(_017_));
 sky130_fd_sc_hd__and2_0 _525_ (.A(\uart_rx_inst.data_reg[3] ),
    .B(_138_),
    .X(_018_));
 sky130_fd_sc_hd__and2_0 _526_ (.A(\uart_rx_inst.data_reg[4] ),
    .B(_138_),
    .X(_019_));
 sky130_fd_sc_hd__and2_0 _527_ (.A(\uart_rx_inst.data_reg[5] ),
    .B(_138_),
    .X(_020_));
 sky130_fd_sc_hd__and2_0 _528_ (.A(\uart_rx_inst.data_reg[6] ),
    .B(_138_),
    .X(_021_));
 sky130_fd_sc_hd__and2_0 _529_ (.A(\uart_rx_inst.data_reg[7] ),
    .B(_138_),
    .X(_022_));
 sky130_fd_sc_hd__and2_0 _530_ (.A(_118_),
    .B(_138_),
    .X(_023_));
 sky130_fd_sc_hd__nand3_1 _531_ (.A(_425_),
    .B(_123_),
    .C(_085_),
    .Y(_149_));
 sky130_fd_sc_hd__nor3_1 _532_ (.A(_118_),
    .B(_099_),
    .C(_149_),
    .Y(_024_));
 sky130_fd_sc_hd__nand4_1 _533_ (.A(_118_),
    .B(\uart_rx_inst.bit_cnt[0] ),
    .C(_123_),
    .D(_085_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_8 _534_ (.A(net41),
    .B(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__mux2i_1 _535_ (.A0(net25),
    .A1(\uart_rx_inst.data_reg[0] ),
    .S(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(_117_),
    .B(_152_),
    .Y(_025_));
 sky130_fd_sc_hd__mux2i_1 _537_ (.A0(net26),
    .A1(\uart_rx_inst.data_reg[1] ),
    .S(_151_),
    .Y(_153_));
 sky130_fd_sc_hd__nor2_1 _538_ (.A(_117_),
    .B(_153_),
    .Y(_026_));
 sky130_fd_sc_hd__mux2i_1 _539_ (.A0(net27),
    .A1(\uart_rx_inst.data_reg[2] ),
    .S(_151_),
    .Y(_154_));
 sky130_fd_sc_hd__nor2_1 _540_ (.A(_117_),
    .B(_154_),
    .Y(_027_));
 sky130_fd_sc_hd__mux2i_1 _541_ (.A0(net28),
    .A1(\uart_rx_inst.data_reg[3] ),
    .S(_151_),
    .Y(_155_));
 sky130_fd_sc_hd__nor2_1 _542_ (.A(_117_),
    .B(_155_),
    .Y(_028_));
 sky130_fd_sc_hd__mux2i_1 _543_ (.A0(net29),
    .A1(\uart_rx_inst.data_reg[4] ),
    .S(_151_),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_1 _544_ (.A(_117_),
    .B(_156_),
    .Y(_029_));
 sky130_fd_sc_hd__mux2i_1 _545_ (.A0(net30),
    .A1(\uart_rx_inst.data_reg[5] ),
    .S(_151_),
    .Y(_157_));
 sky130_fd_sc_hd__nor2_1 _546_ (.A(_117_),
    .B(_157_),
    .Y(_030_));
 sky130_fd_sc_hd__mux2i_1 _547_ (.A0(net31),
    .A1(\uart_rx_inst.data_reg[6] ),
    .S(_151_),
    .Y(_158_));
 sky130_fd_sc_hd__nor2_1 _548_ (.A(_117_),
    .B(_158_),
    .Y(_031_));
 sky130_fd_sc_hd__mux2i_1 _549_ (.A0(net32),
    .A1(\uart_rx_inst.data_reg[7] ),
    .S(_151_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _550_ (.A(_117_),
    .B(_159_),
    .Y(_032_));
 sky130_fd_sc_hd__nand4_1 _551_ (.A(_118_),
    .B(_425_),
    .C(_123_),
    .D(_085_),
    .Y(_160_));
 sky130_fd_sc_hd__inv_1 _552_ (.A(net33),
    .Y(_161_));
 sky130_fd_sc_hd__o32a_1 _553_ (.A1(net2),
    .A2(_098_),
    .A3(_160_),
    .B1(net1),
    .B2(_161_),
    .X(_162_));
 sky130_fd_sc_hd__nor2_1 _554_ (.A(_140_),
    .B(_162_),
    .Y(_033_));
 sky130_fd_sc_hd__nor3_1 _555_ (.A(_161_),
    .B(_099_),
    .C(_160_),
    .Y(_034_));
 sky130_fd_sc_hd__a21o_1 _556_ (.A1(_087_),
    .A2(_134_),
    .B1(net14),
    .X(_163_));
 sky130_fd_sc_hd__buf_6 _557_ (.A(_163_),
    .X(_164_));
 sky130_fd_sc_hd__buf_8 _558_ (.A(_164_),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_4 _559_ (.A(net2),
    .X(_166_));
 sky130_fd_sc_hd__nor2_1 _560_ (.A(_147_),
    .B(_121_),
    .Y(_167_));
 sky130_fd_sc_hd__a21oi_1 _561_ (.A1(_411_),
    .A2(_166_),
    .B1(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__nor2_1 _562_ (.A(_165_),
    .B(_168_),
    .Y(_035_));
 sky130_fd_sc_hd__and3b_1 _563_ (.A_N(\uart_rx_inst.prescale_reg[5] ),
    .B(_413_),
    .C(_091_),
    .X(_169_));
 sky130_fd_sc_hd__nand2_2 _564_ (.A(_093_),
    .B(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__xor2_1 _565_ (.A(\uart_rx_inst.prescale_reg[10] ),
    .B(_170_),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_4 _566_ (.A(prescale[4]),
    .X(_172_));
 sky130_fd_sc_hd__buf_2 _567_ (.A(prescale[5]),
    .X(_173_));
 sky130_fd_sc_hd__buf_2 _568_ (.A(prescale[3]),
    .X(_174_));
 sky130_fd_sc_hd__or3b_4 _569_ (.A(net10),
    .B(_174_),
    .C_N(_417_),
    .X(_175_));
 sky130_fd_sc_hd__nor3_4 _570_ (.A(_175_),
    .B(_173_),
    .C(_172_),
    .Y(_176_));
 sky130_fd_sc_hd__buf_2 _571_ (.A(prescale[6]),
    .X(_177_));
 sky130_fd_sc_hd__nor2_1 _572_ (.A(_177_),
    .B(net11),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _573_ (.A(_176_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__xor2_1 _574_ (.A(net12),
    .B(_179_),
    .X(_180_));
 sky130_fd_sc_hd__nor3_2 _575_ (.A(_174_),
    .B(_172_),
    .C(_173_),
    .Y(_181_));
 sky130_fd_sc_hd__nor3_4 _576_ (.A(net3),
    .B(net10),
    .C(net9),
    .Y(_182_));
 sky130_fd_sc_hd__nand2_1 _577_ (.A(_181_),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__nor2_1 _578_ (.A(_177_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__xnor2_1 _579_ (.A(net11),
    .B(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__o221a_1 _580_ (.A1(_130_),
    .A2(_180_),
    .B1(_185_),
    .B2(_120_),
    .C1(net47),
    .X(_186_));
 sky130_fd_sc_hd__a211oi_1 _581_ (.A1(_166_),
    .A2(_171_),
    .B1(_186_),
    .C1(_165_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _582_ (.A(\uart_rx_inst.prescale_reg[10] ),
    .B(_094_),
    .Y(_187_));
 sky130_fd_sc_hd__xnor2_1 _583_ (.A(net43),
    .B(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__nand4b_1 _584_ (.A_N(net12),
    .B(_181_),
    .C(_178_),
    .D(_182_),
    .Y(_189_));
 sky130_fd_sc_hd__xor2_1 _585_ (.A(net13),
    .B(_189_),
    .X(_190_));
 sky130_fd_sc_hd__o221a_1 _586_ (.A1(_120_),
    .A2(_180_),
    .B1(_190_),
    .B2(_131_),
    .C1(_135_),
    .X(_191_));
 sky130_fd_sc_hd__nor3_1 _587_ (.A(_164_),
    .B(_188_),
    .C(_191_),
    .Y(_037_));
 sky130_fd_sc_hd__nor3_1 _588_ (.A(net44),
    .B(\uart_rx_inst.prescale_reg[10] ),
    .C(_170_),
    .Y(_192_));
 sky130_fd_sc_hd__xnor2_1 _589_ (.A(\uart_rx_inst.prescale_reg[12] ),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__nor3b_2 _590_ (.A(net10),
    .B(_174_),
    .C_N(_417_),
    .Y(_194_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_172_),
    .B(_173_),
    .Y(_195_));
 sky130_fd_sc_hd__nor4_4 _592_ (.A(_177_),
    .B(net11),
    .C(net12),
    .D(net13),
    .Y(_196_));
 sky130_fd_sc_hd__nand3_1 _593_ (.A(_194_),
    .B(_195_),
    .C(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__xor2_1 _594_ (.A(net4),
    .B(_197_),
    .X(_198_));
 sky130_fd_sc_hd__o22ai_1 _595_ (.A1(_120_),
    .A2(_190_),
    .B1(_198_),
    .B2(_131_),
    .Y(_199_));
 sky130_fd_sc_hd__nor2_1 _596_ (.A(_147_),
    .B(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__a211oi_1 _597_ (.A1(_166_),
    .A2(_193_),
    .B1(_200_),
    .C1(_164_),
    .Y(_038_));
 sky130_fd_sc_hd__nor4_1 _598_ (.A(net49),
    .B(\uart_rx_inst.prescale_reg[12] ),
    .C(\uart_rx_inst.prescale_reg[10] ),
    .D(_094_),
    .Y(_201_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(net42),
    .B(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__clkbuf_2 _600_ (.A(prescale[11]),
    .X(_203_));
 sky130_fd_sc_hd__nand4b_4 _601_ (.A_N(net4),
    .B(_181_),
    .C(_182_),
    .D(_196_),
    .Y(_204_));
 sky130_fd_sc_hd__xor2_1 _602_ (.A(_203_),
    .B(_204_),
    .X(_205_));
 sky130_fd_sc_hd__o22ai_1 _603_ (.A1(_121_),
    .A2(_198_),
    .B1(_205_),
    .B2(_131_),
    .Y(_206_));
 sky130_fd_sc_hd__nor2_1 _604_ (.A(_166_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__nor3_1 _605_ (.A(_164_),
    .B(_202_),
    .C(_207_),
    .Y(_039_));
 sky130_fd_sc_hd__nor2_1 _606_ (.A(_088_),
    .B(_170_),
    .Y(_208_));
 sky130_fd_sc_hd__xnor2_1 _607_ (.A(\uart_rx_inst.prescale_reg[14] ),
    .B(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__nor2_1 _608_ (.A(net4),
    .B(_203_),
    .Y(_210_));
 sky130_fd_sc_hd__nand4_1 _609_ (.A(_194_),
    .B(_195_),
    .C(_196_),
    .D(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__xor2_1 _610_ (.A(net5),
    .B(_211_),
    .X(_212_));
 sky130_fd_sc_hd__o22ai_1 _611_ (.A1(_120_),
    .A2(_205_),
    .B1(_212_),
    .B2(_131_),
    .Y(_213_));
 sky130_fd_sc_hd__nor2_1 _612_ (.A(_147_),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__a211oi_1 _613_ (.A1(_166_),
    .A2(_209_),
    .B1(_214_),
    .C1(_164_),
    .Y(_040_));
 sky130_fd_sc_hd__nor3_1 _614_ (.A(net4),
    .B(_203_),
    .C(net5),
    .Y(_215_));
 sky130_fd_sc_hd__nand4_1 _615_ (.A(_181_),
    .B(_182_),
    .C(_196_),
    .D(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_1 _616_ (.A(net6),
    .B(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__a21oi_1 _617_ (.A1(_119_),
    .A2(_217_),
    .B1(_090_),
    .Y(_218_));
 sky130_fd_sc_hd__or3_1 _618_ (.A(\uart_rx_inst.prescale_reg[14] ),
    .B(_088_),
    .C(_094_),
    .X(_219_));
 sky130_fd_sc_hd__or3_1 _619_ (.A(\uart_rx_inst.prescale_reg[15] ),
    .B(_218_),
    .C(_219_),
    .X(_220_));
 sky130_fd_sc_hd__nor3_1 _620_ (.A(_147_),
    .B(_121_),
    .C(_212_),
    .Y(_221_));
 sky130_fd_sc_hd__a21oi_1 _621_ (.A1(\uart_rx_inst.prescale_reg[15] ),
    .A2(_219_),
    .B1(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__a21oi_1 _622_ (.A1(_220_),
    .A2(_222_),
    .B1(_165_),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _623_ (.A(_089_),
    .B(_170_),
    .Y(_223_));
 sky130_fd_sc_hd__xnor2_1 _624_ (.A(\uart_rx_inst.prescale_reg[16] ),
    .B(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__nor2b_1 _625_ (.A(net4),
    .B_N(_196_),
    .Y(_225_));
 sky130_fd_sc_hd__nor3_1 _626_ (.A(_203_),
    .B(net5),
    .C(net6),
    .Y(_226_));
 sky130_fd_sc_hd__nand3_1 _627_ (.A(_176_),
    .B(_225_),
    .C(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__xor2_1 _628_ (.A(net7),
    .B(_227_),
    .X(_228_));
 sky130_fd_sc_hd__nor2_1 _629_ (.A(_087_),
    .B(net2),
    .Y(_229_));
 sky130_fd_sc_hd__o21a_1 _630_ (.A1(_130_),
    .A2(_228_),
    .B1(_229_),
    .X(_230_));
 sky130_fd_sc_hd__a31oi_4 _631_ (.A1(_118_),
    .A2(_083_),
    .A3(_097_),
    .B1(_119_),
    .Y(_231_));
 sky130_fd_sc_hd__nand2_1 _632_ (.A(_231_),
    .B(_217_),
    .Y(_232_));
 sky130_fd_sc_hd__a221oi_1 _633_ (.A1(_166_),
    .A2(_224_),
    .B1(_230_),
    .B2(_232_),
    .C1(_164_),
    .Y(_042_));
 sky130_fd_sc_hd__nor2b_1 _634_ (.A(\uart_rx_inst.prescale_reg[17] ),
    .B_N(\uart_rx_inst.prescale_reg[18] ),
    .Y(_233_));
 sky130_fd_sc_hd__or3_1 _635_ (.A(\uart_rx_inst.prescale_reg[16] ),
    .B(_089_),
    .C(_094_),
    .X(_234_));
 sky130_fd_sc_hd__mux2i_1 _636_ (.A0(_233_),
    .A1(\uart_rx_inst.prescale_reg[17] ),
    .S(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__nand2b_1 _637_ (.A_N(net7),
    .B(_226_),
    .Y(_236_));
 sky130_fd_sc_hd__o21ai_0 _638_ (.A1(_204_),
    .A2(_236_),
    .B1(net8),
    .Y(_237_));
 sky130_fd_sc_hd__or3_1 _639_ (.A(net8),
    .B(_204_),
    .C(_236_),
    .X(_238_));
 sky130_fd_sc_hd__a211o_1 _640_ (.A1(_237_),
    .A2(_238_),
    .B1(net2),
    .C1(_130_),
    .X(_239_));
 sky130_fd_sc_hd__or4_1 _641_ (.A(\uart_rx_inst.prescale_reg[17] ),
    .B(_120_),
    .C(_228_),
    .D(_234_),
    .X(_240_));
 sky130_fd_sc_hd__a31oi_1 _642_ (.A1(_235_),
    .A2(_239_),
    .A3(_240_),
    .B1(_165_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _643_ (.A(_176_),
    .B(_225_),
    .Y(_241_));
 sky130_fd_sc_hd__nor4_1 _644_ (.A(net8),
    .B(_130_),
    .C(_241_),
    .D(_236_),
    .Y(_242_));
 sky130_fd_sc_hd__a21oi_1 _645_ (.A1(_237_),
    .A2(_238_),
    .B1(_121_),
    .Y(_243_));
 sky130_fd_sc_hd__o21ai_1 _646_ (.A1(_242_),
    .A2(_243_),
    .B1(net46),
    .Y(_244_));
 sky130_fd_sc_hd__a31oi_1 _647_ (.A1(_091_),
    .A2(_092_),
    .A3(_093_),
    .B1(\uart_rx_inst.prescale_reg[18] ),
    .Y(_245_));
 sky130_fd_sc_hd__nor4_1 _648_ (.A(\uart_rx_inst.prescale_reg[17] ),
    .B(\uart_rx_inst.prescale_reg[16] ),
    .C(_089_),
    .D(_170_),
    .Y(_246_));
 sky130_fd_sc_hd__mux2i_1 _649_ (.A0(\uart_rx_inst.prescale_reg[18] ),
    .A1(_245_),
    .S(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__a21oi_1 _650_ (.A1(_244_),
    .A2(_247_),
    .B1(_165_),
    .Y(_044_));
 sky130_fd_sc_hd__nor2_1 _651_ (.A(_147_),
    .B(_141_),
    .Y(_248_));
 sky130_fd_sc_hd__a211oi_1 _652_ (.A1(_414_),
    .A2(_166_),
    .B1(_164_),
    .C1(_248_),
    .Y(_045_));
 sky130_fd_sc_hd__xnor2_1 _653_ (.A(\uart_rx_inst.prescale_reg[2] ),
    .B(_413_),
    .Y(_249_));
 sky130_fd_sc_hd__a211oi_1 _654_ (.A1(_415_),
    .A2(_119_),
    .B1(_231_),
    .C1(_147_),
    .Y(_250_));
 sky130_fd_sc_hd__a211oi_1 _655_ (.A1(_166_),
    .A2(_249_),
    .B1(_250_),
    .C1(_164_),
    .Y(_046_));
 sky130_fd_sc_hd__o22ai_1 _656_ (.A1(_418_),
    .A2(_131_),
    .B1(_121_),
    .B2(net3),
    .Y(_251_));
 sky130_fd_sc_hd__nor3_1 _657_ (.A(\uart_rx_inst.prescale_reg[2] ),
    .B(\uart_rx_inst.prescale_reg[1] ),
    .C(\uart_rx_inst.prescale_reg[0] ),
    .Y(_252_));
 sky130_fd_sc_hd__xor2_1 _658_ (.A(\uart_rx_inst.prescale_reg[3] ),
    .B(_252_),
    .X(_253_));
 sky130_fd_sc_hd__o21ai_0 _659_ (.A1(_166_),
    .A2(_251_),
    .B1(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__nor2_1 _660_ (.A(_165_),
    .B(_254_),
    .Y(_047_));
 sky130_fd_sc_hd__nor2_1 _661_ (.A(\uart_rx_inst.prescale_reg[3] ),
    .B(\uart_rx_inst.prescale_reg[2] ),
    .Y(_255_));
 sky130_fd_sc_hd__nand2_1 _662_ (.A(_413_),
    .B(_255_),
    .Y(_256_));
 sky130_fd_sc_hd__xnor2_1 _663_ (.A(\uart_rx_inst.prescale_reg[4] ),
    .B(_256_),
    .Y(_257_));
 sky130_fd_sc_hd__xnor2_1 _664_ (.A(net10),
    .B(_417_),
    .Y(_258_));
 sky130_fd_sc_hd__o221ai_1 _665_ (.A1(_418_),
    .A2(_121_),
    .B1(_258_),
    .B2(_131_),
    .C1(_135_),
    .Y(_259_));
 sky130_fd_sc_hd__o21ai_0 _666_ (.A1(net46),
    .A2(_257_),
    .B1(_259_),
    .Y(_260_));
 sky130_fd_sc_hd__nor2_1 _667_ (.A(_165_),
    .B(_260_),
    .Y(_048_));
 sky130_fd_sc_hd__xnor2_1 _668_ (.A(_174_),
    .B(_182_),
    .Y(_261_));
 sky130_fd_sc_hd__nor3_1 _669_ (.A(_128_),
    .B(_119_),
    .C(_258_),
    .Y(_262_));
 sky130_fd_sc_hd__o21bai_1 _670_ (.A1(_130_),
    .A2(_261_),
    .B1_N(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__nand3_1 _671_ (.A(_412_),
    .B(_411_),
    .C(_091_),
    .Y(_264_));
 sky130_fd_sc_hd__a21o_1 _672_ (.A1(_087_),
    .A2(_134_),
    .B1(_264_),
    .X(_265_));
 sky130_fd_sc_hd__nand2_1 _673_ (.A(_091_),
    .B(_092_),
    .Y(_266_));
 sky130_fd_sc_hd__nor2_1 _674_ (.A(_266_),
    .B(_135_),
    .Y(_267_));
 sky130_fd_sc_hd__a221oi_1 _675_ (.A1(_229_),
    .A2(_263_),
    .B1(_265_),
    .B2(\uart_rx_inst.prescale_reg[5] ),
    .C1(_267_),
    .Y(_268_));
 sky130_fd_sc_hd__nor2_1 _676_ (.A(_140_),
    .B(_268_),
    .Y(_049_));
 sky130_fd_sc_hd__xor2_1 _677_ (.A(\uart_rx_inst.prescale_reg[6] ),
    .B(_169_),
    .X(_269_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(_172_),
    .B(_194_),
    .Y(_270_));
 sky130_fd_sc_hd__o221ai_1 _679_ (.A1(_121_),
    .A2(_261_),
    .B1(_270_),
    .B2(_131_),
    .C1(_135_),
    .Y(_271_));
 sky130_fd_sc_hd__o21ai_0 _680_ (.A1(net46),
    .A2(_269_),
    .B1(_271_),
    .Y(_272_));
 sky130_fd_sc_hd__nor2_1 _681_ (.A(_165_),
    .B(_272_),
    .Y(_050_));
 sky130_fd_sc_hd__nor2_1 _682_ (.A(_174_),
    .B(_172_),
    .Y(_273_));
 sky130_fd_sc_hd__nand2_1 _683_ (.A(_273_),
    .B(_182_),
    .Y(_274_));
 sky130_fd_sc_hd__xor2_1 _684_ (.A(_173_),
    .B(_274_),
    .X(_275_));
 sky130_fd_sc_hd__o22ai_1 _685_ (.A1(_121_),
    .A2(_270_),
    .B1(_275_),
    .B2(_131_),
    .Y(_276_));
 sky130_fd_sc_hd__nor2_1 _686_ (.A(\uart_rx_inst.prescale_reg[6] ),
    .B(_266_),
    .Y(_277_));
 sky130_fd_sc_hd__xor2_1 _687_ (.A(\uart_rx_inst.prescale_reg[7] ),
    .B(_277_),
    .X(_278_));
 sky130_fd_sc_hd__o21ai_0 _688_ (.A1(_166_),
    .A2(_276_),
    .B1(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__nor2_1 _689_ (.A(_165_),
    .B(_279_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _690_ (.A(\uart_rx_inst.prescale_reg[7] ),
    .B(\uart_rx_inst.prescale_reg[6] ),
    .Y(_280_));
 sky130_fd_sc_hd__nand2_1 _691_ (.A(_280_),
    .B(_169_),
    .Y(_281_));
 sky130_fd_sc_hd__xnor2_1 _692_ (.A(\uart_rx_inst.prescale_reg[8] ),
    .B(_281_),
    .Y(_282_));
 sky130_fd_sc_hd__nor3_1 _693_ (.A(_147_),
    .B(_121_),
    .C(_275_),
    .Y(_283_));
 sky130_fd_sc_hd__xnor2_1 _694_ (.A(_177_),
    .B(net48),
    .Y(_284_));
 sky130_fd_sc_hd__nor3_1 _695_ (.A(_147_),
    .B(_131_),
    .C(_284_),
    .Y(_285_));
 sky130_fd_sc_hd__a211oi_1 _696_ (.A1(_147_),
    .A2(_282_),
    .B1(_283_),
    .C1(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__nor2_1 _697_ (.A(_165_),
    .B(_286_),
    .Y(_052_));
 sky130_fd_sc_hd__nand2_1 _698_ (.A(_194_),
    .B(_195_),
    .Y(_287_));
 sky130_fd_sc_hd__o32a_1 _699_ (.A1(net11),
    .A2(_130_),
    .A3(_183_),
    .B1(_287_),
    .B2(_120_),
    .X(_288_));
 sky130_fd_sc_hd__inv_1 _700_ (.A(_177_),
    .Y(_289_));
 sky130_fd_sc_hd__inv_1 _701_ (.A(net11),
    .Y(_290_));
 sky130_fd_sc_hd__a311oi_1 _702_ (.A1(_289_),
    .A2(_181_),
    .A3(_182_),
    .B1(_290_),
    .C1(_130_),
    .Y(_291_));
 sky130_fd_sc_hd__a31oi_1 _703_ (.A1(_177_),
    .A2(_231_),
    .A3(_287_),
    .B1(_291_),
    .Y(_292_));
 sky130_fd_sc_hd__o21ai_0 _704_ (.A1(_177_),
    .A2(_288_),
    .B1(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__o41ai_1 _705_ (.A1(\uart_rx_inst.prescale_reg[7] ),
    .A2(\uart_rx_inst.prescale_reg[8] ),
    .A3(\uart_rx_inst.prescale_reg[6] ),
    .A4(_266_),
    .B1(\uart_rx_inst.prescale_reg[9] ),
    .Y(_294_));
 sky130_fd_sc_hd__o21ai_0 _706_ (.A1(_094_),
    .A2(_135_),
    .B1(_294_),
    .Y(_295_));
 sky130_fd_sc_hd__a21oi_1 _707_ (.A1(_229_),
    .A2(_293_),
    .B1(_295_),
    .Y(_296_));
 sky130_fd_sc_hd__nor2_1 _708_ (.A(_140_),
    .B(_296_),
    .Y(_053_));
 sky130_fd_sc_hd__or2_0 _709_ (.A(_100_),
    .B(net15),
    .X(_054_));
 sky130_fd_sc_hd__nor2b_2 _710_ (.A(net24),
    .B_N(_082_),
    .Y(_297_));
 sky130_fd_sc_hd__or2_0 _711_ (.A(_107_),
    .B(_111_),
    .X(_298_));
 sky130_fd_sc_hd__buf_2 _712_ (.A(_298_),
    .X(_299_));
 sky130_fd_sc_hd__nor2_1 _713_ (.A(_297_),
    .B(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__buf_2 _714_ (.A(_300_),
    .X(_301_));
 sky130_fd_sc_hd__buf_2 _715_ (.A(_299_),
    .X(_302_));
 sky130_fd_sc_hd__mux2i_1 _716_ (.A0(_301_),
    .A1(_302_),
    .S(_081_),
    .Y(_303_));
 sky130_fd_sc_hd__nor2_1 _717_ (.A(_140_),
    .B(_303_),
    .Y(_055_));
 sky130_fd_sc_hd__o21ai_0 _718_ (.A1(_081_),
    .A2(_302_),
    .B1(\uart_tx_inst.bit_cnt[1] ),
    .Y(_304_));
 sky130_fd_sc_hd__or4_1 _719_ (.A(\uart_tx_inst.bit_cnt[1] ),
    .B(_081_),
    .C(_082_),
    .D(_299_),
    .X(_305_));
 sky130_fd_sc_hd__a21oi_1 _720_ (.A1(_304_),
    .A2(_305_),
    .B1(_140_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2b_1 _721_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .B_N(\uart_tx_inst.bit_cnt[3] ),
    .Y(_306_));
 sky130_fd_sc_hd__nor3_1 _722_ (.A(\uart_tx_inst.bit_cnt[1] ),
    .B(_081_),
    .C(_299_),
    .Y(_307_));
 sky130_fd_sc_hd__mux2i_1 _723_ (.A0(\uart_tx_inst.bit_cnt[2] ),
    .A1(_306_),
    .S(_307_),
    .Y(_308_));
 sky130_fd_sc_hd__nor2_1 _724_ (.A(_140_),
    .B(_308_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2b_1 _725_ (.A(\uart_tx_inst.bit_cnt[3] ),
    .B_N(net24),
    .Y(_309_));
 sky130_fd_sc_hd__nor4_1 _726_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .B(\uart_tx_inst.bit_cnt[1] ),
    .C(_081_),
    .D(_299_),
    .Y(_310_));
 sky130_fd_sc_hd__mux2i_1 _727_ (.A0(\uart_tx_inst.bit_cnt[3] ),
    .A1(_309_),
    .S(_310_),
    .Y(_311_));
 sky130_fd_sc_hd__nor2_1 _728_ (.A(_140_),
    .B(_311_),
    .Y(_058_));
 sky130_fd_sc_hd__a21o_2 _729_ (.A1(_297_),
    .A2(_113_),
    .B1(_100_),
    .X(_312_));
 sky130_fd_sc_hd__a21oi_1 _730_ (.A1(_002_),
    .A2(_113_),
    .B1(net38),
    .Y(_313_));
 sky130_fd_sc_hd__nor2_1 _731_ (.A(_312_),
    .B(_313_),
    .Y(_059_));
 sky130_fd_sc_hd__nor3_1 _732_ (.A(\uart_tx_inst.bit_cnt[2] ),
    .B(\uart_tx_inst.bit_cnt[3] ),
    .C(\uart_tx_inst.bit_cnt[1] ),
    .Y(_314_));
 sky130_fd_sc_hd__nand2_2 _733_ (.A(_081_),
    .B(_314_),
    .Y(_315_));
 sky130_fd_sc_hd__a21oi_1 _734_ (.A1(_297_),
    .A2(_113_),
    .B1(_100_),
    .Y(_316_));
 sky130_fd_sc_hd__o21ai_2 _735_ (.A1(_299_),
    .A2(_315_),
    .B1(_316_),
    .Y(_317_));
 sky130_fd_sc_hd__nor2_1 _736_ (.A(\uart_tx_inst.prescale_reg[0] ),
    .B(_317_),
    .Y(_060_));
 sky130_fd_sc_hd__and3_1 _737_ (.A(_429_),
    .B(_103_),
    .C(_105_),
    .X(_318_));
 sky130_fd_sc_hd__nand2_1 _738_ (.A(_106_),
    .B(_318_),
    .Y(_319_));
 sky130_fd_sc_hd__o21ai_0 _739_ (.A1(\uart_tx_inst.prescale_reg[9] ),
    .A2(_319_),
    .B1(\uart_tx_inst.prescale_reg[10] ),
    .Y(_320_));
 sky130_fd_sc_hd__or4_1 _740_ (.A(\uart_tx_inst.prescale_reg[10] ),
    .B(\uart_tx_inst.prescale_reg[9] ),
    .C(_112_),
    .D(_319_),
    .X(_321_));
 sky130_fd_sc_hd__nor3_1 _741_ (.A(_177_),
    .B(_116_),
    .C(_183_),
    .Y(_322_));
 sky130_fd_sc_hd__xnor2_1 _742_ (.A(_290_),
    .B(_322_),
    .Y(_323_));
 sky130_fd_sc_hd__nand2_1 _743_ (.A(_301_),
    .B(_323_),
    .Y(_324_));
 sky130_fd_sc_hd__a31oi_1 _744_ (.A1(_320_),
    .A2(_321_),
    .A3(_324_),
    .B1(_101_),
    .Y(_061_));
 sky130_fd_sc_hd__nor4_4 _745_ (.A(_172_),
    .B(_173_),
    .C(_115_),
    .D(_175_),
    .Y(_325_));
 sky130_fd_sc_hd__nand2_1 _746_ (.A(_178_),
    .B(_325_),
    .Y(_326_));
 sky130_fd_sc_hd__xnor2_1 _747_ (.A(net12),
    .B(_326_),
    .Y(_327_));
 sky130_fd_sc_hd__nand2_1 _748_ (.A(_301_),
    .B(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__or3_1 _749_ (.A(\uart_tx_inst.prescale_reg[10] ),
    .B(\uart_tx_inst.prescale_reg[9] ),
    .C(_107_),
    .X(_329_));
 sky130_fd_sc_hd__nand2b_1 _750_ (.A_N(_329_),
    .B(_299_),
    .Y(_330_));
 sky130_fd_sc_hd__xor2_1 _751_ (.A(\uart_tx_inst.prescale_reg[11] ),
    .B(_330_),
    .X(_331_));
 sky130_fd_sc_hd__a21oi_1 _752_ (.A1(_328_),
    .A2(_331_),
    .B1(_140_),
    .Y(_062_));
 sky130_fd_sc_hd__and2_0 _753_ (.A(_106_),
    .B(_318_),
    .X(_332_));
 sky130_fd_sc_hd__a311o_1 _754_ (.A1(_109_),
    .A2(_299_),
    .A3(_332_),
    .B1(_300_),
    .C1(\uart_tx_inst.prescale_reg[12] ),
    .X(_333_));
 sky130_fd_sc_hd__nand2b_1 _755_ (.A_N(_189_),
    .B(_315_),
    .Y(_334_));
 sky130_fd_sc_hd__xor2_1 _756_ (.A(net13),
    .B(_334_),
    .X(_335_));
 sky130_fd_sc_hd__nand2_1 _757_ (.A(_301_),
    .B(_335_),
    .Y(_336_));
 sky130_fd_sc_hd__a31oi_1 _758_ (.A1(\uart_tx_inst.prescale_reg[12] ),
    .A2(_109_),
    .A3(_332_),
    .B1(_100_),
    .Y(_337_));
 sky130_fd_sc_hd__and3_1 _759_ (.A(_333_),
    .B(_336_),
    .C(_337_),
    .X(_063_));
 sky130_fd_sc_hd__and3_1 _760_ (.A(_103_),
    .B(_104_),
    .C(_105_),
    .X(_338_));
 sky130_fd_sc_hd__and2_0 _761_ (.A(_109_),
    .B(_110_),
    .X(_339_));
 sky130_fd_sc_hd__nand3_1 _762_ (.A(_338_),
    .B(_106_),
    .C(_339_),
    .Y(_340_));
 sky130_fd_sc_hd__o31ai_1 _763_ (.A1(\uart_tx_inst.prescale_reg[12] ),
    .A2(\uart_tx_inst.prescale_reg[11] ),
    .A3(_329_),
    .B1(\uart_tx_inst.prescale_reg[13] ),
    .Y(_341_));
 sky130_fd_sc_hd__nand2_1 _764_ (.A(_196_),
    .B(_325_),
    .Y(_342_));
 sky130_fd_sc_hd__xor2_1 _765_ (.A(net4),
    .B(_342_),
    .X(_343_));
 sky130_fd_sc_hd__a221oi_1 _766_ (.A1(_340_),
    .A2(_341_),
    .B1(_343_),
    .B2(_301_),
    .C1(_312_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2_1 _767_ (.A(_116_),
    .B(_204_),
    .Y(_344_));
 sky130_fd_sc_hd__xor2_1 _768_ (.A(_203_),
    .B(_344_),
    .X(_345_));
 sky130_fd_sc_hd__nand2_1 _769_ (.A(_301_),
    .B(_345_),
    .Y(_346_));
 sky130_fd_sc_hd__nand3_1 _770_ (.A(_106_),
    .B(_339_),
    .C(_318_),
    .Y(_347_));
 sky130_fd_sc_hd__nor3_1 _771_ (.A(\uart_tx_inst.prescale_reg[14] ),
    .B(_113_),
    .C(_347_),
    .Y(_348_));
 sky130_fd_sc_hd__a21oi_1 _772_ (.A1(\uart_tx_inst.prescale_reg[14] ),
    .A2(_347_),
    .B1(_348_),
    .Y(_349_));
 sky130_fd_sc_hd__a21oi_1 _773_ (.A1(_346_),
    .A2(_349_),
    .B1(_101_),
    .Y(_065_));
 sky130_fd_sc_hd__nor3_1 _774_ (.A(\uart_tx_inst.prescale_reg[15] ),
    .B(\uart_tx_inst.prescale_reg[14] ),
    .C(_340_),
    .Y(_350_));
 sky130_fd_sc_hd__o41ai_1 _775_ (.A1(\uart_tx_inst.prescale_reg[18] ),
    .A2(\uart_tx_inst.prescale_reg[17] ),
    .A3(\uart_tx_inst.prescale_reg[16] ),
    .A4(_297_),
    .B1(_350_),
    .Y(_351_));
 sky130_fd_sc_hd__o21ai_0 _776_ (.A1(\uart_tx_inst.prescale_reg[14] ),
    .A2(_340_),
    .B1(\uart_tx_inst.prescale_reg[15] ),
    .Y(_352_));
 sky130_fd_sc_hd__nand3_1 _777_ (.A(_196_),
    .B(_210_),
    .C(_325_),
    .Y(_353_));
 sky130_fd_sc_hd__xnor2_1 _778_ (.A(net5),
    .B(_353_),
    .Y(_354_));
 sky130_fd_sc_hd__nand2_1 _779_ (.A(_113_),
    .B(_354_),
    .Y(_355_));
 sky130_fd_sc_hd__a31oi_1 _780_ (.A1(_351_),
    .A2(_352_),
    .A3(_355_),
    .B1(_312_),
    .Y(_066_));
 sky130_fd_sc_hd__nor3_1 _781_ (.A(\uart_tx_inst.prescale_reg[15] ),
    .B(\uart_tx_inst.prescale_reg[14] ),
    .C(_347_),
    .Y(_356_));
 sky130_fd_sc_hd__xnor2_1 _782_ (.A(\uart_tx_inst.prescale_reg[16] ),
    .B(_356_),
    .Y(_357_));
 sky130_fd_sc_hd__nand2_1 _783_ (.A(_113_),
    .B(_316_),
    .Y(_358_));
 sky130_fd_sc_hd__nor4_1 _784_ (.A(_203_),
    .B(net5),
    .C(_116_),
    .D(_204_),
    .Y(_359_));
 sky130_fd_sc_hd__xnor2_1 _785_ (.A(net6),
    .B(_359_),
    .Y(_360_));
 sky130_fd_sc_hd__o32ai_1 _786_ (.A1(_100_),
    .A2(_113_),
    .A3(_357_),
    .B1(_358_),
    .B2(_360_),
    .Y(_067_));
 sky130_fd_sc_hd__nor2_1 _787_ (.A(\uart_tx_inst.prescale_reg[18] ),
    .B(_297_),
    .Y(_361_));
 sky130_fd_sc_hd__nor2_1 _788_ (.A(\uart_tx_inst.prescale_reg[17] ),
    .B(_361_),
    .Y(_362_));
 sky130_fd_sc_hd__nor4_1 _789_ (.A(\uart_tx_inst.prescale_reg[15] ),
    .B(\uart_tx_inst.prescale_reg[16] ),
    .C(\uart_tx_inst.prescale_reg[14] ),
    .D(_340_),
    .Y(_363_));
 sky130_fd_sc_hd__mux2i_1 _790_ (.A0(\uart_tx_inst.prescale_reg[17] ),
    .A1(_362_),
    .S(_363_),
    .Y(_364_));
 sky130_fd_sc_hd__nand3_1 _791_ (.A(_225_),
    .B(_226_),
    .C(_325_),
    .Y(_365_));
 sky130_fd_sc_hd__xnor2_1 _792_ (.A(net7),
    .B(_365_),
    .Y(_366_));
 sky130_fd_sc_hd__nand2_1 _793_ (.A(_113_),
    .B(_366_),
    .Y(_367_));
 sky130_fd_sc_hd__a21oi_1 _794_ (.A1(_364_),
    .A2(_367_),
    .B1(_312_),
    .Y(_068_));
 sky130_fd_sc_hd__nand3_1 _795_ (.A(_108_),
    .B(_339_),
    .C(_332_),
    .Y(_368_));
 sky130_fd_sc_hd__nor4b_1 _796_ (.A(\uart_tx_inst.prescale_reg[18] ),
    .B(_338_),
    .C(_347_),
    .D_N(_108_),
    .Y(_369_));
 sky130_fd_sc_hd__a21oi_1 _797_ (.A1(\uart_tx_inst.prescale_reg[18] ),
    .A2(_368_),
    .B1(_369_),
    .Y(_370_));
 sky130_fd_sc_hd__nor3_1 _798_ (.A(_116_),
    .B(_204_),
    .C(_236_),
    .Y(_371_));
 sky130_fd_sc_hd__xnor2_1 _799_ (.A(net8),
    .B(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__o22ai_1 _800_ (.A1(_312_),
    .A2(_370_),
    .B1(_372_),
    .B2(_358_),
    .Y(_069_));
 sky130_fd_sc_hd__a21oi_1 _801_ (.A1(_430_),
    .A2(_302_),
    .B1(_317_),
    .Y(_070_));
 sky130_fd_sc_hd__xnor2_1 _802_ (.A(\uart_tx_inst.prescale_reg[2] ),
    .B(_429_),
    .Y(_373_));
 sky130_fd_sc_hd__a21oi_1 _803_ (.A1(_302_),
    .A2(_373_),
    .B1(_317_),
    .Y(_071_));
 sky130_fd_sc_hd__or3_1 _804_ (.A(\uart_tx_inst.prescale_reg[1] ),
    .B(\uart_tx_inst.prescale_reg[2] ),
    .C(\uart_tx_inst.prescale_reg[0] ),
    .X(_374_));
 sky130_fd_sc_hd__nor2_1 _805_ (.A(_374_),
    .B(_112_),
    .Y(_375_));
 sky130_fd_sc_hd__nand2_1 _806_ (.A(_415_),
    .B(_116_),
    .Y(_376_));
 sky130_fd_sc_hd__nand2_1 _807_ (.A(net3),
    .B(_315_),
    .Y(_377_));
 sky130_fd_sc_hd__a311oi_1 _808_ (.A1(_300_),
    .A2(_376_),
    .A3(_377_),
    .B1(_375_),
    .C1(\uart_tx_inst.prescale_reg[3] ),
    .Y(_378_));
 sky130_fd_sc_hd__a211oi_1 _809_ (.A1(\uart_tx_inst.prescale_reg[3] ),
    .A2(_375_),
    .B1(_378_),
    .C1(_101_),
    .Y(_072_));
 sky130_fd_sc_hd__and3_1 _810_ (.A(_429_),
    .B(_105_),
    .C(_299_),
    .X(_379_));
 sky130_fd_sc_hd__nand2_1 _811_ (.A(net9),
    .B(_116_),
    .Y(_380_));
 sky130_fd_sc_hd__o21ai_0 _812_ (.A1(_418_),
    .A2(_116_),
    .B1(_380_),
    .Y(_381_));
 sky130_fd_sc_hd__a211oi_1 _813_ (.A1(_301_),
    .A2(_381_),
    .B1(_379_),
    .C1(\uart_tx_inst.prescale_reg[4] ),
    .Y(_382_));
 sky130_fd_sc_hd__a211oi_1 _814_ (.A1(\uart_tx_inst.prescale_reg[4] ),
    .A2(_379_),
    .B1(_382_),
    .C1(_101_),
    .Y(_073_));
 sky130_fd_sc_hd__o41ai_1 _815_ (.A1(\uart_tx_inst.prescale_reg[4] ),
    .A2(\uart_tx_inst.prescale_reg[3] ),
    .A3(_374_),
    .A4(_113_),
    .B1(\uart_tx_inst.prescale_reg[5] ),
    .Y(_383_));
 sky130_fd_sc_hd__nand2_1 _816_ (.A(_417_),
    .B(_315_),
    .Y(_384_));
 sky130_fd_sc_hd__xnor2_1 _817_ (.A(net10),
    .B(_384_),
    .Y(_385_));
 sky130_fd_sc_hd__a22oi_1 _818_ (.A1(_338_),
    .A2(_302_),
    .B1(_301_),
    .B2(_385_),
    .Y(_386_));
 sky130_fd_sc_hd__a21oi_1 _819_ (.A1(_383_),
    .A2(_386_),
    .B1(_101_),
    .Y(_074_));
 sky130_fd_sc_hd__nand3_1 _820_ (.A(_429_),
    .B(_103_),
    .C(_105_),
    .Y(_387_));
 sky130_fd_sc_hd__nor2_1 _821_ (.A(_112_),
    .B(_387_),
    .Y(_388_));
 sky130_fd_sc_hd__nand2_1 _822_ (.A(_315_),
    .B(_182_),
    .Y(_389_));
 sky130_fd_sc_hd__xnor2_1 _823_ (.A(_174_),
    .B(_389_),
    .Y(_390_));
 sky130_fd_sc_hd__a211oi_1 _824_ (.A1(_301_),
    .A2(_390_),
    .B1(_388_),
    .C1(\uart_tx_inst.prescale_reg[6] ),
    .Y(_391_));
 sky130_fd_sc_hd__a211oi_1 _825_ (.A1(\uart_tx_inst.prescale_reg[6] ),
    .A2(_388_),
    .B1(_391_),
    .C1(_101_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _826_ (.A(_116_),
    .B(_175_),
    .Y(_392_));
 sky130_fd_sc_hd__xor2_1 _827_ (.A(_172_),
    .B(_392_),
    .X(_393_));
 sky130_fd_sc_hd__a21oi_1 _828_ (.A1(_102_),
    .A2(_393_),
    .B1(_302_),
    .Y(_394_));
 sky130_fd_sc_hd__nor2b_1 _829_ (.A(\uart_tx_inst.prescale_reg[6] ),
    .B_N(_338_),
    .Y(_395_));
 sky130_fd_sc_hd__xnor2_1 _830_ (.A(\uart_tx_inst.prescale_reg[7] ),
    .B(_395_),
    .Y(_396_));
 sky130_fd_sc_hd__nor3_1 _831_ (.A(_101_),
    .B(_394_),
    .C(_396_),
    .Y(_076_));
 sky130_fd_sc_hd__nor3_1 _832_ (.A(\uart_tx_inst.prescale_reg[7] ),
    .B(\uart_tx_inst.prescale_reg[6] ),
    .C(_387_),
    .Y(_397_));
 sky130_fd_sc_hd__xnor2_1 _833_ (.A(\uart_tx_inst.prescale_reg[8] ),
    .B(_397_),
    .Y(_398_));
 sky130_fd_sc_hd__nor2_1 _834_ (.A(_116_),
    .B(_274_),
    .Y(_399_));
 sky130_fd_sc_hd__xor2_1 _835_ (.A(_173_),
    .B(_399_),
    .X(_400_));
 sky130_fd_sc_hd__nor2_1 _836_ (.A(_302_),
    .B(_400_),
    .Y(_401_));
 sky130_fd_sc_hd__a211oi_1 _837_ (.A1(_302_),
    .A2(_398_),
    .B1(_401_),
    .C1(_312_),
    .Y(_077_));
 sky130_fd_sc_hd__xnor2_1 _838_ (.A(_289_),
    .B(_325_),
    .Y(_402_));
 sky130_fd_sc_hd__nand2_1 _839_ (.A(_301_),
    .B(_402_),
    .Y(_403_));
 sky130_fd_sc_hd__or3b_1 _840_ (.A(\uart_tx_inst.prescale_reg[9] ),
    .B(_107_),
    .C_N(_111_),
    .X(_404_));
 sky130_fd_sc_hd__nor2_1 _841_ (.A(_102_),
    .B(_111_),
    .Y(_405_));
 sky130_fd_sc_hd__o21ai_0 _842_ (.A1(_107_),
    .A2(_405_),
    .B1(\uart_tx_inst.prescale_reg[9] ),
    .Y(_406_));
 sky130_fd_sc_hd__a31oi_1 _843_ (.A1(_403_),
    .A2(_404_),
    .A3(_406_),
    .B1(_101_),
    .Y(_078_));
 sky130_fd_sc_hd__nand3_1 _844_ (.A(net24),
    .B(net37),
    .C(_002_),
    .Y(_407_));
 sky130_fd_sc_hd__o21ai_0 _845_ (.A1(net37),
    .A2(_002_),
    .B1(_407_),
    .Y(_408_));
 sky130_fd_sc_hd__nor3_1 _846_ (.A(_101_),
    .B(_302_),
    .C(_408_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2b_1 _847_ (.A_N(_314_),
    .B(\uart_tx_inst.data_reg[0] ),
    .Y(_409_));
 sky130_fd_sc_hd__a21oi_1 _848_ (.A1(_315_),
    .A2(_409_),
    .B1(_302_),
    .Y(_410_));
 sky130_fd_sc_hd__a211o_1 _849_ (.A1(net39),
    .A2(_114_),
    .B1(_410_),
    .C1(_100_),
    .X(_080_));
 sky130_fd_sc_hd__ha_1 _850_ (.A(_411_),
    .B(_412_),
    .COUT(_413_),
    .SUM(_414_));
 sky130_fd_sc_hd__ha_1 _851_ (.A(_415_),
    .B(_416_),
    .COUT(_417_),
    .SUM(_418_));
 sky130_fd_sc_hd__ha_1 _852_ (.A(_419_),
    .B(_420_),
    .COUT(_421_),
    .SUM(_422_));
 sky130_fd_sc_hd__ha_1 _853_ (.A(_419_),
    .B(_420_),
    .COUT(_423_),
    .SUM(_424_));
 sky130_fd_sc_hd__ha_1 _854_ (.A(\uart_rx_inst.bit_cnt[0] ),
    .B(_420_),
    .COUT(_425_),
    .SUM(_426_));
 sky130_fd_sc_hd__ha_1 _855_ (.A(_427_),
    .B(_428_),
    .COUT(_429_),
    .SUM(_430_));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.bit_cnt[0]$_SDFFE_PP0P_  (.D(_011_),
    .Q(\uart_rx_inst.bit_cnt[0] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.bit_cnt[1]$_SDFFE_PP0P_  (.D(_012_),
    .Q(\uart_rx_inst.bit_cnt[1] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.bit_cnt[2]$_SDFFE_PP0P_  (.D(_013_),
    .Q(\uart_rx_inst.bit_cnt[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.bit_cnt[3]$_SDFFE_PP0P_  (.D(_014_),
    .Q(\uart_rx_inst.bit_cnt[3] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.busy_reg$_SDFFE_PP0P_  (.D(_015_),
    .Q(net34),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[0]$_SDFFCE_PP0P_  (.D(_016_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[1]$_SDFFCE_PP0P_  (.D(_017_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[2]$_SDFFCE_PP0P_  (.D(_018_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[2] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[3]$_SDFFCE_PP0P_  (.D(_019_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[3] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[4]$_SDFFCE_PP0P_  (.D(_020_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[4] ),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[5]$_SDFFCE_PP0P_  (.D(_021_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[5] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[6]$_SDFFCE_PP0P_  (.D(_022_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[6] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_rx_inst.data_reg[7]$_SDFFCE_PP0P_  (.D(_023_),
    .DE(_001_),
    .Q(\uart_rx_inst.data_reg[7] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.frame_error_reg$_SDFF_PP0_  (.D(_024_),
    .Q(net35),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[0]$_SDFFE_PP0P_  (.D(_025_),
    .Q(net25),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[1]$_SDFFE_PP0P_  (.D(_026_),
    .Q(net26),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[2]$_SDFFE_PP0P_  (.D(_027_),
    .Q(net27),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[3]$_SDFFE_PP0P_  (.D(_028_),
    .Q(net28),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[4]$_SDFFE_PP0P_  (.D(_029_),
    .Q(net29),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[5]$_SDFFE_PP0P_  (.D(_030_),
    .Q(net30),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[6]$_SDFFE_PP0P_  (.D(_031_),
    .Q(net31),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tdata_reg[7]$_SDFFE_PP0P_  (.D(_032_),
    .Q(net32),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.m_axis_tvalid_reg$_SDFF_PP0_  (.D(_033_),
    .Q(net33),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.overrun_error_reg$_SDFF_PP0_  (.D(_034_),
    .Q(net36),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[0]$_SDFFE_PP0P_  (.D(_035_),
    .Q(\uart_rx_inst.prescale_reg[0] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[10]$_SDFFE_PP0P_  (.D(_036_),
    .Q(\uart_rx_inst.prescale_reg[10] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \uart_rx_inst.prescale_reg[11]$_SDFFE_PP0P_  (.D(_037_),
    .Q(\uart_rx_inst.prescale_reg[11] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[12]$_SDFFE_PP0P_  (.D(_038_),
    .Q(\uart_rx_inst.prescale_reg[12] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \uart_rx_inst.prescale_reg[13]$_SDFFE_PP0P_  (.D(_039_),
    .Q(\uart_rx_inst.prescale_reg[13] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[14]$_SDFFE_PP0P_  (.D(_040_),
    .Q(\uart_rx_inst.prescale_reg[14] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[15]$_SDFFE_PP0P_  (.D(_041_),
    .Q(\uart_rx_inst.prescale_reg[15] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[16]$_SDFFE_PP0P_  (.D(_042_),
    .Q(\uart_rx_inst.prescale_reg[16] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[17]$_SDFFE_PP0P_  (.D(_043_),
    .Q(\uart_rx_inst.prescale_reg[17] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[18]$_SDFFE_PP0P_  (.D(_044_),
    .Q(\uart_rx_inst.prescale_reg[18] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[1]$_SDFFE_PP0P_  (.D(_045_),
    .Q(\uart_rx_inst.prescale_reg[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[2]$_SDFFE_PP0P_  (.D(_046_),
    .Q(\uart_rx_inst.prescale_reg[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[3]$_SDFFE_PP0P_  (.D(_047_),
    .Q(\uart_rx_inst.prescale_reg[3] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[4]$_SDFFE_PP0P_  (.D(_048_),
    .Q(\uart_rx_inst.prescale_reg[4] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[5]$_SDFFE_PP0P_  (.D(_049_),
    .Q(\uart_rx_inst.prescale_reg[5] ),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[6]$_SDFFE_PP0P_  (.D(_050_),
    .Q(\uart_rx_inst.prescale_reg[6] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[7]$_SDFFE_PP0P_  (.D(_051_),
    .Q(\uart_rx_inst.prescale_reg[7] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[8]$_SDFFE_PP0P_  (.D(_052_),
    .Q(\uart_rx_inst.prescale_reg[8] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.prescale_reg[9]$_SDFFE_PP0P_  (.D(_053_),
    .Q(\uart_rx_inst.prescale_reg[9] ),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_rx_inst.rxd_reg$_SDFF_PP1_  (.D(_054_),
    .Q(\uart_rx_inst.rxd_reg ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.bit_cnt[0]$_SDFFE_PP0P_  (.D(_055_),
    .Q(\uart_tx_inst.bit_cnt[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \uart_tx_inst.bit_cnt[1]$_SDFFE_PP0P_  (.D(_056_),
    .Q(\uart_tx_inst.bit_cnt[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \uart_tx_inst.bit_cnt[2]$_SDFFE_PP0P_  (.D(_057_),
    .Q(\uart_tx_inst.bit_cnt[2] ),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfxtp_2 \uart_tx_inst.bit_cnt[3]$_SDFFE_PP0P_  (.D(_058_),
    .Q(\uart_tx_inst.bit_cnt[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.busy_reg$_SDFFE_PP0P_  (.D(_059_),
    .Q(net38),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[0]$_DFFE_PP_  (.D(_003_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[1]$_DFFE_PP_  (.D(_004_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[2]$_DFFE_PP_  (.D(_005_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[3]$_DFFE_PP_  (.D(_006_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[3] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[4]$_DFFE_PP_  (.D(_007_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[4] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[5]$_DFFE_PP_  (.D(_008_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[5] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[6]$_DFFE_PP_  (.D(_009_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[6] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[7]$_DFFE_PP_  (.D(_010_),
    .DE(net45),
    .Q(\uart_tx_inst.data_reg[7] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \uart_tx_inst.data_reg[8]$_DFFE_PP_  (.D(_002_),
    .DE(_000_),
    .Q(\uart_tx_inst.data_reg[8] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[0]$_SDFFE_PP0P_  (.D(_060_),
    .Q(\uart_tx_inst.prescale_reg[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[10]$_SDFFE_PP0P_  (.D(_061_),
    .Q(\uart_tx_inst.prescale_reg[10] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[11]$_SDFFE_PP0P_  (.D(_062_),
    .Q(\uart_tx_inst.prescale_reg[11] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[12]$_SDFFE_PP0P_  (.D(_063_),
    .Q(\uart_tx_inst.prescale_reg[12] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[13]$_SDFFE_PP0P_  (.D(_064_),
    .Q(\uart_tx_inst.prescale_reg[13] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[14]$_SDFFE_PP0P_  (.D(_065_),
    .Q(\uart_tx_inst.prescale_reg[14] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[15]$_SDFFE_PP0P_  (.D(_066_),
    .Q(\uart_tx_inst.prescale_reg[15] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[16]$_SDFFE_PP0P_  (.D(_067_),
    .Q(\uart_tx_inst.prescale_reg[16] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[17]$_SDFFE_PP0P_  (.D(_068_),
    .Q(\uart_tx_inst.prescale_reg[17] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[18]$_SDFFE_PP0P_  (.D(_069_),
    .Q(\uart_tx_inst.prescale_reg[18] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[1]$_SDFFE_PP0P_  (.D(_070_),
    .Q(\uart_tx_inst.prescale_reg[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[2]$_SDFFE_PP0P_  (.D(_071_),
    .Q(\uart_tx_inst.prescale_reg[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[3]$_SDFFE_PP0P_  (.D(_072_),
    .Q(\uart_tx_inst.prescale_reg[3] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[4]$_SDFFE_PP0P_  (.D(_073_),
    .Q(\uart_tx_inst.prescale_reg[4] ),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[5]$_SDFFE_PP0P_  (.D(_074_),
    .Q(\uart_tx_inst.prescale_reg[5] ),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[6]$_SDFFE_PP0P_  (.D(_075_),
    .Q(\uart_tx_inst.prescale_reg[6] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[7]$_SDFFE_PP0P_  (.D(_076_),
    .Q(\uart_tx_inst.prescale_reg[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[8]$_SDFFE_PP0P_  (.D(_077_),
    .Q(\uart_tx_inst.prescale_reg[8] ),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.prescale_reg[9]$_SDFFE_PP0P_  (.D(_078_),
    .Q(\uart_tx_inst.prescale_reg[9] ),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.s_axis_tready_reg$_SDFFE_PP0P_  (.D(_079_),
    .Q(net37),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \uart_tx_inst.txd_reg$_SDFFE_PP1P_  (.D(_080_),
    .Q(net39),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 clone2 (.A(_095_),
    .X(net2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_139 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(m_axis_tready),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(prescale[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(prescale[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(prescale[12]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(prescale[13]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(prescale[14]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(prescale[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(prescale[1]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input9 (.A(prescale[2]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input10 (.A(prescale[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(prescale[8]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(prescale[9]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(rst),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(rxd),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(s_axis_tdata[0]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(s_axis_tdata[1]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(s_axis_tdata[2]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(s_axis_tdata[3]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(s_axis_tdata[4]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(s_axis_tdata[5]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(s_axis_tdata[6]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(s_axis_tdata[7]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(s_axis_tvalid),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(m_axis_tdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(m_axis_tdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(m_axis_tdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(m_axis_tdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(m_axis_tdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(m_axis_tdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(m_axis_tdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(m_axis_tdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(m_axis_tvalid));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(rx_busy));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(rx_frame_error));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(rx_overrun_error));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(s_axis_tready));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(tx_busy));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(txd));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_089_),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(\uart_rx_inst.prescale_reg[13] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net49),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net49),
    .X(net44));
 sky130_fd_sc_hd__buf_6 rebuffer6 (.A(_000_),
    .X(net45));
 sky130_fd_sc_hd__buf_2 clone7 (.A(_134_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(_134_),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(_176_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(\uart_rx_inst.prescale_reg[11] ),
    .X(net49));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_7 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_227 ();
endmodule
