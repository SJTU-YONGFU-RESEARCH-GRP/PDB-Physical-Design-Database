module configurable_carry_skip_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sky130_fd_sc_hd__inv_1 _225_ (.A(net65),
    .Y(_053_));
 sky130_fd_sc_hd__inv_1 _226_ (.A(net25),
    .Y(_030_));
 sky130_fd_sc_hd__inv_1 _227_ (.A(net57),
    .Y(_031_));
 sky130_fd_sc_hd__nand4_2 _228_ (.A(_102_),
    .B(_106_),
    .C(_110_),
    .D(_114_),
    .Y(_000_));
 sky130_fd_sc_hd__mux2i_4 _229_ (.A0(net65),
    .A1(_035_),
    .S(_000_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _230_ (.A(_001_),
    .Y(_037_));
 sky130_fd_sc_hd__and4_1 _231_ (.A(_118_),
    .B(_122_),
    .C(_126_),
    .D(_130_),
    .X(_002_));
 sky130_fd_sc_hd__nor2_1 _232_ (.A(_044_),
    .B(_002_),
    .Y(_003_));
 sky130_fd_sc_hd__a21oi_1 _233_ (.A1(_001_),
    .A2(_002_),
    .B1(_003_),
    .Y(_046_));
 sky130_fd_sc_hd__nand4_1 _234_ (.A(_134_),
    .B(_138_),
    .C(_142_),
    .D(_146_),
    .Y(_004_));
 sky130_fd_sc_hd__a211oi_2 _235_ (.A1(_001_),
    .A2(_002_),
    .B1(_003_),
    .C1(_004_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _236_ (.A(_057_),
    .B(_004_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2b_1 _237_ (.A_N(_005_),
    .B(_006_),
    .Y(_059_));
 sky130_fd_sc_hd__and4_1 _238_ (.A(_150_),
    .B(_154_),
    .C(_158_),
    .D(_162_),
    .X(_007_));
 sky130_fd_sc_hd__nand2_1 _239_ (.A(_006_),
    .B(_007_),
    .Y(_008_));
 sky130_fd_sc_hd__o22a_1 _240_ (.A1(_066_),
    .A2(_007_),
    .B1(_008_),
    .B2(_005_),
    .X(_068_));
 sky130_fd_sc_hd__inv_1 _241_ (.A(_054_),
    .Y(_077_));
 sky130_fd_sc_hd__nand4_2 _242_ (.A(_166_),
    .B(_170_),
    .C(_174_),
    .D(_178_),
    .Y(_009_));
 sky130_fd_sc_hd__mux2_1 _243_ (.A0(_068_),
    .A1(_075_),
    .S(_009_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_1 _244_ (.A(_066_),
    .B(_007_),
    .Y(_010_));
 sky130_fd_sc_hd__nand4_1 _245_ (.A(_182_),
    .B(_186_),
    .C(_190_),
    .D(_194_),
    .Y(_011_));
 sky130_fd_sc_hd__nor3_1 _246_ (.A(_010_),
    .B(_009_),
    .C(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__o21ai_1 _247_ (.A1(_005_),
    .A2(_008_),
    .B1(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _248_ (.A(_075_),
    .B(_009_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(_086_),
    .B(_011_),
    .Y(_015_));
 sky130_fd_sc_hd__o21ai_1 _250_ (.A1(_014_),
    .A2(_011_),
    .B1(_015_),
    .Y(_016_));
 sky130_fd_sc_hd__inv_1 _251_ (.A(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__nand2_1 _252_ (.A(_013_),
    .B(_017_),
    .Y(_088_));
 sky130_fd_sc_hd__nand4_1 _253_ (.A(_198_),
    .B(_202_),
    .C(_206_),
    .D(_210_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _254_ (.A(_016_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__nor2b_1 _255_ (.A(_095_),
    .B_N(_018_),
    .Y(_020_));
 sky130_fd_sc_hd__a21oi_1 _256_ (.A1(_013_),
    .A2(_019_),
    .B1(_020_),
    .Y(_097_));
 sky130_fd_sc_hd__inv_1 _257_ (.A(_026_),
    .Y(net89));
 sky130_fd_sc_hd__inv_1 _258_ (.A(_029_),
    .Y(net90));
 sky130_fd_sc_hd__inv_1 _259_ (.A(_034_),
    .Y(net91));
 sky130_fd_sc_hd__inv_1 _260_ (.A(_036_),
    .Y(net92));
 sky130_fd_sc_hd__inv_1 _261_ (.A(_039_),
    .Y(net93));
 sky130_fd_sc_hd__inv_1 _262_ (.A(_041_),
    .Y(net94));
 sky130_fd_sc_hd__inv_1 _263_ (.A(_043_),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _264_ (.A(_045_),
    .Y(net96));
 sky130_fd_sc_hd__inv_1 _265_ (.A(_048_),
    .Y(net97));
 sky130_fd_sc_hd__inv_1 _266_ (.A(_050_),
    .Y(net98));
 sky130_fd_sc_hd__inv_1 _267_ (.A(_056_),
    .Y(net68));
 sky130_fd_sc_hd__inv_1 _268_ (.A(_058_),
    .Y(net69));
 sky130_fd_sc_hd__inv_1 _269_ (.A(_061_),
    .Y(net70));
 sky130_fd_sc_hd__inv_1 _270_ (.A(_063_),
    .Y(net71));
 sky130_fd_sc_hd__inv_1 _271_ (.A(_065_),
    .Y(net72));
 sky130_fd_sc_hd__inv_1 _272_ (.A(_067_),
    .Y(net73));
 sky130_fd_sc_hd__inv_1 _273_ (.A(_070_),
    .Y(net74));
 sky130_fd_sc_hd__inv_1 _274_ (.A(_072_),
    .Y(net75));
 sky130_fd_sc_hd__inv_1 _275_ (.A(_074_),
    .Y(net76));
 sky130_fd_sc_hd__inv_1 _276_ (.A(_076_),
    .Y(net77));
 sky130_fd_sc_hd__inv_1 _277_ (.A(_078_),
    .Y(net78));
 sky130_fd_sc_hd__inv_1 _278_ (.A(_081_),
    .Y(net79));
 sky130_fd_sc_hd__inv_1 _279_ (.A(_083_),
    .Y(net80));
 sky130_fd_sc_hd__inv_1 _280_ (.A(_085_),
    .Y(net81));
 sky130_fd_sc_hd__inv_1 _281_ (.A(_087_),
    .Y(net82));
 sky130_fd_sc_hd__inv_1 _282_ (.A(_090_),
    .Y(net83));
 sky130_fd_sc_hd__inv_1 _283_ (.A(_092_),
    .Y(net84));
 sky130_fd_sc_hd__inv_1 _284_ (.A(_094_),
    .Y(net85));
 sky130_fd_sc_hd__inv_1 _285_ (.A(_096_),
    .Y(net86));
 sky130_fd_sc_hd__inv_1 _286_ (.A(_099_),
    .Y(net87));
 sky130_fd_sc_hd__inv_1 _287_ (.A(_100_),
    .Y(net88));
 sky130_fd_sc_hd__inv_1 _288_ (.A(_028_),
    .Y(_032_));
 sky130_fd_sc_hd__inv_1 _289_ (.A(net1),
    .Y(_051_));
 sky130_fd_sc_hd__inv_1 _290_ (.A(net12),
    .Y(_103_));
 sky130_fd_sc_hd__inv_1 _291_ (.A(net23),
    .Y(_107_));
 sky130_fd_sc_hd__inv_1 _292_ (.A(net26),
    .Y(_111_));
 sky130_fd_sc_hd__inv_1 _293_ (.A(net27),
    .Y(_115_));
 sky130_fd_sc_hd__inv_1 _294_ (.A(net28),
    .Y(_119_));
 sky130_fd_sc_hd__inv_1 _295_ (.A(net29),
    .Y(_123_));
 sky130_fd_sc_hd__inv_1 _296_ (.A(net30),
    .Y(_127_));
 sky130_fd_sc_hd__inv_1 _297_ (.A(net31),
    .Y(_131_));
 sky130_fd_sc_hd__inv_1 _298_ (.A(net32),
    .Y(_135_));
 sky130_fd_sc_hd__inv_1 _299_ (.A(net2),
    .Y(_139_));
 sky130_fd_sc_hd__inv_1 _300_ (.A(net3),
    .Y(_143_));
 sky130_fd_sc_hd__inv_1 _301_ (.A(net4),
    .Y(_147_));
 sky130_fd_sc_hd__inv_1 _302_ (.A(net5),
    .Y(_151_));
 sky130_fd_sc_hd__inv_1 _303_ (.A(net6),
    .Y(_155_));
 sky130_fd_sc_hd__inv_1 _304_ (.A(net7),
    .Y(_159_));
 sky130_fd_sc_hd__inv_1 _305_ (.A(net8),
    .Y(_163_));
 sky130_fd_sc_hd__inv_1 _306_ (.A(net9),
    .Y(_167_));
 sky130_fd_sc_hd__inv_1 _307_ (.A(net10),
    .Y(_171_));
 sky130_fd_sc_hd__inv_1 _308_ (.A(net11),
    .Y(_175_));
 sky130_fd_sc_hd__inv_1 _309_ (.A(net13),
    .Y(_179_));
 sky130_fd_sc_hd__inv_1 _310_ (.A(net14),
    .Y(_183_));
 sky130_fd_sc_hd__inv_1 _311_ (.A(net15),
    .Y(_187_));
 sky130_fd_sc_hd__inv_1 _312_ (.A(net16),
    .Y(_191_));
 sky130_fd_sc_hd__inv_1 _313_ (.A(net17),
    .Y(_195_));
 sky130_fd_sc_hd__inv_1 _314_ (.A(net18),
    .Y(_199_));
 sky130_fd_sc_hd__inv_1 _315_ (.A(net19),
    .Y(_203_));
 sky130_fd_sc_hd__inv_1 _316_ (.A(net20),
    .Y(_207_));
 sky130_fd_sc_hd__inv_1 _317_ (.A(net21),
    .Y(_211_));
 sky130_fd_sc_hd__inv_1 _318_ (.A(net22),
    .Y(_215_));
 sky130_fd_sc_hd__inv_1 _319_ (.A(net24),
    .Y(_219_));
 sky130_fd_sc_hd__inv_1 _320_ (.A(net33),
    .Y(_052_));
 sky130_fd_sc_hd__inv_1 _321_ (.A(net44),
    .Y(_104_));
 sky130_fd_sc_hd__inv_1 _322_ (.A(net55),
    .Y(_108_));
 sky130_fd_sc_hd__inv_1 _323_ (.A(net58),
    .Y(_112_));
 sky130_fd_sc_hd__inv_1 _324_ (.A(net59),
    .Y(_116_));
 sky130_fd_sc_hd__inv_1 _325_ (.A(net60),
    .Y(_120_));
 sky130_fd_sc_hd__inv_1 _326_ (.A(net61),
    .Y(_124_));
 sky130_fd_sc_hd__inv_1 _327_ (.A(net62),
    .Y(_128_));
 sky130_fd_sc_hd__inv_1 _328_ (.A(net63),
    .Y(_132_));
 sky130_fd_sc_hd__inv_1 _329_ (.A(net64),
    .Y(_136_));
 sky130_fd_sc_hd__inv_1 _330_ (.A(net34),
    .Y(_140_));
 sky130_fd_sc_hd__inv_1 _331_ (.A(net35),
    .Y(_144_));
 sky130_fd_sc_hd__inv_1 _332_ (.A(net36),
    .Y(_148_));
 sky130_fd_sc_hd__inv_1 _333_ (.A(net37),
    .Y(_152_));
 sky130_fd_sc_hd__inv_1 _334_ (.A(net38),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _335_ (.A(net39),
    .Y(_160_));
 sky130_fd_sc_hd__inv_1 _336_ (.A(net40),
    .Y(_164_));
 sky130_fd_sc_hd__inv_1 _337_ (.A(net41),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _338_ (.A(net42),
    .Y(_172_));
 sky130_fd_sc_hd__inv_1 _339_ (.A(net43),
    .Y(_176_));
 sky130_fd_sc_hd__inv_1 _340_ (.A(net45),
    .Y(_180_));
 sky130_fd_sc_hd__inv_1 _341_ (.A(net46),
    .Y(_184_));
 sky130_fd_sc_hd__inv_1 _342_ (.A(net47),
    .Y(_188_));
 sky130_fd_sc_hd__inv_1 _343_ (.A(net48),
    .Y(_192_));
 sky130_fd_sc_hd__inv_1 _344_ (.A(net49),
    .Y(_196_));
 sky130_fd_sc_hd__inv_1 _345_ (.A(net50),
    .Y(_200_));
 sky130_fd_sc_hd__inv_1 _346_ (.A(net51),
    .Y(_204_));
 sky130_fd_sc_hd__inv_1 _347_ (.A(net52),
    .Y(_208_));
 sky130_fd_sc_hd__inv_1 _348_ (.A(net53),
    .Y(_212_));
 sky130_fd_sc_hd__inv_1 _349_ (.A(net54),
    .Y(_216_));
 sky130_fd_sc_hd__inv_1 _350_ (.A(net56),
    .Y(_220_));
 sky130_fd_sc_hd__nand4_1 _351_ (.A(_214_),
    .B(_218_),
    .C(_222_),
    .D(_224_),
    .Y(_021_));
 sky130_fd_sc_hd__nor3_1 _352_ (.A(_016_),
    .B(_018_),
    .C(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(_020_),
    .A1(_033_),
    .S(_021_),
    .X(_023_));
 sky130_fd_sc_hd__a21oi_1 _354_ (.A1(_013_),
    .A2(_022_),
    .B1(_023_),
    .Y(net66));
 sky130_fd_sc_hd__fa_1 _355_ (.A(net23),
    .B(net55),
    .CIN(_024_),
    .COUT(_025_),
    .SUM(_026_));
 sky130_fd_sc_hd__fa_1 _356_ (.A(net24),
    .B(net56),
    .CIN(_027_),
    .COUT(_028_),
    .SUM(_029_));
 sky130_fd_sc_hd__fa_1 _357_ (.A(_030_),
    .B(_031_),
    .CIN(_032_),
    .COUT(_033_),
    .SUM(_034_));
 sky130_fd_sc_hd__fa_1 _358_ (.A(net26),
    .B(net58),
    .CIN(_025_),
    .COUT(_035_),
    .SUM(_036_));
 sky130_fd_sc_hd__fa_1 _359_ (.A(net27),
    .B(net59),
    .CIN(_037_),
    .COUT(_038_),
    .SUM(_039_));
 sky130_fd_sc_hd__fa_1 _360_ (.A(net28),
    .B(net60),
    .CIN(_038_),
    .COUT(_040_),
    .SUM(_041_));
 sky130_fd_sc_hd__fa_1 _361_ (.A(net29),
    .B(net61),
    .CIN(_040_),
    .COUT(_042_),
    .SUM(_043_));
 sky130_fd_sc_hd__fa_1 _362_ (.A(net30),
    .B(net62),
    .CIN(_042_),
    .COUT(_044_),
    .SUM(_045_));
 sky130_fd_sc_hd__fa_1 _363_ (.A(net31),
    .B(net63),
    .CIN(_046_),
    .COUT(_047_),
    .SUM(_048_));
 sky130_fd_sc_hd__fa_1 _364_ (.A(net32),
    .B(net64),
    .CIN(_047_),
    .COUT(_049_),
    .SUM(_050_));
 sky130_fd_sc_hd__fa_1 _365_ (.A(_051_),
    .B(_052_),
    .CIN(_053_),
    .COUT(_054_),
    .SUM(net67));
 sky130_fd_sc_hd__fa_1 _366_ (.A(net2),
    .B(net34),
    .CIN(_049_),
    .COUT(_055_),
    .SUM(_056_));
 sky130_fd_sc_hd__fa_1 _367_ (.A(net3),
    .B(net35),
    .CIN(_055_),
    .COUT(_057_),
    .SUM(_058_));
 sky130_fd_sc_hd__fa_1 _368_ (.A(net4),
    .B(net36),
    .CIN(_059_),
    .COUT(_060_),
    .SUM(_061_));
 sky130_fd_sc_hd__fa_1 _369_ (.A(net5),
    .B(net37),
    .CIN(_060_),
    .COUT(_062_),
    .SUM(_063_));
 sky130_fd_sc_hd__fa_1 _370_ (.A(net6),
    .B(net38),
    .CIN(_062_),
    .COUT(_064_),
    .SUM(_065_));
 sky130_fd_sc_hd__fa_1 _371_ (.A(net7),
    .B(net39),
    .CIN(_064_),
    .COUT(_066_),
    .SUM(_067_));
 sky130_fd_sc_hd__fa_1 _372_ (.A(net8),
    .B(net40),
    .CIN(_068_),
    .COUT(_069_),
    .SUM(_070_));
 sky130_fd_sc_hd__fa_1 _373_ (.A(net9),
    .B(net41),
    .CIN(_069_),
    .COUT(_071_),
    .SUM(_072_));
 sky130_fd_sc_hd__fa_1 _374_ (.A(net10),
    .B(net42),
    .CIN(_071_),
    .COUT(_073_),
    .SUM(_074_));
 sky130_fd_sc_hd__fa_1 _375_ (.A(net11),
    .B(net43),
    .CIN(_073_),
    .COUT(_075_),
    .SUM(_076_));
 sky130_fd_sc_hd__fa_1 _376_ (.A(net12),
    .B(net44),
    .CIN(_077_),
    .COUT(_024_),
    .SUM(_078_));
 sky130_fd_sc_hd__fa_1 _377_ (.A(net13),
    .B(net45),
    .CIN(_079_),
    .COUT(_080_),
    .SUM(_081_));
 sky130_fd_sc_hd__fa_1 _378_ (.A(net14),
    .B(net46),
    .CIN(_080_),
    .COUT(_082_),
    .SUM(_083_));
 sky130_fd_sc_hd__fa_1 _379_ (.A(net15),
    .B(net47),
    .CIN(_082_),
    .COUT(_084_),
    .SUM(_085_));
 sky130_fd_sc_hd__fa_1 _380_ (.A(net16),
    .B(net48),
    .CIN(_084_),
    .COUT(_086_),
    .SUM(_087_));
 sky130_fd_sc_hd__fa_1 _381_ (.A(net17),
    .B(net49),
    .CIN(_088_),
    .COUT(_089_),
    .SUM(_090_));
 sky130_fd_sc_hd__fa_1 _382_ (.A(net18),
    .B(net50),
    .CIN(_089_),
    .COUT(_091_),
    .SUM(_092_));
 sky130_fd_sc_hd__fa_1 _383_ (.A(net19),
    .B(net51),
    .CIN(_091_),
    .COUT(_093_),
    .SUM(_094_));
 sky130_fd_sc_hd__fa_1 _384_ (.A(net20),
    .B(net52),
    .CIN(_093_),
    .COUT(_095_),
    .SUM(_096_));
 sky130_fd_sc_hd__fa_1 _385_ (.A(net21),
    .B(net53),
    .CIN(_097_),
    .COUT(_098_),
    .SUM(_099_));
 sky130_fd_sc_hd__fa_1 _386_ (.A(net22),
    .B(net54),
    .CIN(_098_),
    .COUT(_027_),
    .SUM(_100_));
 sky130_fd_sc_hd__ha_1 _387_ (.A(_051_),
    .B(_052_),
    .COUT(_101_),
    .SUM(_102_));
 sky130_fd_sc_hd__ha_1 _388_ (.A(_103_),
    .B(_104_),
    .COUT(_105_),
    .SUM(_106_));
 sky130_fd_sc_hd__ha_1 _389_ (.A(_107_),
    .B(_108_),
    .COUT(_109_),
    .SUM(_110_));
 sky130_fd_sc_hd__ha_1 _390_ (.A(_111_),
    .B(_112_),
    .COUT(_113_),
    .SUM(_114_));
 sky130_fd_sc_hd__ha_1 _391_ (.A(_115_),
    .B(_116_),
    .COUT(_117_),
    .SUM(_118_));
 sky130_fd_sc_hd__ha_1 _392_ (.A(_119_),
    .B(_120_),
    .COUT(_121_),
    .SUM(_122_));
 sky130_fd_sc_hd__ha_1 _393_ (.A(_123_),
    .B(_124_),
    .COUT(_125_),
    .SUM(_126_));
 sky130_fd_sc_hd__ha_1 _394_ (.A(_127_),
    .B(_128_),
    .COUT(_129_),
    .SUM(_130_));
 sky130_fd_sc_hd__ha_1 _395_ (.A(_131_),
    .B(_132_),
    .COUT(_133_),
    .SUM(_134_));
 sky130_fd_sc_hd__ha_1 _396_ (.A(_135_),
    .B(_136_),
    .COUT(_137_),
    .SUM(_138_));
 sky130_fd_sc_hd__ha_1 _397_ (.A(_139_),
    .B(_140_),
    .COUT(_141_),
    .SUM(_142_));
 sky130_fd_sc_hd__ha_1 _398_ (.A(_143_),
    .B(_144_),
    .COUT(_145_),
    .SUM(_146_));
 sky130_fd_sc_hd__ha_1 _399_ (.A(_147_),
    .B(_148_),
    .COUT(_149_),
    .SUM(_150_));
 sky130_fd_sc_hd__ha_1 _400_ (.A(_151_),
    .B(_152_),
    .COUT(_153_),
    .SUM(_154_));
 sky130_fd_sc_hd__ha_1 _401_ (.A(_155_),
    .B(_156_),
    .COUT(_157_),
    .SUM(_158_));
 sky130_fd_sc_hd__ha_1 _402_ (.A(_159_),
    .B(_160_),
    .COUT(_161_),
    .SUM(_162_));
 sky130_fd_sc_hd__ha_1 _403_ (.A(_163_),
    .B(_164_),
    .COUT(_165_),
    .SUM(_166_));
 sky130_fd_sc_hd__ha_1 _404_ (.A(_167_),
    .B(_168_),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__ha_1 _405_ (.A(_171_),
    .B(_172_),
    .COUT(_173_),
    .SUM(_174_));
 sky130_fd_sc_hd__ha_1 _406_ (.A(_175_),
    .B(_176_),
    .COUT(_177_),
    .SUM(_178_));
 sky130_fd_sc_hd__ha_1 _407_ (.A(_179_),
    .B(_180_),
    .COUT(_181_),
    .SUM(_182_));
 sky130_fd_sc_hd__ha_1 _408_ (.A(_183_),
    .B(_184_),
    .COUT(_185_),
    .SUM(_186_));
 sky130_fd_sc_hd__ha_1 _409_ (.A(_187_),
    .B(_188_),
    .COUT(_189_),
    .SUM(_190_));
 sky130_fd_sc_hd__ha_1 _410_ (.A(_191_),
    .B(_192_),
    .COUT(_193_),
    .SUM(_194_));
 sky130_fd_sc_hd__ha_1 _411_ (.A(_195_),
    .B(_196_),
    .COUT(_197_),
    .SUM(_198_));
 sky130_fd_sc_hd__ha_1 _412_ (.A(_199_),
    .B(_200_),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__ha_1 _413_ (.A(_203_),
    .B(_204_),
    .COUT(_205_),
    .SUM(_206_));
 sky130_fd_sc_hd__ha_1 _414_ (.A(_207_),
    .B(_208_),
    .COUT(_209_),
    .SUM(_210_));
 sky130_fd_sc_hd__ha_1 _415_ (.A(_211_),
    .B(_212_),
    .COUT(_213_),
    .SUM(_214_));
 sky130_fd_sc_hd__ha_1 _416_ (.A(_215_),
    .B(_216_),
    .COUT(_217_),
    .SUM(_218_));
 sky130_fd_sc_hd__ha_1 _417_ (.A(_219_),
    .B(_220_),
    .COUT(_221_),
    .SUM(_222_));
 sky130_fd_sc_hd__ha_1 _418_ (.A(_030_),
    .B(_031_),
    .COUT(_223_),
    .SUM(_224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_30 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(sum[9]));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_112 ();
endmodule
