module gray_counter (clk,
    direction,
    enable,
    load,
    rst_n,
    binary_out,
    data_in,
    gray_out);
 input clk;
 input direction;
 input enable;
 input load;
 input rst_n;
 output [3:0] binary_out;
 input [3:0] data_in;
 output [3:0] gray_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net17;

 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _43_ (.A1(net7),
    .A2(net9),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _44_ (.I(net8),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _45_ (.I0(_07_),
    .I1(net2),
    .S(_08_),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _46_ (.I0(net10),
    .I1(_38_),
    .S(net7),
    .Z(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _47_ (.I0(_09_),
    .I1(net3),
    .S(_08_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _48_ (.A1(_42_),
    .A2(_37_),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _49_ (.I0(net11),
    .I1(_10_),
    .S(net7),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _50_ (.I0(_11_),
    .I1(net4),
    .S(_08_),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _51_ (.A1(net9),
    .A2(_42_),
    .A3(_40_),
    .Z(_12_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _52_ (.A1(_42_),
    .A2(_39_),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_4 _53_ (.A1(_41_),
    .A2(_12_),
    .A3(_13_),
    .B(net6),
    .ZN(_14_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _54_ (.A1(net6),
    .A2(_41_),
    .A3(_12_),
    .A4(_13_),
    .Z(_15_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _55_ (.I(net12),
    .ZN(_16_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _56_ (.A1(_14_),
    .A2(_15_),
    .B(_08_),
    .C(_16_),
    .ZN(_17_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _57_ (.I(net7),
    .ZN(_18_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _58_ (.A1(_08_),
    .A2(_18_),
    .ZN(_19_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _59_ (.A1(_16_),
    .A2(_14_),
    .A3(_15_),
    .A4(_19_),
    .Z(_20_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _60_ (.A1(net8),
    .A2(net7),
    .ZN(_21_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _61_ (.A1(_08_),
    .A2(net5),
    .B1(_21_),
    .B2(net12),
    .ZN(_22_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _62_ (.I(_22_),
    .ZN(_23_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _63_ (.A1(_17_),
    .A2(_20_),
    .A3(_23_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _64_ (.A1(net9),
    .A2(_38_),
    .ZN(_24_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _65_ (.I0(net13),
    .I1(_24_),
    .S(net7),
    .Z(_25_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _66_ (.A1(net2),
    .A2(net3),
    .Z(_26_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _67_ (.I0(_25_),
    .I1(_26_),
    .S(_08_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _68_ (.A1(_38_),
    .A2(_10_),
    .Z(_27_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _69_ (.I0(net14),
    .I1(_27_),
    .S(net7),
    .Z(_28_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _70_ (.A1(net3),
    .A2(net4),
    .Z(_29_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _71_ (.I0(_28_),
    .I1(_29_),
    .S(_08_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _72_ (.A1(net12),
    .A2(_42_),
    .A3(_37_),
    .ZN(_30_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _73_ (.A1(_14_),
    .A2(_15_),
    .A3(_19_),
    .A4(_30_),
    .Z(_31_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _74_ (.A1(_08_),
    .A2(_18_),
    .A3(_30_),
    .Z(_32_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _75_ (.A1(_14_),
    .A2(_15_),
    .B(_32_),
    .ZN(_33_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _76_ (.A1(net4),
    .A2(net5),
    .Z(_34_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _77_ (.A1(net15),
    .A2(_21_),
    .B1(_34_),
    .B2(_08_),
    .ZN(_35_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _78_ (.I(_35_),
    .ZN(_36_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _79_ (.A1(_31_),
    .A2(_33_),
    .A3(_36_),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _80_ (.A(net9),
    .B(net10),
    .CI(net6),
    .CO(_37_),
    .S(_38_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _81_ (.A(net10),
    .B(net6),
    .CO(_39_),
    .S(_40_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _82_ (.A(net11),
    .B(net6),
    .CO(_41_),
    .S(_42_));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 _83_ (.I(net12),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \binary_count[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \binary_count[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \binary_count[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net11));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \binary_count[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gray_out[0]$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gray_out[1]$_DFFE_PN0P_  (.D(_05_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \gray_out[2]$_DFFE_PN0P_  (.D(_06_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 hold1 (.I(net17),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_86 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_87 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_88 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_89 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_90 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_91 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_92 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_93 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_94 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_95 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_96 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_98 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_99 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_100 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_101 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_102 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_103 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_104 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(data_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(data_in[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input3 (.I(data_in[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(data_in[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input5 (.I(direction),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input6 (.I(enable),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input7 (.I(load),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output8 (.I(net9),
    .Z(binary_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output9 (.I(net10),
    .Z(binary_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output10 (.I(net11),
    .Z(binary_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(binary_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(gray_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(gray_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(gray_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(gray_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload0 (.I(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_390 ();
endmodule
