module bist_controller (bist_done,
    bist_pass,
    bist_start,
    clk,
    mem_enable,
    mem_write,
    rst_n,
    error_addr,
    error_count,
    mem_addr,
    mem_rdata,
    mem_wdata);
 output bist_done;
 output bist_pass;
 input bist_start;
 input clk;
 output mem_enable;
 output mem_write;
 input rst_n;
 output [4:0] error_addr;
 output [31:0] error_count;
 output [4:0] mem_addr;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire phase_complete;
 wire read_phase;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net113;

 sky130_fd_sc_hd__clkbuf_2 _361_ (.A(net77),
    .X(_051_));
 sky130_fd_sc_hd__nand3_1 _362_ (.A(_051_),
    .B(net76),
    .C(_352_),
    .Y(_355_));
 sky130_fd_sc_hd__inv_1 _363_ (.A(_355_),
    .Y(_358_));
 sky130_fd_sc_hd__inv_1 _364_ (.A(net78),
    .Y(_354_));
 sky130_fd_sc_hd__inv_1 _365_ (.A(net42),
    .Y(_342_));
 sky130_fd_sc_hd__inv_1 _366_ (.A(net74),
    .Y(_348_));
 sky130_fd_sc_hd__inv_1 _367_ (.A(net53),
    .Y(_343_));
 sky130_fd_sc_hd__inv_1 _368_ (.A(net75),
    .Y(_349_));
 sky130_fd_sc_hd__buf_2 _369_ (.A(phase_complete),
    .X(_052_));
 sky130_fd_sc_hd__buf_4 _370_ (.A(\state[2] ),
    .X(_053_));
 sky130_fd_sc_hd__buf_2 _371_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__clkbuf_2 _372_ (.A(\state[0] ),
    .X(_055_));
 sky130_fd_sc_hd__buf_2 _373_ (.A(\state[1] ),
    .X(_056_));
 sky130_fd_sc_hd__a21bo_1 _374_ (.A1(_055_),
    .A2(_056_),
    .B1_N(net112),
    .X(_057_));
 sky130_fd_sc_hd__nand3_1 _375_ (.A(read_phase),
    .B(_055_),
    .C(_056_),
    .Y(_058_));
 sky130_fd_sc_hd__nor4bb_1 _376_ (.A(\state[2] ),
    .B(net112),
    .C_N(_055_),
    .D_N(_056_),
    .Y(_059_));
 sky130_fd_sc_hd__a31oi_1 _377_ (.A1(_054_),
    .A2(_057_),
    .A3(_058_),
    .B1(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__and2_0 _378_ (.A(read_phase),
    .B(_053_),
    .X(_061_));
 sky130_fd_sc_hd__nor3_1 _379_ (.A(_056_),
    .B(_053_),
    .C(net2),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _380_ (.A(_055_),
    .Y(_063_));
 sky130_fd_sc_hd__o21ai_0 _381_ (.A1(_061_),
    .A2(_062_),
    .B1(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__nor2b_1 _382_ (.A(_056_),
    .B_N(_053_),
    .Y(_065_));
 sky130_fd_sc_hd__and3b_1 _383_ (.A_N(_053_),
    .B(_056_),
    .C(_055_),
    .X(_066_));
 sky130_fd_sc_hd__o21ai_0 _384_ (.A1(_065_),
    .A2(_066_),
    .B1(read_phase),
    .Y(_067_));
 sky130_fd_sc_hd__clkbuf_4 _385_ (.A(\state[3] ),
    .X(_068_));
 sky130_fd_sc_hd__clkinv_4 _386_ (.A(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__o2111ai_2 _387_ (.A1(_052_),
    .A2(_060_),
    .B1(_064_),
    .C1(_067_),
    .D1(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2b_1 _388_ (.A(_053_),
    .B_N(net112),
    .Y(_071_));
 sky130_fd_sc_hd__and2_2 _389_ (.A(_055_),
    .B(\state[1] ),
    .X(_072_));
 sky130_fd_sc_hd__o21ai_1 _390_ (.A1(_061_),
    .A2(_071_),
    .B1(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__buf_2 _391_ (.A(_055_),
    .X(_074_));
 sky130_fd_sc_hd__buf_2 _392_ (.A(_056_),
    .X(_075_));
 sky130_fd_sc_hd__nand2_1 _393_ (.A(_074_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__nand3_1 _394_ (.A(_054_),
    .B(net112),
    .C(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a21oi_1 _395_ (.A1(_073_),
    .A2(_077_),
    .B1(_068_),
    .Y(_078_));
 sky130_fd_sc_hd__or2_1 _396_ (.A(_070_),
    .B(_078_),
    .X(_079_));
 sky130_fd_sc_hd__o21ai_4 _397_ (.A1(\state[1] ),
    .A2(\state[2] ),
    .B1(_069_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2_2 _398_ (.A(_074_),
    .B(_056_),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _399_ (.A(_052_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__or3_2 _400_ (.A(_079_),
    .B(_080_),
    .C(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_1 _401_ (.A(_051_),
    .B(net76),
    .Y(_084_));
 sky130_fd_sc_hd__nand2b_2 _402_ (.A_N(_068_),
    .B(_053_),
    .Y(_085_));
 sky130_fd_sc_hd__a311oi_4 _403_ (.A1(_350_),
    .A2(_354_),
    .A3(_084_),
    .B1(_085_),
    .C1(_081_),
    .Y(_086_));
 sky130_fd_sc_hd__or3b_1 _404_ (.A(_074_),
    .B(_075_),
    .C_N(_054_),
    .X(_087_));
 sky130_fd_sc_hd__or3b_1 _405_ (.A(_054_),
    .B(_359_),
    .C_N(_075_),
    .X(_088_));
 sky130_fd_sc_hd__a21oi_2 _406_ (.A1(_087_),
    .A2(_088_),
    .B1(_068_),
    .Y(_089_));
 sky130_fd_sc_hd__o21ai_0 _407_ (.A1(_086_),
    .A2(_089_),
    .B1(_348_),
    .Y(_090_));
 sky130_fd_sc_hd__or2_0 _408_ (.A(_052_),
    .B(_081_),
    .X(_091_));
 sky130_fd_sc_hd__nor2b_1 _409_ (.A(_068_),
    .B_N(_054_),
    .Y(_092_));
 sky130_fd_sc_hd__and3_1 _410_ (.A(_359_),
    .B(_081_),
    .C(_092_),
    .X(_093_));
 sky130_fd_sc_hd__inv_1 _411_ (.A(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__a21oi_1 _412_ (.A1(_091_),
    .A2(_094_),
    .B1(_080_),
    .Y(_095_));
 sky130_fd_sc_hd__o21ai_0 _413_ (.A1(_079_),
    .A2(_095_),
    .B1(net74),
    .Y(_096_));
 sky130_fd_sc_hd__o21ai_0 _414_ (.A1(_083_),
    .A2(_090_),
    .B1(_096_),
    .Y(_000_));
 sky130_fd_sc_hd__o21bai_1 _415_ (.A1(_080_),
    .A2(_091_),
    .B1_N(_079_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _416_ (.A(_093_),
    .B(_086_),
    .Y(_098_));
 sky130_fd_sc_hd__nor2_1 _417_ (.A(_351_),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _418_ (.A1(_351_),
    .A2(_089_),
    .B1(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__o2bb2ai_1 _419_ (.A1_N(net75),
    .A2_N(_097_),
    .B1(_083_),
    .B2(_100_),
    .Y(_001_));
 sky130_fd_sc_hd__a22oi_1 _420_ (.A1(_350_),
    .A2(_086_),
    .B1(_089_),
    .B2(_352_),
    .Y(_101_));
 sky130_fd_sc_hd__nand3b_1 _421_ (.A_N(_352_),
    .B(_089_),
    .C(net76),
    .Y(_102_));
 sky130_fd_sc_hd__o21ai_0 _422_ (.A1(net76),
    .A2(_101_),
    .B1(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__nor2_1 _423_ (.A(_093_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__or3_1 _424_ (.A(_350_),
    .B(_081_),
    .C(_085_),
    .X(_105_));
 sky130_fd_sc_hd__a21oi_1 _425_ (.A1(_091_),
    .A2(_105_),
    .B1(_080_),
    .Y(_106_));
 sky130_fd_sc_hd__o21ai_0 _426_ (.A1(_079_),
    .A2(_106_),
    .B1(net76),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _427_ (.A1(_083_),
    .A2(_104_),
    .B1(_107_),
    .Y(_002_));
 sky130_fd_sc_hd__nand3_1 _428_ (.A(net76),
    .B(net74),
    .C(net75),
    .Y(_108_));
 sky130_fd_sc_hd__xnor2_1 _429_ (.A(_051_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nor3_1 _430_ (.A(net76),
    .B(net74),
    .C(net75),
    .Y(_110_));
 sky130_fd_sc_hd__xor2_1 _431_ (.A(_051_),
    .B(_110_),
    .X(_111_));
 sky130_fd_sc_hd__a22o_1 _432_ (.A1(_089_),
    .A2(_109_),
    .B1(_111_),
    .B2(_086_),
    .X(_112_));
 sky130_fd_sc_hd__nor2_1 _433_ (.A(_093_),
    .B(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__o2bb2ai_1 _434_ (.A1_N(_051_),
    .A2_N(_097_),
    .B1(_113_),
    .B2(_083_),
    .Y(_003_));
 sky130_fd_sc_hd__buf_2 _435_ (.A(_068_),
    .X(_114_));
 sky130_fd_sc_hd__buf_2 _436_ (.A(_054_),
    .X(_115_));
 sky130_fd_sc_hd__inv_1 _437_ (.A(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2_1 _438_ (.A(_356_),
    .B(_087_),
    .Y(_117_));
 sky130_fd_sc_hd__a31oi_1 _439_ (.A1(_075_),
    .A2(_116_),
    .A3(_357_),
    .B1(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__a211oi_1 _440_ (.A1(_350_),
    .A2(_084_),
    .B1(_085_),
    .C1(_081_),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(_082_),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_1 _442_ (.A(_080_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__o21ai_0 _443_ (.A1(_079_),
    .A2(_121_),
    .B1(net78),
    .Y(_122_));
 sky130_fd_sc_hd__o31ai_1 _444_ (.A1(_114_),
    .A2(_083_),
    .A3(_118_),
    .B1(_122_),
    .Y(_004_));
 sky130_fd_sc_hd__nor3_1 _445_ (.A(_074_),
    .B(_075_),
    .C(_115_),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(_114_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(net2),
    .B(_123_),
    .Y(_125_));
 sky130_fd_sc_hd__nand2_1 _448_ (.A(net35),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(_124_),
    .B(_126_),
    .Y(_005_));
 sky130_fd_sc_hd__nor4b_1 _450_ (.A(net60),
    .B(net65),
    .C(net66),
    .D_N(_344_),
    .Y(_127_));
 sky130_fd_sc_hd__nor4_1 _451_ (.A(net51),
    .B(net61),
    .C(net62),
    .D(net63),
    .Y(_128_));
 sky130_fd_sc_hd__clkbuf_2 _452_ (.A(net57),
    .X(_129_));
 sky130_fd_sc_hd__nor4_1 _453_ (.A(net56),
    .B(_129_),
    .C(net58),
    .D(net59),
    .Y(_130_));
 sky130_fd_sc_hd__nor3_1 _454_ (.A(net52),
    .B(net54),
    .C(net55),
    .Y(_131_));
 sky130_fd_sc_hd__nand4_1 _455_ (.A(_127_),
    .B(_128_),
    .C(_130_),
    .D(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__clkbuf_2 _456_ (.A(net72),
    .X(_133_));
 sky130_fd_sc_hd__nor4_1 _457_ (.A(net70),
    .B(net71),
    .C(_133_),
    .D(net73),
    .Y(_134_));
 sky130_fd_sc_hd__buf_2 _458_ (.A(net68),
    .X(_135_));
 sky130_fd_sc_hd__nor4_1 _459_ (.A(net64),
    .B(net67),
    .C(_135_),
    .D(net69),
    .Y(_136_));
 sky130_fd_sc_hd__nor4_1 _460_ (.A(net43),
    .B(net47),
    .C(net48),
    .D(net49),
    .Y(_137_));
 sky130_fd_sc_hd__nor4_1 _461_ (.A(net44),
    .B(net45),
    .C(net46),
    .D(net50),
    .Y(_138_));
 sky130_fd_sc_hd__nand4_1 _462_ (.A(_134_),
    .B(_136_),
    .C(_137_),
    .D(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_0 _463_ (.A1(_114_),
    .A2(net2),
    .B1(_123_),
    .Y(_140_));
 sky130_fd_sc_hd__nand2_1 _464_ (.A(net36),
    .B(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__o31ai_1 _465_ (.A1(_124_),
    .A2(_132_),
    .A3(_139_),
    .B1(_141_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(_063_),
    .B(_092_),
    .Y(_142_));
 sky130_fd_sc_hd__nor4_1 _467_ (.A(net11),
    .B(net15),
    .C(net18),
    .D(net17),
    .Y(_143_));
 sky130_fd_sc_hd__nor4_1 _468_ (.A(net10),
    .B(net13),
    .C(net12),
    .D(net16),
    .Y(_144_));
 sky130_fd_sc_hd__nor4_1 _469_ (.A(net20),
    .B(net23),
    .C(net27),
    .D(net26),
    .Y(_145_));
 sky130_fd_sc_hd__nor4_1 _470_ (.A(net19),
    .B(net22),
    .C(net21),
    .D(net24),
    .Y(_146_));
 sky130_fd_sc_hd__nand4_1 _471_ (.A(_143_),
    .B(_144_),
    .C(_145_),
    .D(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__nor4_1 _472_ (.A(net30),
    .B(net29),
    .C(net32),
    .D(net8),
    .Y(_148_));
 sky130_fd_sc_hd__nor4_1 _473_ (.A(net14),
    .B(net3),
    .C(net28),
    .D(net25),
    .Y(_149_));
 sky130_fd_sc_hd__nor4_1 _474_ (.A(net31),
    .B(net7),
    .C(net6),
    .D(net9),
    .Y(_150_));
 sky130_fd_sc_hd__nor4_1 _475_ (.A(net34),
    .B(net33),
    .C(net5),
    .D(net4),
    .Y(_151_));
 sky130_fd_sc_hd__nand4_1 _476_ (.A(_148_),
    .B(_149_),
    .C(_150_),
    .D(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__o21ai_0 _477_ (.A1(_147_),
    .A2(_152_),
    .B1(read_phase),
    .Y(_153_));
 sky130_fd_sc_hd__o21ai_4 _478_ (.A1(_054_),
    .A2(_072_),
    .B1(_069_),
    .Y(_154_));
 sky130_fd_sc_hd__nand4_1 _479_ (.A(net11),
    .B(net15),
    .C(net18),
    .D(net17),
    .Y(_155_));
 sky130_fd_sc_hd__nand4_1 _480_ (.A(net10),
    .B(net13),
    .C(net12),
    .D(net16),
    .Y(_156_));
 sky130_fd_sc_hd__nand4_1 _481_ (.A(net20),
    .B(net23),
    .C(net27),
    .D(net26),
    .Y(_157_));
 sky130_fd_sc_hd__nand4_1 _482_ (.A(net19),
    .B(net22),
    .C(net21),
    .D(net24),
    .Y(_158_));
 sky130_fd_sc_hd__nor4_1 _483_ (.A(_155_),
    .B(_156_),
    .C(_157_),
    .D(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__nand4_1 _484_ (.A(net30),
    .B(net29),
    .C(net32),
    .D(net8),
    .Y(_160_));
 sky130_fd_sc_hd__nand4_1 _485_ (.A(net14),
    .B(net3),
    .C(net28),
    .D(net25),
    .Y(_161_));
 sky130_fd_sc_hd__nand4_1 _486_ (.A(net31),
    .B(net7),
    .C(net6),
    .D(net9),
    .Y(_162_));
 sky130_fd_sc_hd__nand4_1 _487_ (.A(net34),
    .B(net33),
    .C(net5),
    .D(net4),
    .Y(_163_));
 sky130_fd_sc_hd__nor4_1 _488_ (.A(_160_),
    .B(_161_),
    .C(_162_),
    .D(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__a21boi_2 _489_ (.A1(_159_),
    .A2(_164_),
    .B1_N(read_phase),
    .Y(_165_));
 sky130_fd_sc_hd__nand3b_1 _490_ (.A_N(net112),
    .B(\state[1] ),
    .C(_055_),
    .Y(_166_));
 sky130_fd_sc_hd__nand2b_1 _491_ (.A_N(net112),
    .B(\state[2] ),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _492_ (.A(\state[1] ),
    .B(\state[2] ),
    .Y(_168_));
 sky130_fd_sc_hd__or2_0 _493_ (.A(read_phase),
    .B(_052_),
    .X(_169_));
 sky130_fd_sc_hd__a31oi_1 _494_ (.A1(_166_),
    .A2(_167_),
    .A3(_168_),
    .B1(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__a21oi_1 _495_ (.A1(_063_),
    .A2(\state[2] ),
    .B1(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__nor3_1 _496_ (.A(_068_),
    .B(_165_),
    .C(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__a211o_1 _497_ (.A1(_142_),
    .A2(_153_),
    .B1(_154_),
    .C1(_172_),
    .X(_173_));
 sky130_fd_sc_hd__buf_2 _498_ (.A(_173_),
    .X(_174_));
 sky130_fd_sc_hd__clkbuf_4 _499_ (.A(_174_),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _500_ (.A0(net74),
    .A1(net37),
    .S(_175_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _501_ (.A0(net75),
    .A1(net38),
    .S(_174_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(net76),
    .A1(net39),
    .S(_174_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(_051_),
    .A1(net40),
    .S(_174_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _504_ (.A0(net78),
    .A1(net41),
    .S(_174_),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_4 _505_ (.A(_174_),
    .X(_176_));
 sky130_fd_sc_hd__inv_1 _506_ (.A(_056_),
    .Y(_177_));
 sky130_fd_sc_hd__a21oi_1 _507_ (.A1(_177_),
    .A2(net2),
    .B1(_053_),
    .Y(_178_));
 sky130_fd_sc_hd__o21ai_0 _508_ (.A1(_053_),
    .A2(_072_),
    .B1(read_phase),
    .Y(_179_));
 sky130_fd_sc_hd__o21ai_1 _509_ (.A1(_055_),
    .A2(_178_),
    .B1(_179_),
    .Y(_180_));
 sky130_fd_sc_hd__or4_1 _510_ (.A(_063_),
    .B(_080_),
    .C(_147_),
    .D(_152_),
    .X(_181_));
 sky130_fd_sc_hd__o2111ai_4 _511_ (.A1(_165_),
    .A2(_171_),
    .B1(_180_),
    .C1(_181_),
    .D1(_069_),
    .Y(_182_));
 sky130_fd_sc_hd__buf_2 _512_ (.A(_182_),
    .X(_183_));
 sky130_fd_sc_hd__nand2_1 _513_ (.A(net42),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__o21ai_0 _514_ (.A1(net42),
    .A2(_176_),
    .B1(_184_),
    .Y(_012_));
 sky130_fd_sc_hd__and3_1 _515_ (.A(_346_),
    .B(net64),
    .C(net67),
    .X(_185_));
 sky130_fd_sc_hd__and2_0 _516_ (.A(net70),
    .B(net71),
    .X(_186_));
 sky130_fd_sc_hd__nand4_4 _517_ (.A(_135_),
    .B(net69),
    .C(_185_),
    .D(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(_133_),
    .B(net73),
    .Y(_188_));
 sky130_fd_sc_hd__nand3_1 _519_ (.A(_346_),
    .B(net64),
    .C(net67),
    .Y(_189_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_135_),
    .B(net69),
    .Y(_190_));
 sky130_fd_sc_hd__nor3b_2 _521_ (.A(_189_),
    .B(_190_),
    .C_N(_186_),
    .Y(_191_));
 sky130_fd_sc_hd__clkbuf_4 _522_ (.A(_154_),
    .X(_192_));
 sky130_fd_sc_hd__a31oi_1 _523_ (.A1(_133_),
    .A2(net73),
    .A3(_191_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__o21ai_0 _524_ (.A1(_183_),
    .A2(_193_),
    .B1(net43),
    .Y(_194_));
 sky130_fd_sc_hd__o41ai_1 _525_ (.A1(net43),
    .A2(_175_),
    .A3(_187_),
    .A4(_188_),
    .B1(_194_),
    .Y(_013_));
 sky130_fd_sc_hd__inv_1 _526_ (.A(net71),
    .Y(_195_));
 sky130_fd_sc_hd__nand3_1 _527_ (.A(net64),
    .B(net67),
    .C(_135_),
    .Y(_196_));
 sky130_fd_sc_hd__nand2_1 _528_ (.A(net42),
    .B(net53),
    .Y(_197_));
 sky130_fd_sc_hd__nand2_1 _529_ (.A(net69),
    .B(net70),
    .Y(_198_));
 sky130_fd_sc_hd__or4_1 _530_ (.A(_195_),
    .B(_196_),
    .C(_197_),
    .D(_198_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_2 _531_ (.A(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand3_1 _532_ (.A(_133_),
    .B(net73),
    .C(net43),
    .Y(_201_));
 sky130_fd_sc_hd__clkbuf_4 _533_ (.A(_154_),
    .X(_202_));
 sky130_fd_sc_hd__nor2_1 _534_ (.A(_200_),
    .B(_201_),
    .Y(_203_));
 sky130_fd_sc_hd__nor2_1 _535_ (.A(_202_),
    .B(_203_),
    .Y(_204_));
 sky130_fd_sc_hd__o21ai_0 _536_ (.A1(_183_),
    .A2(_204_),
    .B1(net44),
    .Y(_205_));
 sky130_fd_sc_hd__o41ai_1 _537_ (.A1(net44),
    .A2(_175_),
    .A3(_200_),
    .A4(_201_),
    .B1(_205_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _538_ (.A(net43),
    .B(net44),
    .Y(_206_));
 sky130_fd_sc_hd__nor3_1 _539_ (.A(_187_),
    .B(_188_),
    .C(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__nand2b_1 _540_ (.A_N(net45),
    .B(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__buf_2 _541_ (.A(_182_),
    .X(_209_));
 sky130_fd_sc_hd__nor2_1 _542_ (.A(_192_),
    .B(_207_),
    .Y(_210_));
 sky130_fd_sc_hd__o21ai_0 _543_ (.A1(_209_),
    .A2(_210_),
    .B1(net45),
    .Y(_211_));
 sky130_fd_sc_hd__o21ai_0 _544_ (.A1(_176_),
    .A2(_208_),
    .B1(_211_),
    .Y(_015_));
 sky130_fd_sc_hd__nor3_2 _545_ (.A(_196_),
    .B(_197_),
    .C(_198_),
    .Y(_212_));
 sky130_fd_sc_hd__nand3_1 _546_ (.A(net43),
    .B(net44),
    .C(net45),
    .Y(_213_));
 sky130_fd_sc_hd__nor2_1 _547_ (.A(_188_),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__nand3_1 _548_ (.A(net71),
    .B(_212_),
    .C(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__buf_2 _549_ (.A(_182_),
    .X(_216_));
 sky130_fd_sc_hd__a31oi_1 _550_ (.A1(net71),
    .A2(_212_),
    .A3(_214_),
    .B1(_192_),
    .Y(_217_));
 sky130_fd_sc_hd__o21ai_0 _551_ (.A1(_216_),
    .A2(_217_),
    .B1(net46),
    .Y(_218_));
 sky130_fd_sc_hd__o31ai_1 _552_ (.A1(net46),
    .A2(_176_),
    .A3(_215_),
    .B1(_218_),
    .Y(_016_));
 sky130_fd_sc_hd__nand3_1 _553_ (.A(net46),
    .B(_191_),
    .C(_214_),
    .Y(_219_));
 sky130_fd_sc_hd__a31oi_1 _554_ (.A1(net46),
    .A2(_191_),
    .A3(_214_),
    .B1(_192_),
    .Y(_220_));
 sky130_fd_sc_hd__o21ai_0 _555_ (.A1(_216_),
    .A2(_220_),
    .B1(net47),
    .Y(_221_));
 sky130_fd_sc_hd__o31ai_1 _556_ (.A1(net47),
    .A2(_176_),
    .A3(_219_),
    .B1(_221_),
    .Y(_017_));
 sky130_fd_sc_hd__and2_0 _557_ (.A(net46),
    .B(net47),
    .X(_222_));
 sky130_fd_sc_hd__or3b_1 _558_ (.A(_188_),
    .B(_213_),
    .C_N(_222_),
    .X(_223_));
 sky130_fd_sc_hd__buf_2 _559_ (.A(_223_),
    .X(_224_));
 sky130_fd_sc_hd__nor2_2 _560_ (.A(_200_),
    .B(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__nor2_1 _561_ (.A(_202_),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__o21ai_0 _562_ (.A1(_183_),
    .A2(_226_),
    .B1(net48),
    .Y(_227_));
 sky130_fd_sc_hd__o41ai_1 _563_ (.A1(net48),
    .A2(_175_),
    .A3(_200_),
    .A4(_224_),
    .B1(_227_),
    .Y(_018_));
 sky130_fd_sc_hd__nand4_1 _564_ (.A(net45),
    .B(net48),
    .C(_207_),
    .D(_222_),
    .Y(_228_));
 sky130_fd_sc_hd__clkbuf_4 _565_ (.A(_154_),
    .X(_229_));
 sky130_fd_sc_hd__a41oi_1 _566_ (.A1(net45),
    .A2(net48),
    .A3(_207_),
    .A4(_222_),
    .B1(_229_),
    .Y(_230_));
 sky130_fd_sc_hd__o21ai_0 _567_ (.A1(_216_),
    .A2(_230_),
    .B1(net49),
    .Y(_231_));
 sky130_fd_sc_hd__o31ai_1 _568_ (.A1(net49),
    .A2(_176_),
    .A3(_228_),
    .B1(_231_),
    .Y(_019_));
 sky130_fd_sc_hd__and2_0 _569_ (.A(net48),
    .B(net49),
    .X(_232_));
 sky130_fd_sc_hd__clkbuf_2 _570_ (.A(_232_),
    .X(_233_));
 sky130_fd_sc_hd__nand2_1 _571_ (.A(_225_),
    .B(_233_),
    .Y(_234_));
 sky130_fd_sc_hd__a21oi_1 _572_ (.A1(_225_),
    .A2(_233_),
    .B1(_202_),
    .Y(_235_));
 sky130_fd_sc_hd__o21ai_0 _573_ (.A1(_216_),
    .A2(_235_),
    .B1(net50),
    .Y(_236_));
 sky130_fd_sc_hd__o31ai_1 _574_ (.A1(net50),
    .A2(_176_),
    .A3(_234_),
    .B1(_236_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_2 _575_ (.A(_187_),
    .B(_224_),
    .Y(_237_));
 sky130_fd_sc_hd__nand3_1 _576_ (.A(net50),
    .B(_233_),
    .C(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__a31oi_1 _577_ (.A1(net50),
    .A2(_233_),
    .A3(_237_),
    .B1(_229_),
    .Y(_239_));
 sky130_fd_sc_hd__o21ai_0 _578_ (.A1(_216_),
    .A2(_239_),
    .B1(net51),
    .Y(_240_));
 sky130_fd_sc_hd__o31ai_1 _579_ (.A1(net51),
    .A2(_176_),
    .A3(_238_),
    .B1(_240_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _580_ (.A(net50),
    .B(net51),
    .Y(_241_));
 sky130_fd_sc_hd__a41oi_1 _581_ (.A1(net50),
    .A2(net51),
    .A3(_225_),
    .A4(_233_),
    .B1(_229_),
    .Y(_242_));
 sky130_fd_sc_hd__o21ai_0 _582_ (.A1(_183_),
    .A2(_242_),
    .B1(net52),
    .Y(_243_));
 sky130_fd_sc_hd__o41ai_1 _583_ (.A1(net52),
    .A2(_175_),
    .A3(_234_),
    .A4(_241_),
    .B1(_243_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_1 _584_ (.A(_345_),
    .Y(_244_));
 sky130_fd_sc_hd__nand2_1 _585_ (.A(net53),
    .B(_183_),
    .Y(_245_));
 sky130_fd_sc_hd__o31ai_1 _586_ (.A1(_244_),
    .A2(_202_),
    .A3(_183_),
    .B1(_245_),
    .Y(_023_));
 sky130_fd_sc_hd__buf_2 _587_ (.A(_174_),
    .X(_246_));
 sky130_fd_sc_hd__and3_1 _588_ (.A(net50),
    .B(net51),
    .C(net52),
    .X(_247_));
 sky130_fd_sc_hd__nand3_1 _589_ (.A(_233_),
    .B(_237_),
    .C(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__a31oi_1 _590_ (.A1(_233_),
    .A2(_237_),
    .A3(_247_),
    .B1(_229_),
    .Y(_249_));
 sky130_fd_sc_hd__o21ai_0 _591_ (.A1(_216_),
    .A2(_249_),
    .B1(net54),
    .Y(_250_));
 sky130_fd_sc_hd__o31ai_1 _592_ (.A1(net54),
    .A2(_246_),
    .A3(_248_),
    .B1(_250_),
    .Y(_024_));
 sky130_fd_sc_hd__and3_1 _593_ (.A(net48),
    .B(net49),
    .C(net54),
    .X(_251_));
 sky130_fd_sc_hd__and2_0 _594_ (.A(_247_),
    .B(_251_),
    .X(_252_));
 sky130_fd_sc_hd__nand2_1 _595_ (.A(_225_),
    .B(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__a21oi_1 _596_ (.A1(_225_),
    .A2(_252_),
    .B1(_202_),
    .Y(_254_));
 sky130_fd_sc_hd__o21ai_0 _597_ (.A1(_216_),
    .A2(_254_),
    .B1(net55),
    .Y(_255_));
 sky130_fd_sc_hd__o31ai_1 _598_ (.A1(net55),
    .A2(_246_),
    .A3(_253_),
    .B1(_255_),
    .Y(_025_));
 sky130_fd_sc_hd__nand3_1 _599_ (.A(net55),
    .B(_237_),
    .C(_252_),
    .Y(_256_));
 sky130_fd_sc_hd__a31oi_1 _600_ (.A1(net55),
    .A2(_237_),
    .A3(_252_),
    .B1(_229_),
    .Y(_257_));
 sky130_fd_sc_hd__o21ai_0 _601_ (.A1(_216_),
    .A2(_257_),
    .B1(net56),
    .Y(_258_));
 sky130_fd_sc_hd__o31ai_1 _602_ (.A1(net56),
    .A2(_246_),
    .A3(_256_),
    .B1(_258_),
    .Y(_026_));
 sky130_fd_sc_hd__nand4_4 _603_ (.A(net55),
    .B(net56),
    .C(_247_),
    .D(_251_),
    .Y(_259_));
 sky130_fd_sc_hd__nor3_4 _604_ (.A(_200_),
    .B(_224_),
    .C(_259_),
    .Y(_260_));
 sky130_fd_sc_hd__nand2b_1 _605_ (.A_N(_129_),
    .B(_260_),
    .Y(_261_));
 sky130_fd_sc_hd__nor2_1 _606_ (.A(_192_),
    .B(_260_),
    .Y(_262_));
 sky130_fd_sc_hd__o21ai_0 _607_ (.A1(_182_),
    .A2(_262_),
    .B1(_129_),
    .Y(_263_));
 sky130_fd_sc_hd__o21ai_0 _608_ (.A1(_176_),
    .A2(_261_),
    .B1(_263_),
    .Y(_027_));
 sky130_fd_sc_hd__nor3_4 _609_ (.A(_187_),
    .B(_224_),
    .C(_259_),
    .Y(_264_));
 sky130_fd_sc_hd__nand2_1 _610_ (.A(_129_),
    .B(_264_),
    .Y(_265_));
 sky130_fd_sc_hd__a21oi_1 _611_ (.A1(_129_),
    .A2(_264_),
    .B1(_192_),
    .Y(_266_));
 sky130_fd_sc_hd__o21ai_0 _612_ (.A1(_216_),
    .A2(_266_),
    .B1(net58),
    .Y(_267_));
 sky130_fd_sc_hd__o31ai_1 _613_ (.A1(net58),
    .A2(_246_),
    .A3(_265_),
    .B1(_267_),
    .Y(_028_));
 sky130_fd_sc_hd__nand3_1 _614_ (.A(_129_),
    .B(net58),
    .C(_260_),
    .Y(_268_));
 sky130_fd_sc_hd__a31oi_1 _615_ (.A1(_129_),
    .A2(net58),
    .A3(_260_),
    .B1(_229_),
    .Y(_269_));
 sky130_fd_sc_hd__o21ai_0 _616_ (.A1(_209_),
    .A2(_269_),
    .B1(net59),
    .Y(_270_));
 sky130_fd_sc_hd__o31ai_1 _617_ (.A1(net59),
    .A2(_246_),
    .A3(_268_),
    .B1(_270_),
    .Y(_029_));
 sky130_fd_sc_hd__nand4_1 _618_ (.A(_129_),
    .B(net58),
    .C(net59),
    .D(_264_),
    .Y(_271_));
 sky130_fd_sc_hd__a41oi_1 _619_ (.A1(_129_),
    .A2(net58),
    .A3(net59),
    .A4(_264_),
    .B1(_229_),
    .Y(_272_));
 sky130_fd_sc_hd__o21ai_0 _620_ (.A1(_209_),
    .A2(_272_),
    .B1(net60),
    .Y(_273_));
 sky130_fd_sc_hd__o31ai_1 _621_ (.A1(net60),
    .A2(_246_),
    .A3(_271_),
    .B1(_273_),
    .Y(_030_));
 sky130_fd_sc_hd__and4_1 _622_ (.A(_129_),
    .B(net58),
    .C(net59),
    .D(net60),
    .X(_274_));
 sky130_fd_sc_hd__nand2_1 _623_ (.A(_260_),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__a21oi_1 _624_ (.A1(_260_),
    .A2(_274_),
    .B1(_192_),
    .Y(_276_));
 sky130_fd_sc_hd__o21ai_0 _625_ (.A1(_209_),
    .A2(_276_),
    .B1(net61),
    .Y(_277_));
 sky130_fd_sc_hd__o31ai_1 _626_ (.A1(net61),
    .A2(_246_),
    .A3(_275_),
    .B1(_277_),
    .Y(_031_));
 sky130_fd_sc_hd__nand3_1 _627_ (.A(net61),
    .B(_264_),
    .C(_274_),
    .Y(_278_));
 sky130_fd_sc_hd__a31oi_1 _628_ (.A1(net61),
    .A2(_264_),
    .A3(_274_),
    .B1(_229_),
    .Y(_279_));
 sky130_fd_sc_hd__o21ai_0 _629_ (.A1(_209_),
    .A2(_279_),
    .B1(net62),
    .Y(_280_));
 sky130_fd_sc_hd__o31ai_1 _630_ (.A1(net62),
    .A2(_246_),
    .A3(_278_),
    .B1(_280_),
    .Y(_032_));
 sky130_fd_sc_hd__and3_1 _631_ (.A(net61),
    .B(net62),
    .C(_274_),
    .X(_281_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _632_ (.A(_281_),
    .X(_282_));
 sky130_fd_sc_hd__nand2_1 _633_ (.A(_260_),
    .B(_282_),
    .Y(_283_));
 sky130_fd_sc_hd__a21oi_1 _634_ (.A1(_260_),
    .A2(_282_),
    .B1(_192_),
    .Y(_284_));
 sky130_fd_sc_hd__o21ai_0 _635_ (.A1(_209_),
    .A2(_284_),
    .B1(net63),
    .Y(_285_));
 sky130_fd_sc_hd__o31ai_1 _636_ (.A1(net63),
    .A2(_246_),
    .A3(_283_),
    .B1(_285_),
    .Y(_033_));
 sky130_fd_sc_hd__nand2b_1 _637_ (.A_N(net64),
    .B(_346_),
    .Y(_286_));
 sky130_fd_sc_hd__nor2_1 _638_ (.A(_346_),
    .B(_202_),
    .Y(_287_));
 sky130_fd_sc_hd__o21ai_0 _639_ (.A1(_182_),
    .A2(_287_),
    .B1(net64),
    .Y(_288_));
 sky130_fd_sc_hd__o21ai_0 _640_ (.A1(_176_),
    .A2(_286_),
    .B1(_288_),
    .Y(_034_));
 sky130_fd_sc_hd__nand3_1 _641_ (.A(net63),
    .B(_264_),
    .C(_282_),
    .Y(_289_));
 sky130_fd_sc_hd__a31oi_1 _642_ (.A1(net63),
    .A2(_264_),
    .A3(_282_),
    .B1(_229_),
    .Y(_290_));
 sky130_fd_sc_hd__o21ai_0 _643_ (.A1(_209_),
    .A2(_290_),
    .B1(net65),
    .Y(_291_));
 sky130_fd_sc_hd__o31ai_1 _644_ (.A1(net65),
    .A2(_246_),
    .A3(_289_),
    .B1(_291_),
    .Y(_035_));
 sky130_fd_sc_hd__nand4_1 _645_ (.A(net63),
    .B(net65),
    .C(_260_),
    .D(_282_),
    .Y(_292_));
 sky130_fd_sc_hd__a41oi_1 _646_ (.A1(net63),
    .A2(net65),
    .A3(_260_),
    .A4(_282_),
    .B1(_154_),
    .Y(_293_));
 sky130_fd_sc_hd__o21ai_0 _647_ (.A1(_209_),
    .A2(_293_),
    .B1(net66),
    .Y(_294_));
 sky130_fd_sc_hd__o31ai_1 _648_ (.A1(net66),
    .A2(_175_),
    .A3(_292_),
    .B1(_294_),
    .Y(_036_));
 sky130_fd_sc_hd__nand3_1 _649_ (.A(net42),
    .B(net64),
    .C(net53),
    .Y(_295_));
 sky130_fd_sc_hd__nand2_1 _650_ (.A(net67),
    .B(_295_),
    .Y(_296_));
 sky130_fd_sc_hd__nand2_1 _651_ (.A(net67),
    .B(_183_),
    .Y(_297_));
 sky130_fd_sc_hd__or4_1 _652_ (.A(net67),
    .B(_154_),
    .C(_182_),
    .D(_295_),
    .X(_298_));
 sky130_fd_sc_hd__o211ai_1 _653_ (.A1(_202_),
    .A2(_296_),
    .B1(_297_),
    .C1(_298_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _654_ (.A(_135_),
    .B(_189_),
    .Y(_299_));
 sky130_fd_sc_hd__nand2_1 _655_ (.A(_135_),
    .B(_183_),
    .Y(_300_));
 sky130_fd_sc_hd__or4_1 _656_ (.A(_135_),
    .B(_154_),
    .C(_182_),
    .D(_189_),
    .X(_301_));
 sky130_fd_sc_hd__o211ai_1 _657_ (.A1(_202_),
    .A2(_299_),
    .B1(_300_),
    .C1(_301_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _658_ (.A(_196_),
    .B(_197_),
    .Y(_302_));
 sky130_fd_sc_hd__nor2_1 _659_ (.A(_202_),
    .B(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__o21ai_0 _660_ (.A1(_183_),
    .A2(_303_),
    .B1(net69),
    .Y(_304_));
 sky130_fd_sc_hd__o41ai_1 _661_ (.A1(net69),
    .A2(_175_),
    .A3(_196_),
    .A4(_197_),
    .B1(_304_),
    .Y(_039_));
 sky130_fd_sc_hd__a31oi_1 _662_ (.A1(_135_),
    .A2(net69),
    .A3(_185_),
    .B1(_192_),
    .Y(_305_));
 sky130_fd_sc_hd__o21ai_0 _663_ (.A1(_216_),
    .A2(_305_),
    .B1(net70),
    .Y(_306_));
 sky130_fd_sc_hd__o41ai_1 _664_ (.A1(net70),
    .A2(_175_),
    .A3(_189_),
    .A4(_190_),
    .B1(_306_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _665_ (.A(_195_),
    .B(_212_),
    .Y(_307_));
 sky130_fd_sc_hd__nor2_1 _666_ (.A(_192_),
    .B(_212_),
    .Y(_308_));
 sky130_fd_sc_hd__o21ai_0 _667_ (.A1(_182_),
    .A2(_308_),
    .B1(net71),
    .Y(_309_));
 sky130_fd_sc_hd__o21ai_0 _668_ (.A1(_176_),
    .A2(_307_),
    .B1(_309_),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_1 _669_ (.A(_202_),
    .B(_191_),
    .Y(_310_));
 sky130_fd_sc_hd__o21ai_0 _670_ (.A1(_209_),
    .A2(_310_),
    .B1(_133_),
    .Y(_311_));
 sky130_fd_sc_hd__o31ai_1 _671_ (.A1(_133_),
    .A2(_175_),
    .A3(_187_),
    .B1(_311_),
    .Y(_042_));
 sky130_fd_sc_hd__nand3_1 _672_ (.A(net71),
    .B(_133_),
    .C(_212_),
    .Y(_312_));
 sky130_fd_sc_hd__a31oi_1 _673_ (.A1(net71),
    .A2(_133_),
    .A3(_212_),
    .B1(_229_),
    .Y(_313_));
 sky130_fd_sc_hd__o21ai_0 _674_ (.A1(_209_),
    .A2(_313_),
    .B1(net73),
    .Y(_314_));
 sky130_fd_sc_hd__o31ai_1 _675_ (.A1(net73),
    .A2(_175_),
    .A3(_312_),
    .B1(_314_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _676_ (.A(_115_),
    .B(net112),
    .Y(_315_));
 sky130_fd_sc_hd__o21a_1 _677_ (.A1(_115_),
    .A2(_052_),
    .B1(_315_),
    .X(_316_));
 sky130_fd_sc_hd__o221a_1 _678_ (.A1(_075_),
    .A2(_315_),
    .B1(_316_),
    .B2(_074_),
    .C1(_073_),
    .X(_317_));
 sky130_fd_sc_hd__nand2_1 _679_ (.A(_052_),
    .B(_070_),
    .Y(_318_));
 sky130_fd_sc_hd__o31ai_1 _680_ (.A1(_070_),
    .A2(_080_),
    .A3(_317_),
    .B1(_318_),
    .Y(_044_));
 sky130_fd_sc_hd__a21boi_0 _681_ (.A1(_115_),
    .A2(_057_),
    .B1_N(_166_),
    .Y(_319_));
 sky130_fd_sc_hd__and2_0 _682_ (.A(_063_),
    .B(_178_),
    .X(_320_));
 sky130_fd_sc_hd__o21ai_0 _683_ (.A1(_114_),
    .A2(_320_),
    .B1(read_phase),
    .Y(_321_));
 sky130_fd_sc_hd__o41ai_1 _684_ (.A1(_114_),
    .A2(_169_),
    .A3(_319_),
    .A4(_320_),
    .B1(_321_),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_0 _685_ (.A1(_054_),
    .A2(_359_),
    .B1(_052_),
    .Y(_322_));
 sky130_fd_sc_hd__and3b_1 _686_ (.A_N(_052_),
    .B(_053_),
    .C(_074_),
    .X(_323_));
 sky130_fd_sc_hd__nor4_1 _687_ (.A(_074_),
    .B(_056_),
    .C(_054_),
    .D(net2),
    .Y(_324_));
 sky130_fd_sc_hd__a211o_1 _688_ (.A1(_075_),
    .A2(_322_),
    .B1(_323_),
    .C1(_324_),
    .X(_325_));
 sky130_fd_sc_hd__and2_0 _689_ (.A(_052_),
    .B(_359_),
    .X(_326_));
 sky130_fd_sc_hd__nand3b_1 _690_ (.A_N(_054_),
    .B(net2),
    .C(_068_),
    .Y(_327_));
 sky130_fd_sc_hd__o21ai_0 _691_ (.A1(_085_),
    .A2(_326_),
    .B1(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__a221o_1 _692_ (.A1(_069_),
    .A2(_325_),
    .B1(_328_),
    .B2(_081_),
    .C1(_086_),
    .X(_329_));
 sky130_fd_sc_hd__nand2b_1 _693_ (.A_N(_329_),
    .B(_069_),
    .Y(_330_));
 sky130_fd_sc_hd__nand2_1 _694_ (.A(_074_),
    .B(_329_),
    .Y(_331_));
 sky130_fd_sc_hd__o21ai_0 _695_ (.A1(_074_),
    .A2(_330_),
    .B1(_331_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _696_ (.A(_074_),
    .B(_114_),
    .Y(_332_));
 sky130_fd_sc_hd__o21ai_0 _697_ (.A1(_329_),
    .A2(_332_),
    .B1(_075_),
    .Y(_333_));
 sky130_fd_sc_hd__o31ai_1 _698_ (.A1(_063_),
    .A2(_075_),
    .A3(_330_),
    .B1(_333_),
    .Y(_047_));
 sky130_fd_sc_hd__nor3_1 _699_ (.A(_115_),
    .B(_076_),
    .C(_329_),
    .Y(_334_));
 sky130_fd_sc_hd__a21oi_1 _700_ (.A1(_115_),
    .A2(_076_),
    .B1(_334_),
    .Y(_335_));
 sky130_fd_sc_hd__nand2_1 _701_ (.A(_115_),
    .B(_329_),
    .Y(_336_));
 sky130_fd_sc_hd__o21ai_0 _702_ (.A1(_114_),
    .A2(_335_),
    .B1(_336_),
    .Y(_048_));
 sky130_fd_sc_hd__nand3_1 _703_ (.A(_114_),
    .B(net2),
    .C(_123_),
    .Y(_337_));
 sky130_fd_sc_hd__o41ai_1 _704_ (.A1(_114_),
    .A2(_116_),
    .A3(_076_),
    .A4(_329_),
    .B1(_337_),
    .Y(_049_));
 sky130_fd_sc_hd__a211oi_1 _705_ (.A1(_115_),
    .A2(_072_),
    .B1(_324_),
    .C1(_114_),
    .Y(_338_));
 sky130_fd_sc_hd__nand2_1 _706_ (.A(_075_),
    .B(_052_),
    .Y(_339_));
 sky130_fd_sc_hd__maj3_1 _707_ (.A(read_phase),
    .B(_115_),
    .C(_072_),
    .X(_340_));
 sky130_fd_sc_hd__a21oi_1 _708_ (.A1(_320_),
    .A2(_339_),
    .B1(_340_),
    .Y(_341_));
 sky130_fd_sc_hd__a2bb2oi_1 _709_ (.A1_N(net112),
    .A2_N(_338_),
    .B1(_341_),
    .B2(_069_),
    .Y(_050_));
 sky130_fd_sc_hd__o211ai_1 _710_ (.A1(_063_),
    .A2(_069_),
    .B1(_116_),
    .C1(_177_),
    .Y(net79));
 sky130_fd_sc_hd__nand2b_4 _711_ (.A_N(_080_),
    .B(_063_),
    .Y(net104));
 sky130_fd_sc_hd__ha_1 _712_ (.A(_342_),
    .B(_343_),
    .COUT(_344_),
    .SUM(_345_));
 sky130_fd_sc_hd__ha_1 _713_ (.A(net42),
    .B(net53),
    .COUT(_346_),
    .SUM(_347_));
 sky130_fd_sc_hd__ha_1 _714_ (.A(_348_),
    .B(_349_),
    .COUT(_350_),
    .SUM(_351_));
 sky130_fd_sc_hd__ha_1 _715_ (.A(net74),
    .B(net75),
    .COUT(_352_),
    .SUM(_353_));
 sky130_fd_sc_hd__ha_1 _716_ (.A(_354_),
    .B(_355_),
    .COUT(_356_),
    .SUM(_357_));
 sky130_fd_sc_hd__ha_1 _717_ (.A(net78),
    .B(_358_),
    .COUT(_359_),
    .SUM(_360_));
 sky130_fd_sc_hd__clkbuf_1 _718_ (.A(net104),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _719_ (.A(net104),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _720_ (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _721_ (.A(net104),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _722_ (.A(net104),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _723_ (.A(net104),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 _724_ (.A(net104),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _725_ (.A(net104),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _726_ (.A(net104),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 _727_ (.A(net104),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 _728_ (.A(net104),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _729_ (.A(net104),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _730_ (.A(net104),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _731_ (.A(net104),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _732_ (.A(net104),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _733_ (.A(net104),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _734_ (.A(net104),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _735_ (.A(net104),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _736_ (.A(net104),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _737_ (.A(net104),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _738_ (.A(net104),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _739_ (.A(net104),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _740_ (.A(net104),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _741_ (.A(net104),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _742_ (.A(net104),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _743_ (.A(net104),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _744_ (.A(net104),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _745_ (.A(net104),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _746_ (.A(net104),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _747_ (.A(net104),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _748_ (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__dfrtp_2 \addr_counter[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(net74),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \addr_counter[1]$_DFFE_PN0P_  (.D(_001_),
    .Q(net75),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \addr_counter[2]$_DFFE_PN0P_  (.D(_002_),
    .Q(net76),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \addr_counter[3]$_DFFE_PN0P_  (.D(_003_),
    .Q(net77),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \addr_counter[4]$_DFFE_PN0P_  (.D(_004_),
    .Q(net78),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \bist_done$_DFFE_PN0P_  (.D(_005_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \bist_pass$_DFFE_PN0P_  (.D(_006_),
    .Q(net36),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_addr[0]$_DFFE_PN0P_  (.D(_007_),
    .Q(net37),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_addr[1]$_DFFE_PN0P_  (.D(_008_),
    .Q(net38),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_addr[2]$_DFFE_PN0P_  (.D(_009_),
    .Q(net39),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_addr[3]$_DFFE_PN0P_  (.D(_010_),
    .Q(net40),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_addr[4]$_DFFE_PN0P_  (.D(_011_),
    .Q(net41),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[0]$_DFFE_PN0P_  (.D(_012_),
    .Q(net42),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[10]$_DFFE_PN0P_  (.D(_013_),
    .Q(net43),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[11]$_DFFE_PN0P_  (.D(_014_),
    .Q(net44),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[12]$_DFFE_PN0P_  (.D(_015_),
    .Q(net45),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[13]$_DFFE_PN0P_  (.D(_016_),
    .Q(net46),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[14]$_DFFE_PN0P_  (.D(_017_),
    .Q(net47),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[15]$_DFFE_PN0P_  (.D(_018_),
    .Q(net48),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[16]$_DFFE_PN0P_  (.D(_019_),
    .Q(net49),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[17]$_DFFE_PN0P_  (.D(_020_),
    .Q(net50),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[18]$_DFFE_PN0P_  (.D(_021_),
    .Q(net51),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[19]$_DFFE_PN0P_  (.D(_022_),
    .Q(net52),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(net53),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[20]$_DFFE_PN0P_  (.D(_024_),
    .Q(net54),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[21]$_DFFE_PN0P_  (.D(_025_),
    .Q(net55),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[22]$_DFFE_PN0P_  (.D(_026_),
    .Q(net56),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[23]$_DFFE_PN0P_  (.D(_027_),
    .Q(net57),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[24]$_DFFE_PN0P_  (.D(_028_),
    .Q(net58),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[25]$_DFFE_PN0P_  (.D(_029_),
    .Q(net59),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[26]$_DFFE_PN0P_  (.D(_030_),
    .Q(net60),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[27]$_DFFE_PN0P_  (.D(_031_),
    .Q(net61),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[28]$_DFFE_PN0P_  (.D(_032_),
    .Q(net62),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \error_count[29]$_DFFE_PN0P_  (.D(_033_),
    .Q(net63),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[2]$_DFFE_PN0P_  (.D(_034_),
    .Q(net64),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[30]$_DFFE_PN0P_  (.D(_035_),
    .Q(net65),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[31]$_DFFE_PN0P_  (.D(_036_),
    .Q(net66),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[3]$_DFFE_PN0P_  (.D(_037_),
    .Q(net67),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[4]$_DFFE_PN0P_  (.D(_038_),
    .Q(net68),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \error_count[5]$_DFFE_PN0P_  (.D(_039_),
    .Q(net69),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[6]$_DFFE_PN0P_  (.D(_040_),
    .Q(net70),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[7]$_DFFE_PN0P_  (.D(_041_),
    .Q(net71),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[8]$_DFFE_PN0P_  (.D(_042_),
    .Q(net72),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[9]$_DFFE_PN0P_  (.D(_043_),
    .Q(net73),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \phase_complete$_DFFE_PN0P_  (.D(_044_),
    .Q(phase_complete),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \read_phase$_DFFE_PN0P_  (.D(_045_),
    .Q(read_phase),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_046_),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_047_),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \state[2]$_DFFE_PN0P_  (.D(_048_),
    .Q(\state[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[3]$_DFFE_PN0P_  (.D(_049_),
    .Q(\state[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \write_phase$_DFFE_PN0P_  (.D(_050_),
    .Q(net112),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net113),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_76 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(bist_start),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(mem_rdata[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(mem_rdata[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(mem_rdata[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(mem_rdata[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(mem_rdata[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(mem_rdata[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(mem_rdata[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(mem_rdata[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(mem_rdata[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(mem_rdata[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(mem_rdata[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(mem_rdata[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(mem_rdata[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(mem_rdata[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(mem_rdata[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(mem_rdata[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(mem_rdata[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(mem_rdata[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(mem_rdata[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(mem_rdata[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(mem_rdata[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(mem_rdata[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(mem_rdata[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(mem_rdata[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(mem_rdata[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(mem_rdata[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(mem_rdata[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(mem_rdata[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(mem_rdata[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(mem_rdata[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(mem_rdata[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(mem_rdata[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(bist_done));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(bist_pass));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(error_addr[0]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(error_addr[1]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(error_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(error_addr[3]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(error_addr[4]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(error_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(error_count[10]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(error_count[11]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(error_count[12]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(error_count[13]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(error_count[14]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(error_count[15]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(error_count[16]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(error_count[17]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(error_count[18]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(error_count[19]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(error_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(error_count[20]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net55),
    .X(error_count[21]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net56),
    .X(error_count[22]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net57),
    .X(error_count[23]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net58),
    .X(error_count[24]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net59),
    .X(error_count[25]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net60),
    .X(error_count[26]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net61),
    .X(error_count[27]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net62),
    .X(error_count[28]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net63),
    .X(error_count[29]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net64),
    .X(error_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net65),
    .X(error_count[30]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net66),
    .X(error_count[31]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net67),
    .X(error_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(error_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(error_count[5]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(error_count[6]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(error_count[7]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(error_count[8]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(error_count[9]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(mem_enable));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net100),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net101),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net105),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net106),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net107),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net108),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net109),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net110),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net111),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net112),
    .X(mem_write));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net113));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_174 ();
endmodule
