module configurable_brent_kung_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 INV_X1 _070_ (.A(net1),
    .ZN(_000_));
 INV_X1 _071_ (.A(net25),
    .ZN(_052_));
 INV_X1 _072_ (.A(net33),
    .ZN(_001_));
 INV_X1 _073_ (.A(net57),
    .ZN(_053_));
 INV_X1 _074_ (.A(net65),
    .ZN(_002_));
 INV_X1 _075_ (.A(_006_),
    .ZN(net68));
 INV_X1 _076_ (.A(_008_),
    .ZN(net69));
 INV_X1 _077_ (.A(_010_),
    .ZN(net70));
 INV_X1 _078_ (.A(_012_),
    .ZN(net71));
 INV_X1 _079_ (.A(_014_),
    .ZN(net72));
 INV_X1 _080_ (.A(_016_),
    .ZN(net73));
 INV_X1 _081_ (.A(_018_),
    .ZN(net74));
 INV_X1 _082_ (.A(_020_),
    .ZN(net75));
 INV_X1 _083_ (.A(_022_),
    .ZN(net76));
 INV_X1 _084_ (.A(_024_),
    .ZN(net77));
 INV_X1 _085_ (.A(_027_),
    .ZN(net78));
 INV_X1 _086_ (.A(_029_),
    .ZN(net79));
 INV_X1 _087_ (.A(_031_),
    .ZN(net80));
 INV_X1 _088_ (.A(_033_),
    .ZN(net81));
 INV_X1 _089_ (.A(_035_),
    .ZN(net82));
 INV_X1 _090_ (.A(_037_),
    .ZN(net83));
 INV_X1 _091_ (.A(_039_),
    .ZN(net84));
 INV_X1 _092_ (.A(_041_),
    .ZN(net85));
 INV_X1 _093_ (.A(_043_),
    .ZN(net86));
 INV_X1 _094_ (.A(_045_),
    .ZN(net87));
 INV_X1 _095_ (.A(_047_),
    .ZN(net88));
 INV_X1 _096_ (.A(_049_),
    .ZN(net89));
 INV_X1 _097_ (.A(_051_),
    .ZN(net90));
 INV_X1 _098_ (.A(_056_),
    .ZN(net91));
 INV_X1 _099_ (.A(_058_),
    .ZN(net92));
 INV_X1 _100_ (.A(_060_),
    .ZN(net93));
 INV_X1 _101_ (.A(_062_),
    .ZN(net94));
 INV_X1 _102_ (.A(_064_),
    .ZN(net95));
 INV_X1 _103_ (.A(_066_),
    .ZN(net96));
 INV_X1 _104_ (.A(_068_),
    .ZN(net97));
 INV_X1 _105_ (.A(_069_),
    .ZN(net98));
 INV_X1 _106_ (.A(_050_),
    .ZN(_054_));
 INV_X1 _107_ (.A(_055_),
    .ZN(net66));
 INV_X1 _108_ (.A(_003_),
    .ZN(_025_));
 FA_X1 _109_ (.A(_000_),
    .B(_001_),
    .CI(_002_),
    .CO(_003_),
    .S(net67));
 FA_X1 _110_ (.A(net2),
    .B(net34),
    .CI(_004_),
    .CO(_005_),
    .S(_006_));
 FA_X1 _111_ (.A(net3),
    .B(net35),
    .CI(_005_),
    .CO(_007_),
    .S(_008_));
 FA_X1 _112_ (.A(net4),
    .B(net36),
    .CI(_007_),
    .CO(_009_),
    .S(_010_));
 FA_X1 _113_ (.A(net5),
    .B(net37),
    .CI(_009_),
    .CO(_011_),
    .S(_012_));
 FA_X1 _114_ (.A(net6),
    .B(net38),
    .CI(_011_),
    .CO(_013_),
    .S(_014_));
 FA_X1 _115_ (.A(net7),
    .B(net39),
    .CI(_013_),
    .CO(_015_),
    .S(_016_));
 FA_X1 _116_ (.A(net8),
    .B(net40),
    .CI(_015_),
    .CO(_017_),
    .S(_018_));
 FA_X1 _117_ (.A(net9),
    .B(net41),
    .CI(_017_),
    .CO(_019_),
    .S(_020_));
 FA_X1 _118_ (.A(net10),
    .B(net42),
    .CI(_019_),
    .CO(_021_),
    .S(_022_));
 FA_X1 _119_ (.A(net11),
    .B(net43),
    .CI(_021_),
    .CO(_023_),
    .S(_024_));
 FA_X1 _120_ (.A(net12),
    .B(net44),
    .CI(_025_),
    .CO(_026_),
    .S(_027_));
 FA_X1 _121_ (.A(net13),
    .B(net45),
    .CI(_023_),
    .CO(_028_),
    .S(_029_));
 FA_X1 _122_ (.A(net14),
    .B(net46),
    .CI(_028_),
    .CO(_030_),
    .S(_031_));
 FA_X1 _123_ (.A(net15),
    .B(net47),
    .CI(_030_),
    .CO(_032_),
    .S(_033_));
 FA_X1 _124_ (.A(net16),
    .B(net48),
    .CI(_032_),
    .CO(_034_),
    .S(_035_));
 FA_X1 _125_ (.A(net17),
    .B(net49),
    .CI(_034_),
    .CO(_036_),
    .S(_037_));
 FA_X1 _126_ (.A(net18),
    .B(net50),
    .CI(_036_),
    .CO(_038_),
    .S(_039_));
 FA_X1 _127_ (.A(net19),
    .B(net51),
    .CI(_038_),
    .CO(_040_),
    .S(_041_));
 FA_X1 _128_ (.A(net20),
    .B(net52),
    .CI(_040_),
    .CO(_042_),
    .S(_043_));
 FA_X1 _129_ (.A(net21),
    .B(net53),
    .CI(_042_),
    .CO(_044_),
    .S(_045_));
 FA_X1 _130_ (.A(net22),
    .B(net54),
    .CI(_044_),
    .CO(_046_),
    .S(_047_));
 FA_X1 _131_ (.A(net23),
    .B(net55),
    .CI(_026_),
    .CO(_048_),
    .S(_049_));
 FA_X1 _132_ (.A(net24),
    .B(net56),
    .CI(_046_),
    .CO(_050_),
    .S(_051_));
 FA_X1 _133_ (.A(_052_),
    .B(_053_),
    .CI(_054_),
    .CO(_055_),
    .S(_056_));
 FA_X1 _134_ (.A(net26),
    .B(net58),
    .CI(_048_),
    .CO(_057_),
    .S(_058_));
 FA_X1 _135_ (.A(net27),
    .B(net59),
    .CI(_057_),
    .CO(_059_),
    .S(_060_));
 FA_X1 _136_ (.A(net28),
    .B(net60),
    .CI(_059_),
    .CO(_061_),
    .S(_062_));
 FA_X1 _137_ (.A(net29),
    .B(net61),
    .CI(_061_),
    .CO(_063_),
    .S(_064_));
 FA_X1 _138_ (.A(net30),
    .B(net62),
    .CI(_063_),
    .CO(_065_),
    .S(_066_));
 FA_X1 _139_ (.A(net31),
    .B(net63),
    .CI(_065_),
    .CO(_067_),
    .S(_068_));
 FA_X1 _140_ (.A(net32),
    .B(net64),
    .CI(_067_),
    .CO(_004_),
    .S(_069_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_111 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 BUF_X1 input2 (.A(a[10]),
    .Z(net2));
 BUF_X1 input3 (.A(a[11]),
    .Z(net3));
 BUF_X1 input4 (.A(a[12]),
    .Z(net4));
 BUF_X1 input5 (.A(a[13]),
    .Z(net5));
 BUF_X1 input6 (.A(a[14]),
    .Z(net6));
 BUF_X1 input7 (.A(a[15]),
    .Z(net7));
 BUF_X1 input8 (.A(a[16]),
    .Z(net8));
 BUF_X1 input9 (.A(a[17]),
    .Z(net9));
 BUF_X1 input10 (.A(a[18]),
    .Z(net10));
 BUF_X1 input11 (.A(a[19]),
    .Z(net11));
 BUF_X1 input12 (.A(a[1]),
    .Z(net12));
 BUF_X1 input13 (.A(a[20]),
    .Z(net13));
 BUF_X1 input14 (.A(a[21]),
    .Z(net14));
 BUF_X1 input15 (.A(a[22]),
    .Z(net15));
 BUF_X1 input16 (.A(a[23]),
    .Z(net16));
 BUF_X1 input17 (.A(a[24]),
    .Z(net17));
 BUF_X1 input18 (.A(a[25]),
    .Z(net18));
 BUF_X1 input19 (.A(a[26]),
    .Z(net19));
 BUF_X1 input20 (.A(a[27]),
    .Z(net20));
 BUF_X1 input21 (.A(a[28]),
    .Z(net21));
 BUF_X1 input22 (.A(a[29]),
    .Z(net22));
 BUF_X1 input23 (.A(a[2]),
    .Z(net23));
 BUF_X1 input24 (.A(a[30]),
    .Z(net24));
 BUF_X1 input25 (.A(a[31]),
    .Z(net25));
 BUF_X1 input26 (.A(a[3]),
    .Z(net26));
 BUF_X1 input27 (.A(a[4]),
    .Z(net27));
 BUF_X1 input28 (.A(a[5]),
    .Z(net28));
 BUF_X1 input29 (.A(a[6]),
    .Z(net29));
 BUF_X1 input30 (.A(a[7]),
    .Z(net30));
 BUF_X1 input31 (.A(a[8]),
    .Z(net31));
 BUF_X1 input32 (.A(a[9]),
    .Z(net32));
 BUF_X1 input33 (.A(b[0]),
    .Z(net33));
 BUF_X1 input34 (.A(b[10]),
    .Z(net34));
 BUF_X1 input35 (.A(b[11]),
    .Z(net35));
 BUF_X1 input36 (.A(b[12]),
    .Z(net36));
 BUF_X1 input37 (.A(b[13]),
    .Z(net37));
 BUF_X1 input38 (.A(b[14]),
    .Z(net38));
 BUF_X1 input39 (.A(b[15]),
    .Z(net39));
 BUF_X1 input40 (.A(b[16]),
    .Z(net40));
 BUF_X1 input41 (.A(b[17]),
    .Z(net41));
 BUF_X1 input42 (.A(b[18]),
    .Z(net42));
 BUF_X1 input43 (.A(b[19]),
    .Z(net43));
 BUF_X1 input44 (.A(b[1]),
    .Z(net44));
 BUF_X1 input45 (.A(b[20]),
    .Z(net45));
 BUF_X1 input46 (.A(b[21]),
    .Z(net46));
 BUF_X1 input47 (.A(b[22]),
    .Z(net47));
 BUF_X1 input48 (.A(b[23]),
    .Z(net48));
 BUF_X1 input49 (.A(b[24]),
    .Z(net49));
 BUF_X1 input50 (.A(b[25]),
    .Z(net50));
 BUF_X1 input51 (.A(b[26]),
    .Z(net51));
 BUF_X1 input52 (.A(b[27]),
    .Z(net52));
 BUF_X1 input53 (.A(b[28]),
    .Z(net53));
 BUF_X1 input54 (.A(b[29]),
    .Z(net54));
 BUF_X1 input55 (.A(b[2]),
    .Z(net55));
 BUF_X1 input56 (.A(b[30]),
    .Z(net56));
 BUF_X1 input57 (.A(b[31]),
    .Z(net57));
 BUF_X1 input58 (.A(b[3]),
    .Z(net58));
 BUF_X1 input59 (.A(b[4]),
    .Z(net59));
 BUF_X1 input60 (.A(b[5]),
    .Z(net60));
 BUF_X1 input61 (.A(b[6]),
    .Z(net61));
 BUF_X1 input62 (.A(b[7]),
    .Z(net62));
 BUF_X1 input63 (.A(b[8]),
    .Z(net63));
 BUF_X1 input64 (.A(b[9]),
    .Z(net64));
 BUF_X1 input65 (.A(cin),
    .Z(net65));
 BUF_X1 output66 (.A(net66),
    .Z(cout));
 BUF_X1 output67 (.A(net67),
    .Z(sum[0]));
 BUF_X1 output68 (.A(net68),
    .Z(sum[10]));
 BUF_X1 output69 (.A(net69),
    .Z(sum[11]));
 BUF_X1 output70 (.A(net70),
    .Z(sum[12]));
 BUF_X1 output71 (.A(net71),
    .Z(sum[13]));
 BUF_X1 output72 (.A(net72),
    .Z(sum[14]));
 BUF_X1 output73 (.A(net73),
    .Z(sum[15]));
 BUF_X1 output74 (.A(net74),
    .Z(sum[16]));
 BUF_X1 output75 (.A(net75),
    .Z(sum[17]));
 BUF_X1 output76 (.A(net76),
    .Z(sum[18]));
 BUF_X1 output77 (.A(net77),
    .Z(sum[19]));
 BUF_X1 output78 (.A(net78),
    .Z(sum[1]));
 BUF_X1 output79 (.A(net79),
    .Z(sum[20]));
 BUF_X1 output80 (.A(net80),
    .Z(sum[21]));
 BUF_X1 output81 (.A(net81),
    .Z(sum[22]));
 BUF_X1 output82 (.A(net82),
    .Z(sum[23]));
 BUF_X1 output83 (.A(net83),
    .Z(sum[24]));
 BUF_X1 output84 (.A(net84),
    .Z(sum[25]));
 BUF_X1 output85 (.A(net85),
    .Z(sum[26]));
 BUF_X1 output86 (.A(net86),
    .Z(sum[27]));
 BUF_X1 output87 (.A(net87),
    .Z(sum[28]));
 BUF_X1 output88 (.A(net88),
    .Z(sum[29]));
 BUF_X1 output89 (.A(net89),
    .Z(sum[2]));
 BUF_X1 output90 (.A(net90),
    .Z(sum[30]));
 BUF_X1 output91 (.A(net91),
    .Z(sum[31]));
 BUF_X1 output92 (.A(net92),
    .Z(sum[3]));
 BUF_X1 output93 (.A(net93),
    .Z(sum[4]));
 BUF_X1 output94 (.A(net94),
    .Z(sum[5]));
 BUF_X1 output95 (.A(net95),
    .Z(sum[6]));
 BUF_X1 output96 (.A(net96),
    .Z(sum[7]));
 BUF_X1 output97 (.A(net97),
    .Z(sum[8]));
 BUF_X1 output98 (.A(net98),
    .Z(sum[9]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X2 FILLER_0_417 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X2 FILLER_1_417 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X2 FILLER_2_417 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X2 FILLER_3_417 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X2 FILLER_4_417 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X2 FILLER_5_417 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X2 FILLER_6_417 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X2 FILLER_7_417 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X2 FILLER_8_417 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X2 FILLER_9_417 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X2 FILLER_10_417 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X2 FILLER_11_417 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X2 FILLER_12_417 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X2 FILLER_13_417 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X2 FILLER_14_417 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_417 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X4 FILLER_16_385 ();
 FILLCELL_X1 FILLER_16_389 ();
 FILLCELL_X2 FILLER_16_406 ();
 FILLCELL_X8 FILLER_16_410 ();
 FILLCELL_X1 FILLER_16_418 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X4 FILLER_17_385 ();
 FILLCELL_X2 FILLER_17_389 ();
 FILLCELL_X2 FILLER_17_407 ();
 FILLCELL_X1 FILLER_17_409 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X2 FILLER_18_385 ();
 FILLCELL_X1 FILLER_18_406 ();
 FILLCELL_X1 FILLER_18_409 ();
 FILLCELL_X1 FILLER_18_415 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X8 FILLER_19_385 ();
 FILLCELL_X2 FILLER_19_393 ();
 FILLCELL_X1 FILLER_19_395 ();
 FILLCELL_X8 FILLER_19_399 ();
 FILLCELL_X4 FILLER_19_407 ();
 FILLCELL_X2 FILLER_19_416 ();
 FILLCELL_X1 FILLER_19_418 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X8 FILLER_20_385 ();
 FILLCELL_X4 FILLER_20_393 ();
 FILLCELL_X1 FILLER_20_397 ();
 FILLCELL_X8 FILLER_20_401 ();
 FILLCELL_X2 FILLER_20_412 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_5 ();
 FILLCELL_X1 FILLER_21_7 ();
 FILLCELL_X32 FILLER_21_27 ();
 FILLCELL_X32 FILLER_21_59 ();
 FILLCELL_X32 FILLER_21_91 ();
 FILLCELL_X32 FILLER_21_123 ();
 FILLCELL_X32 FILLER_21_155 ();
 FILLCELL_X32 FILLER_21_187 ();
 FILLCELL_X32 FILLER_21_219 ();
 FILLCELL_X32 FILLER_21_251 ();
 FILLCELL_X32 FILLER_21_283 ();
 FILLCELL_X32 FILLER_21_315 ();
 FILLCELL_X32 FILLER_21_347 ();
 FILLCELL_X8 FILLER_21_379 ();
 FILLCELL_X4 FILLER_21_387 ();
 FILLCELL_X2 FILLER_21_407 ();
 FILLCELL_X1 FILLER_21_412 ();
 FILLCELL_X1 FILLER_21_415 ();
 FILLCELL_X1 FILLER_22_28 ();
 FILLCELL_X4 FILLER_22_31 ();
 FILLCELL_X2 FILLER_22_35 ();
 FILLCELL_X1 FILLER_22_37 ();
 FILLCELL_X32 FILLER_22_41 ();
 FILLCELL_X32 FILLER_22_73 ();
 FILLCELL_X32 FILLER_22_105 ();
 FILLCELL_X32 FILLER_22_137 ();
 FILLCELL_X32 FILLER_22_169 ();
 FILLCELL_X32 FILLER_22_201 ();
 FILLCELL_X32 FILLER_22_233 ();
 FILLCELL_X32 FILLER_22_265 ();
 FILLCELL_X32 FILLER_22_297 ();
 FILLCELL_X32 FILLER_22_329 ();
 FILLCELL_X16 FILLER_22_361 ();
 FILLCELL_X2 FILLER_22_377 ();
 FILLCELL_X1 FILLER_22_379 ();
 FILLCELL_X4 FILLER_22_396 ();
 FILLCELL_X1 FILLER_22_400 ();
 FILLCELL_X2 FILLER_22_404 ();
 FILLCELL_X1 FILLER_22_406 ();
 FILLCELL_X4 FILLER_22_415 ();
 FILLCELL_X2 FILLER_23_9 ();
 FILLCELL_X4 FILLER_23_30 ();
 FILLCELL_X1 FILLER_23_34 ();
 FILLCELL_X32 FILLER_23_51 ();
 FILLCELL_X32 FILLER_23_83 ();
 FILLCELL_X32 FILLER_23_115 ();
 FILLCELL_X32 FILLER_23_147 ();
 FILLCELL_X32 FILLER_23_179 ();
 FILLCELL_X32 FILLER_23_211 ();
 FILLCELL_X32 FILLER_23_243 ();
 FILLCELL_X32 FILLER_23_275 ();
 FILLCELL_X32 FILLER_23_307 ();
 FILLCELL_X32 FILLER_23_339 ();
 FILLCELL_X4 FILLER_23_371 ();
 FILLCELL_X1 FILLER_23_375 ();
 FILLCELL_X1 FILLER_23_415 ();
 FILLCELL_X32 FILLER_24_30 ();
 FILLCELL_X32 FILLER_24_62 ();
 FILLCELL_X32 FILLER_24_94 ();
 FILLCELL_X32 FILLER_24_126 ();
 FILLCELL_X32 FILLER_24_158 ();
 FILLCELL_X32 FILLER_24_190 ();
 FILLCELL_X32 FILLER_24_222 ();
 FILLCELL_X32 FILLER_24_254 ();
 FILLCELL_X32 FILLER_24_286 ();
 FILLCELL_X32 FILLER_24_318 ();
 FILLCELL_X32 FILLER_24_350 ();
 FILLCELL_X4 FILLER_24_382 ();
 FILLCELL_X1 FILLER_24_386 ();
 FILLCELL_X16 FILLER_24_392 ();
 FILLCELL_X2 FILLER_24_408 ();
 FILLCELL_X2 FILLER_24_413 ();
 FILLCELL_X1 FILLER_24_415 ();
 FILLCELL_X1 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_5 ();
 FILLCELL_X1 FILLER_25_12 ();
 FILLCELL_X32 FILLER_25_16 ();
 FILLCELL_X32 FILLER_25_48 ();
 FILLCELL_X32 FILLER_25_80 ();
 FILLCELL_X32 FILLER_25_112 ();
 FILLCELL_X32 FILLER_25_144 ();
 FILLCELL_X32 FILLER_25_176 ();
 FILLCELL_X32 FILLER_25_208 ();
 FILLCELL_X32 FILLER_25_240 ();
 FILLCELL_X32 FILLER_25_272 ();
 FILLCELL_X32 FILLER_25_304 ();
 FILLCELL_X32 FILLER_25_336 ();
 FILLCELL_X32 FILLER_25_368 ();
 FILLCELL_X1 FILLER_25_403 ();
 FILLCELL_X8 FILLER_25_407 ();
 FILLCELL_X4 FILLER_25_415 ();
 FILLCELL_X8 FILLER_26_1 ();
 FILLCELL_X1 FILLER_26_9 ();
 FILLCELL_X32 FILLER_26_13 ();
 FILLCELL_X32 FILLER_26_45 ();
 FILLCELL_X32 FILLER_26_77 ();
 FILLCELL_X32 FILLER_26_109 ();
 FILLCELL_X32 FILLER_26_141 ();
 FILLCELL_X8 FILLER_26_173 ();
 FILLCELL_X32 FILLER_26_183 ();
 FILLCELL_X32 FILLER_26_215 ();
 FILLCELL_X32 FILLER_26_247 ();
 FILLCELL_X32 FILLER_26_279 ();
 FILLCELL_X32 FILLER_26_311 ();
 FILLCELL_X32 FILLER_26_343 ();
 FILLCELL_X8 FILLER_26_375 ();
 FILLCELL_X4 FILLER_26_383 ();
 FILLCELL_X2 FILLER_26_387 ();
 FILLCELL_X4 FILLER_26_405 ();
 FILLCELL_X1 FILLER_26_409 ();
 FILLCELL_X1 FILLER_26_413 ();
 FILLCELL_X2 FILLER_27_7 ();
 FILLCELL_X1 FILLER_27_28 ();
 FILLCELL_X32 FILLER_27_31 ();
 FILLCELL_X32 FILLER_27_63 ();
 FILLCELL_X32 FILLER_27_95 ();
 FILLCELL_X32 FILLER_27_127 ();
 FILLCELL_X32 FILLER_27_159 ();
 FILLCELL_X32 FILLER_27_191 ();
 FILLCELL_X32 FILLER_27_223 ();
 FILLCELL_X32 FILLER_27_255 ();
 FILLCELL_X32 FILLER_27_287 ();
 FILLCELL_X32 FILLER_27_319 ();
 FILLCELL_X32 FILLER_27_351 ();
 FILLCELL_X16 FILLER_27_383 ();
 FILLCELL_X4 FILLER_27_399 ();
 FILLCELL_X8 FILLER_27_408 ();
 FILLCELL_X32 FILLER_28_20 ();
 FILLCELL_X32 FILLER_28_52 ();
 FILLCELL_X32 FILLER_28_84 ();
 FILLCELL_X32 FILLER_28_116 ();
 FILLCELL_X32 FILLER_28_148 ();
 FILLCELL_X32 FILLER_28_180 ();
 FILLCELL_X32 FILLER_28_212 ();
 FILLCELL_X32 FILLER_28_244 ();
 FILLCELL_X32 FILLER_28_276 ();
 FILLCELL_X32 FILLER_28_308 ();
 FILLCELL_X32 FILLER_28_340 ();
 FILLCELL_X8 FILLER_28_372 ();
 FILLCELL_X4 FILLER_28_380 ();
 FILLCELL_X2 FILLER_28_384 ();
 FILLCELL_X1 FILLER_28_386 ();
 FILLCELL_X2 FILLER_28_406 ();
 FILLCELL_X4 FILLER_28_414 ();
 FILLCELL_X1 FILLER_28_418 ();
 FILLCELL_X32 FILLER_29_28 ();
 FILLCELL_X32 FILLER_29_60 ();
 FILLCELL_X32 FILLER_29_92 ();
 FILLCELL_X32 FILLER_29_124 ();
 FILLCELL_X32 FILLER_29_156 ();
 FILLCELL_X32 FILLER_29_188 ();
 FILLCELL_X32 FILLER_29_220 ();
 FILLCELL_X32 FILLER_29_252 ();
 FILLCELL_X32 FILLER_29_284 ();
 FILLCELL_X32 FILLER_29_316 ();
 FILLCELL_X32 FILLER_29_348 ();
 FILLCELL_X8 FILLER_29_380 ();
 FILLCELL_X2 FILLER_29_388 ();
 FILLCELL_X1 FILLER_29_390 ();
 FILLCELL_X1 FILLER_29_410 ();
 FILLCELL_X1 FILLER_30_6 ();
 FILLCELL_X1 FILLER_30_10 ();
 FILLCELL_X32 FILLER_30_27 ();
 FILLCELL_X32 FILLER_30_59 ();
 FILLCELL_X32 FILLER_30_91 ();
 FILLCELL_X32 FILLER_30_123 ();
 FILLCELL_X32 FILLER_30_155 ();
 FILLCELL_X32 FILLER_30_187 ();
 FILLCELL_X32 FILLER_30_219 ();
 FILLCELL_X32 FILLER_30_251 ();
 FILLCELL_X32 FILLER_30_283 ();
 FILLCELL_X32 FILLER_30_315 ();
 FILLCELL_X32 FILLER_30_347 ();
 FILLCELL_X16 FILLER_30_379 ();
 FILLCELL_X2 FILLER_30_395 ();
 FILLCELL_X4 FILLER_30_415 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X2 FILLER_31_5 ();
 FILLCELL_X1 FILLER_31_7 ();
 FILLCELL_X32 FILLER_31_11 ();
 FILLCELL_X32 FILLER_31_43 ();
 FILLCELL_X32 FILLER_31_75 ();
 FILLCELL_X32 FILLER_31_107 ();
 FILLCELL_X32 FILLER_31_139 ();
 FILLCELL_X32 FILLER_31_171 ();
 FILLCELL_X32 FILLER_31_203 ();
 FILLCELL_X32 FILLER_31_235 ();
 FILLCELL_X32 FILLER_31_267 ();
 FILLCELL_X32 FILLER_31_299 ();
 FILLCELL_X32 FILLER_31_331 ();
 FILLCELL_X16 FILLER_31_363 ();
 FILLCELL_X8 FILLER_31_379 ();
 FILLCELL_X4 FILLER_31_387 ();
 FILLCELL_X1 FILLER_31_391 ();
 FILLCELL_X8 FILLER_31_395 ();
 FILLCELL_X4 FILLER_31_403 ();
 FILLCELL_X2 FILLER_31_407 ();
 FILLCELL_X1 FILLER_31_409 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_6 ();
 FILLCELL_X2 FILLER_32_14 ();
 FILLCELL_X1 FILLER_32_27 ();
 FILLCELL_X1 FILLER_32_35 ();
 FILLCELL_X32 FILLER_32_54 ();
 FILLCELL_X32 FILLER_32_86 ();
 FILLCELL_X32 FILLER_32_118 ();
 FILLCELL_X32 FILLER_32_150 ();
 FILLCELL_X32 FILLER_32_182 ();
 FILLCELL_X32 FILLER_32_214 ();
 FILLCELL_X32 FILLER_32_246 ();
 FILLCELL_X32 FILLER_32_278 ();
 FILLCELL_X32 FILLER_32_310 ();
 FILLCELL_X32 FILLER_32_342 ();
 FILLCELL_X4 FILLER_32_374 ();
 FILLCELL_X1 FILLER_33_1 ();
 FILLCELL_X2 FILLER_33_11 ();
 FILLCELL_X2 FILLER_33_15 ();
 FILLCELL_X1 FILLER_33_22 ();
 FILLCELL_X1 FILLER_33_39 ();
 FILLCELL_X32 FILLER_33_42 ();
 FILLCELL_X32 FILLER_33_74 ();
 FILLCELL_X32 FILLER_33_106 ();
 FILLCELL_X32 FILLER_33_138 ();
 FILLCELL_X32 FILLER_33_170 ();
 FILLCELL_X32 FILLER_33_202 ();
 FILLCELL_X32 FILLER_33_234 ();
 FILLCELL_X32 FILLER_33_266 ();
 FILLCELL_X32 FILLER_33_298 ();
 FILLCELL_X32 FILLER_33_330 ();
 FILLCELL_X16 FILLER_33_362 ();
 FILLCELL_X8 FILLER_33_378 ();
 FILLCELL_X4 FILLER_33_386 ();
 FILLCELL_X2 FILLER_33_411 ();
 FILLCELL_X32 FILLER_34_20 ();
 FILLCELL_X32 FILLER_34_52 ();
 FILLCELL_X32 FILLER_34_84 ();
 FILLCELL_X32 FILLER_34_116 ();
 FILLCELL_X32 FILLER_34_148 ();
 FILLCELL_X32 FILLER_34_180 ();
 FILLCELL_X32 FILLER_34_212 ();
 FILLCELL_X32 FILLER_34_244 ();
 FILLCELL_X32 FILLER_34_276 ();
 FILLCELL_X32 FILLER_34_308 ();
 FILLCELL_X32 FILLER_34_340 ();
 FILLCELL_X8 FILLER_34_372 ();
 FILLCELL_X4 FILLER_34_380 ();
 FILLCELL_X2 FILLER_34_384 ();
 FILLCELL_X1 FILLER_34_386 ();
 FILLCELL_X1 FILLER_34_410 ();
 FILLCELL_X1 FILLER_34_415 ();
 FILLCELL_X2 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_3 ();
 FILLCELL_X2 FILLER_35_7 ();
 FILLCELL_X2 FILLER_35_12 ();
 FILLCELL_X1 FILLER_35_14 ();
 FILLCELL_X32 FILLER_35_17 ();
 FILLCELL_X32 FILLER_35_49 ();
 FILLCELL_X32 FILLER_35_81 ();
 FILLCELL_X32 FILLER_35_113 ();
 FILLCELL_X32 FILLER_35_145 ();
 FILLCELL_X32 FILLER_35_177 ();
 FILLCELL_X32 FILLER_35_209 ();
 FILLCELL_X32 FILLER_35_241 ();
 FILLCELL_X32 FILLER_35_273 ();
 FILLCELL_X32 FILLER_35_305 ();
 FILLCELL_X32 FILLER_35_337 ();
 FILLCELL_X8 FILLER_35_369 ();
 FILLCELL_X4 FILLER_35_377 ();
 FILLCELL_X2 FILLER_35_381 ();
 FILLCELL_X1 FILLER_35_383 ();
 FILLCELL_X2 FILLER_35_400 ();
 FILLCELL_X1 FILLER_35_402 ();
 FILLCELL_X1 FILLER_35_412 ();
 FILLCELL_X2 FILLER_35_416 ();
 FILLCELL_X1 FILLER_35_418 ();
 FILLCELL_X1 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_24 ();
 FILLCELL_X32 FILLER_36_56 ();
 FILLCELL_X32 FILLER_36_88 ();
 FILLCELL_X32 FILLER_36_120 ();
 FILLCELL_X32 FILLER_36_152 ();
 FILLCELL_X32 FILLER_36_184 ();
 FILLCELL_X32 FILLER_36_216 ();
 FILLCELL_X32 FILLER_36_248 ();
 FILLCELL_X32 FILLER_36_280 ();
 FILLCELL_X32 FILLER_36_312 ();
 FILLCELL_X32 FILLER_36_344 ();
 FILLCELL_X32 FILLER_36_376 ();
 FILLCELL_X8 FILLER_36_408 ();
 FILLCELL_X2 FILLER_36_416 ();
 FILLCELL_X1 FILLER_36_418 ();
 FILLCELL_X8 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_9 ();
 FILLCELL_X1 FILLER_37_14 ();
 FILLCELL_X4 FILLER_37_18 ();
 FILLCELL_X2 FILLER_37_22 ();
 FILLCELL_X32 FILLER_37_26 ();
 FILLCELL_X32 FILLER_37_58 ();
 FILLCELL_X32 FILLER_37_90 ();
 FILLCELL_X32 FILLER_37_122 ();
 FILLCELL_X32 FILLER_37_154 ();
 FILLCELL_X32 FILLER_37_186 ();
 FILLCELL_X32 FILLER_37_218 ();
 FILLCELL_X32 FILLER_37_250 ();
 FILLCELL_X32 FILLER_37_282 ();
 FILLCELL_X32 FILLER_37_314 ();
 FILLCELL_X32 FILLER_37_346 ();
 FILLCELL_X32 FILLER_37_378 ();
 FILLCELL_X8 FILLER_37_410 ();
 FILLCELL_X1 FILLER_37_418 ();
 FILLCELL_X32 FILLER_38_26 ();
 FILLCELL_X32 FILLER_38_58 ();
 FILLCELL_X32 FILLER_38_90 ();
 FILLCELL_X32 FILLER_38_122 ();
 FILLCELL_X32 FILLER_38_154 ();
 FILLCELL_X32 FILLER_38_186 ();
 FILLCELL_X32 FILLER_38_218 ();
 FILLCELL_X32 FILLER_38_250 ();
 FILLCELL_X32 FILLER_38_282 ();
 FILLCELL_X32 FILLER_38_314 ();
 FILLCELL_X32 FILLER_38_346 ();
 FILLCELL_X32 FILLER_38_378 ();
 FILLCELL_X8 FILLER_38_410 ();
 FILLCELL_X1 FILLER_38_418 ();
 FILLCELL_X1 FILLER_39_4 ();
 FILLCELL_X32 FILLER_39_29 ();
 FILLCELL_X32 FILLER_39_61 ();
 FILLCELL_X32 FILLER_39_93 ();
 FILLCELL_X32 FILLER_39_125 ();
 FILLCELL_X32 FILLER_39_157 ();
 FILLCELL_X32 FILLER_39_189 ();
 FILLCELL_X32 FILLER_39_221 ();
 FILLCELL_X32 FILLER_39_253 ();
 FILLCELL_X32 FILLER_39_285 ();
 FILLCELL_X32 FILLER_39_317 ();
 FILLCELL_X32 FILLER_39_349 ();
 FILLCELL_X32 FILLER_39_381 ();
 FILLCELL_X4 FILLER_39_413 ();
 FILLCELL_X2 FILLER_39_417 ();
 FILLCELL_X4 FILLER_40_1 ();
 FILLCELL_X2 FILLER_40_5 ();
 FILLCELL_X2 FILLER_40_9 ();
 FILLCELL_X32 FILLER_40_27 ();
 FILLCELL_X32 FILLER_40_59 ();
 FILLCELL_X32 FILLER_40_91 ();
 FILLCELL_X32 FILLER_40_123 ();
 FILLCELL_X32 FILLER_40_155 ();
 FILLCELL_X32 FILLER_40_187 ();
 FILLCELL_X32 FILLER_40_219 ();
 FILLCELL_X32 FILLER_40_251 ();
 FILLCELL_X32 FILLER_40_283 ();
 FILLCELL_X32 FILLER_40_315 ();
 FILLCELL_X32 FILLER_40_347 ();
 FILLCELL_X32 FILLER_40_379 ();
 FILLCELL_X8 FILLER_40_411 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X2 FILLER_41_417 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X2 FILLER_42_417 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X2 FILLER_43_417 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X2 FILLER_44_417 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X2 FILLER_45_417 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X2 FILLER_46_417 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X2 FILLER_47_417 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X2 FILLER_48_417 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X2 FILLER_49_417 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X2 FILLER_50_417 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X2 FILLER_51_417 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X2 FILLER_52_417 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X2 FILLER_53_417 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X2 FILLER_54_417 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X16 FILLER_55_161 ();
 FILLCELL_X4 FILLER_55_177 ();
 FILLCELL_X2 FILLER_55_181 ();
 FILLCELL_X32 FILLER_55_186 ();
 FILLCELL_X32 FILLER_55_218 ();
 FILLCELL_X32 FILLER_55_250 ();
 FILLCELL_X32 FILLER_55_282 ();
 FILLCELL_X32 FILLER_55_314 ();
 FILLCELL_X32 FILLER_55_346 ();
 FILLCELL_X32 FILLER_55_378 ();
 FILLCELL_X8 FILLER_55_410 ();
 FILLCELL_X1 FILLER_55_418 ();
endmodule
