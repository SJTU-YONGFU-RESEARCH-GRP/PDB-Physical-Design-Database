module parameterized_fft (busy,
    clk,
    data_ready,
    data_valid_in,
    data_valid_out,
    rst_n,
    start,
    data_in_imag,
    data_in_real,
    data_out_imag,
    data_out_real);
 output busy;
 input clk;
 output data_ready;
 input data_valid_in;
 output data_valid_out;
 input rst_n;
 input start;
 input [15:0] data_in_imag;
 input [15:0] data_in_real;
 output [127:0] data_out_imag;
 output [127:0] data_out_real;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire net9;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire net36;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire net8;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire net10;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire net5;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire net27;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire net7;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire net18;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire net6;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire net414;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire net407;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire net58;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire net64;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire net601;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire net41;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire net49;
 wire _03268_;
 wire _03269_;
 wire net51;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire net43;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire net50;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire net46;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire net534;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire net54;
 wire _03925_;
 wire net531;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire net47;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire net66;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire net55;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire net65;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire net40;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire net62;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire net77;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire net67;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire net34;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire net57;
 wire net52;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire net48;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire net56;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire net619;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire net59;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire net649;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire net648;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire clknet_leaf_0_clk;
 wire net385;
 wire \bit_rev_idx[0] ;
 wire \bit_rev_idx[1] ;
 wire \bit_rev_idx[2] ;
 wire \butterfly_count[0] ;
 wire \butterfly_count[1] ;
 wire \butterfly_count[2] ;
 wire \butterfly_in_group[0] ;
 wire \butterfly_in_group[1] ;
 wire \butterfly_in_group[2] ;
 wire \group[0] ;
 wire \group[1] ;
 wire \group[2] ;
 wire \idx1[0] ;
 wire \idx1[1] ;
 wire \idx1[2] ;
 wire \idx2[0] ;
 wire \idx2[1] ;
 wire \idx2[2] ;
 wire \sample_count[0] ;
 wire \sample_count[1] ;
 wire \sample_count[2] ;
 wire \samples_imag[0][0] ;
 wire \samples_imag[0][10] ;
 wire \samples_imag[0][11] ;
 wire \samples_imag[0][12] ;
 wire \samples_imag[0][13] ;
 wire \samples_imag[0][14] ;
 wire \samples_imag[0][15] ;
 wire \samples_imag[0][1] ;
 wire \samples_imag[0][2] ;
 wire \samples_imag[0][3] ;
 wire \samples_imag[0][4] ;
 wire \samples_imag[0][5] ;
 wire \samples_imag[0][6] ;
 wire \samples_imag[0][7] ;
 wire \samples_imag[0][8] ;
 wire \samples_imag[0][9] ;
 wire \samples_imag[1][0] ;
 wire \samples_imag[1][10] ;
 wire \samples_imag[1][11] ;
 wire \samples_imag[1][12] ;
 wire \samples_imag[1][13] ;
 wire \samples_imag[1][14] ;
 wire \samples_imag[1][15] ;
 wire \samples_imag[1][1] ;
 wire \samples_imag[1][2] ;
 wire \samples_imag[1][3] ;
 wire \samples_imag[1][4] ;
 wire \samples_imag[1][5] ;
 wire \samples_imag[1][6] ;
 wire \samples_imag[1][7] ;
 wire \samples_imag[1][8] ;
 wire \samples_imag[1][9] ;
 wire \samples_imag[2][0] ;
 wire \samples_imag[2][10] ;
 wire \samples_imag[2][11] ;
 wire \samples_imag[2][12] ;
 wire \samples_imag[2][13] ;
 wire \samples_imag[2][14] ;
 wire \samples_imag[2][15] ;
 wire \samples_imag[2][1] ;
 wire \samples_imag[2][2] ;
 wire \samples_imag[2][3] ;
 wire \samples_imag[2][4] ;
 wire \samples_imag[2][5] ;
 wire \samples_imag[2][6] ;
 wire \samples_imag[2][7] ;
 wire \samples_imag[2][8] ;
 wire \samples_imag[2][9] ;
 wire \samples_imag[3][0] ;
 wire \samples_imag[3][10] ;
 wire \samples_imag[3][11] ;
 wire \samples_imag[3][12] ;
 wire \samples_imag[3][13] ;
 wire \samples_imag[3][14] ;
 wire \samples_imag[3][15] ;
 wire \samples_imag[3][1] ;
 wire \samples_imag[3][2] ;
 wire \samples_imag[3][3] ;
 wire \samples_imag[3][4] ;
 wire \samples_imag[3][5] ;
 wire \samples_imag[3][6] ;
 wire \samples_imag[3][7] ;
 wire \samples_imag[3][8] ;
 wire \samples_imag[3][9] ;
 wire \samples_imag[4][0] ;
 wire \samples_imag[4][10] ;
 wire \samples_imag[4][11] ;
 wire \samples_imag[4][12] ;
 wire \samples_imag[4][13] ;
 wire \samples_imag[4][14] ;
 wire \samples_imag[4][15] ;
 wire \samples_imag[4][1] ;
 wire \samples_imag[4][2] ;
 wire \samples_imag[4][3] ;
 wire \samples_imag[4][4] ;
 wire \samples_imag[4][5] ;
 wire \samples_imag[4][6] ;
 wire \samples_imag[4][7] ;
 wire \samples_imag[4][8] ;
 wire \samples_imag[4][9] ;
 wire \samples_imag[5][0] ;
 wire \samples_imag[5][10] ;
 wire \samples_imag[5][11] ;
 wire \samples_imag[5][12] ;
 wire \samples_imag[5][13] ;
 wire \samples_imag[5][14] ;
 wire \samples_imag[5][15] ;
 wire \samples_imag[5][1] ;
 wire \samples_imag[5][2] ;
 wire \samples_imag[5][3] ;
 wire \samples_imag[5][4] ;
 wire \samples_imag[5][5] ;
 wire \samples_imag[5][6] ;
 wire \samples_imag[5][7] ;
 wire \samples_imag[5][8] ;
 wire \samples_imag[5][9] ;
 wire \samples_imag[6][0] ;
 wire \samples_imag[6][10] ;
 wire \samples_imag[6][11] ;
 wire \samples_imag[6][12] ;
 wire \samples_imag[6][13] ;
 wire \samples_imag[6][14] ;
 wire \samples_imag[6][15] ;
 wire \samples_imag[6][1] ;
 wire \samples_imag[6][2] ;
 wire \samples_imag[6][3] ;
 wire \samples_imag[6][4] ;
 wire \samples_imag[6][5] ;
 wire \samples_imag[6][6] ;
 wire \samples_imag[6][7] ;
 wire \samples_imag[6][8] ;
 wire \samples_imag[6][9] ;
 wire \samples_imag[7][0] ;
 wire \samples_imag[7][10] ;
 wire \samples_imag[7][11] ;
 wire \samples_imag[7][12] ;
 wire \samples_imag[7][13] ;
 wire \samples_imag[7][14] ;
 wire \samples_imag[7][15] ;
 wire \samples_imag[7][1] ;
 wire \samples_imag[7][2] ;
 wire \samples_imag[7][3] ;
 wire \samples_imag[7][4] ;
 wire \samples_imag[7][5] ;
 wire \samples_imag[7][6] ;
 wire \samples_imag[7][7] ;
 wire \samples_imag[7][8] ;
 wire \samples_imag[7][9] ;
 wire \samples_real[0][0] ;
 wire \samples_real[0][10] ;
 wire \samples_real[0][11] ;
 wire \samples_real[0][12] ;
 wire \samples_real[0][13] ;
 wire \samples_real[0][14] ;
 wire \samples_real[0][15] ;
 wire \samples_real[0][1] ;
 wire \samples_real[0][2] ;
 wire \samples_real[0][3] ;
 wire \samples_real[0][4] ;
 wire \samples_real[0][5] ;
 wire \samples_real[0][6] ;
 wire \samples_real[0][7] ;
 wire \samples_real[0][8] ;
 wire \samples_real[0][9] ;
 wire \samples_real[1][0] ;
 wire \samples_real[1][10] ;
 wire \samples_real[1][11] ;
 wire \samples_real[1][12] ;
 wire \samples_real[1][13] ;
 wire \samples_real[1][14] ;
 wire \samples_real[1][15] ;
 wire \samples_real[1][1] ;
 wire \samples_real[1][2] ;
 wire \samples_real[1][3] ;
 wire \samples_real[1][4] ;
 wire \samples_real[1][5] ;
 wire \samples_real[1][6] ;
 wire \samples_real[1][7] ;
 wire \samples_real[1][8] ;
 wire \samples_real[1][9] ;
 wire \samples_real[2][0] ;
 wire \samples_real[2][10] ;
 wire \samples_real[2][11] ;
 wire \samples_real[2][12] ;
 wire \samples_real[2][13] ;
 wire \samples_real[2][14] ;
 wire \samples_real[2][15] ;
 wire \samples_real[2][1] ;
 wire \samples_real[2][2] ;
 wire \samples_real[2][3] ;
 wire \samples_real[2][4] ;
 wire \samples_real[2][5] ;
 wire \samples_real[2][6] ;
 wire \samples_real[2][7] ;
 wire \samples_real[2][8] ;
 wire \samples_real[2][9] ;
 wire \samples_real[3][0] ;
 wire \samples_real[3][10] ;
 wire \samples_real[3][11] ;
 wire \samples_real[3][12] ;
 wire \samples_real[3][13] ;
 wire \samples_real[3][14] ;
 wire \samples_real[3][15] ;
 wire \samples_real[3][1] ;
 wire \samples_real[3][2] ;
 wire \samples_real[3][3] ;
 wire \samples_real[3][4] ;
 wire \samples_real[3][5] ;
 wire \samples_real[3][6] ;
 wire \samples_real[3][7] ;
 wire \samples_real[3][8] ;
 wire \samples_real[3][9] ;
 wire \samples_real[4][0] ;
 wire \samples_real[4][10] ;
 wire \samples_real[4][11] ;
 wire \samples_real[4][12] ;
 wire \samples_real[4][13] ;
 wire \samples_real[4][14] ;
 wire \samples_real[4][15] ;
 wire \samples_real[4][1] ;
 wire \samples_real[4][2] ;
 wire \samples_real[4][3] ;
 wire \samples_real[4][4] ;
 wire \samples_real[4][5] ;
 wire \samples_real[4][6] ;
 wire \samples_real[4][7] ;
 wire \samples_real[4][8] ;
 wire \samples_real[4][9] ;
 wire \samples_real[5][0] ;
 wire \samples_real[5][10] ;
 wire \samples_real[5][11] ;
 wire \samples_real[5][12] ;
 wire \samples_real[5][13] ;
 wire \samples_real[5][14] ;
 wire \samples_real[5][15] ;
 wire \samples_real[5][1] ;
 wire \samples_real[5][2] ;
 wire \samples_real[5][3] ;
 wire \samples_real[5][4] ;
 wire \samples_real[5][5] ;
 wire \samples_real[5][6] ;
 wire \samples_real[5][7] ;
 wire \samples_real[5][8] ;
 wire \samples_real[5][9] ;
 wire \samples_real[6][0] ;
 wire \samples_real[6][10] ;
 wire \samples_real[6][11] ;
 wire \samples_real[6][12] ;
 wire \samples_real[6][13] ;
 wire \samples_real[6][14] ;
 wire \samples_real[6][15] ;
 wire \samples_real[6][1] ;
 wire \samples_real[6][2] ;
 wire \samples_real[6][3] ;
 wire \samples_real[6][4] ;
 wire \samples_real[6][5] ;
 wire \samples_real[6][6] ;
 wire \samples_real[6][7] ;
 wire \samples_real[6][8] ;
 wire \samples_real[6][9] ;
 wire \samples_real[7][0] ;
 wire \samples_real[7][10] ;
 wire \samples_real[7][11] ;
 wire \samples_real[7][12] ;
 wire \samples_real[7][13] ;
 wire \samples_real[7][14] ;
 wire \samples_real[7][15] ;
 wire \samples_real[7][1] ;
 wire \samples_real[7][2] ;
 wire \samples_real[7][3] ;
 wire \samples_real[7][4] ;
 wire \samples_real[7][5] ;
 wire \samples_real[7][6] ;
 wire \samples_real[7][7] ;
 wire \samples_real[7][8] ;
 wire \samples_real[7][9] ;
 wire \stage[0] ;
 wire \stage[1] ;
 wire \stage[2] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \temp_imag[0] ;
 wire \temp_real[0] ;
 wire \twiddle_idx[0] ;
 wire \twiddle_idx[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net35;
 wire net37;
 wire net38;
 wire net39;
 wire net42;
 wire net44;
 wire net45;
 wire net60;
 wire net61;
 wire net63;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net408;
 wire net409;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net462;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net603;
 wire net528;
 wire net529;
 wire net530;
 wire net532;
 wire net533;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net602;
 wire net600;
 wire net610;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net646;
 wire net647;
 wire net53;
 wire net410;
 wire net411;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net510;
 wire net512;
 wire net513;
 wire net564;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net611;
 wire net612;
 wire net617;

 sky130_fd_sc_hd__inv_1 _08341_ (.A(net93),
    .Y(_00557_));
 sky130_fd_sc_hd__buf_8 _08342_ (.A(\state[3] ),
    .X(_00558_));
 sky130_fd_sc_hd__buf_6 _08343_ (.A(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__clkbuf_4 _08344_ (.A(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__a21o_1 _08345_ (.A1(\state[0] ),
    .A2(_00557_),
    .B1(_00560_),
    .X(_00004_));
 sky130_fd_sc_hd__buf_4 _08346_ (.A(\stage[2] ),
    .X(_00561_));
 sky130_fd_sc_hd__nor2b_4 _08347_ (.A(_00561_),
    .B_N(_07805_),
    .Y(_07667_));
 sky130_fd_sc_hd__clkinv_8 _08348_ (.A(_07667_),
    .Y(_07106_));
 sky130_fd_sc_hd__buf_6 _08349_ (.A(_00561_),
    .X(_00562_));
 sky130_fd_sc_hd__buf_6 _08350_ (.A(_07809_),
    .X(_00563_));
 sky130_fd_sc_hd__nand2_8 _08351_ (.A(_00562_),
    .B(_00563_),
    .Y(_07166_));
 sky130_fd_sc_hd__inv_1 _08352_ (.A(_07166_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_8 _08353_ (.A(_00562_),
    .B(_07811_),
    .Y(_07153_));
 sky130_fd_sc_hd__inv_1 _08354_ (.A(_07153_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand2_8 _08355_ (.A(_00561_),
    .B(_07805_),
    .Y(_07133_));
 sky130_fd_sc_hd__clkinv_2 _08356_ (.A(_07133_),
    .Y(_07702_));
 sky130_fd_sc_hd__inv_4 _08357_ (.A(_00562_),
    .Y(_07817_));
 sky130_fd_sc_hd__nand2_8 _08358_ (.A(_07817_),
    .B(_00563_),
    .Y(_07112_));
 sky130_fd_sc_hd__inv_1 _08359_ (.A(_07112_),
    .Y(_07710_));
 sky130_fd_sc_hd__nand2_8 _08360_ (.A(_07817_),
    .B(_07811_),
    .Y(_05892_));
 sky130_fd_sc_hd__inv_1 _08361_ (.A(_05892_),
    .Y(_05907_));
 sky130_fd_sc_hd__buf_4 _08362_ (.A(_07824_),
    .X(_00564_));
 sky130_fd_sc_hd__inv_6 _08363_ (.A(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__buf_4 _08364_ (.A(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_4 _08365_ (.A(_00566_),
    .X(_00567_));
 sky130_fd_sc_hd__buf_6 _08366_ (.A(_00567_),
    .X(_00568_));
 sky130_fd_sc_hd__buf_4 _08367_ (.A(_00568_),
    .X(_00569_));
 sky130_fd_sc_hd__clkbuf_16 _08368_ (.A(_00569_),
    .X(_07207_));
 sky130_fd_sc_hd__o21ai_1 _08369_ (.A1(_07805_),
    .A2(_07811_),
    .B1(_00561_),
    .Y(_00570_));
 sky130_fd_sc_hd__clkbuf_2 clone9 (.A(_00810_),
    .X(net9));
 sky130_fd_sc_hd__nor3_2 _08371_ (.A(_07821_),
    .B(_00563_),
    .C(_00564_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_00570_),
    .B(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__clkinv_16 _08373_ (.A(_07706_),
    .Y(_07121_));
 sky130_fd_sc_hd__nor3b_2 _08374_ (.A(\butterfly_count[2] ),
    .B(_07690_),
    .C_N(_07799_),
    .Y(_00574_));
 sky130_fd_sc_hd__o21ai_4 _08375_ (.A1(_00563_),
    .A2(_07811_),
    .B1(_00561_),
    .Y(_00575_));
 sky130_fd_sc_hd__mux2i_1 _08376_ (.A0(_00563_),
    .A1(_07805_),
    .S(_00561_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand4_2 _08377_ (.A(_07121_),
    .B(_00574_),
    .C(_00575_),
    .D(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__o21bai_1 _08378_ (.A1(_07805_),
    .A2(_07811_),
    .B1_N(_00562_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_4 _08379_ (.A(_07108_),
    .B(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__a21oi_4 _08380_ (.A1(_00573_),
    .A2(_00577_),
    .B1(_00579_),
    .Y(_07109_));
 sky130_fd_sc_hd__and4_1 _08381_ (.A(_07817_),
    .B(_07110_),
    .C(_07805_),
    .D(_00572_),
    .X(_07116_));
 sky130_fd_sc_hd__o21a_1 _08382_ (.A1(_07532_),
    .A2(_07531_),
    .B1(_07550_),
    .X(_00580_));
 sky130_fd_sc_hd__o21a_1 _08383_ (.A1(_00580_),
    .A2(_07549_),
    .B1(_07547_),
    .X(_00581_));
 sky130_fd_sc_hd__o21a_1 _08384_ (.A1(_07546_),
    .A2(_00581_),
    .B1(_07544_),
    .X(_00582_));
 sky130_fd_sc_hd__o21a_1 _08385_ (.A1(_07543_),
    .A2(_00582_),
    .B1(_07541_),
    .X(_00583_));
 sky130_fd_sc_hd__o21a_1 _08386_ (.A1(_00583_),
    .A2(_07540_),
    .B1(_07538_),
    .X(_00584_));
 sky130_fd_sc_hd__o21a_1 _08387_ (.A1(_07370_),
    .A2(_07369_),
    .B1(_07368_),
    .X(_00585_));
 sky130_fd_sc_hd__o21a_1 _08388_ (.A1(_07367_),
    .A2(_00585_),
    .B1(_07365_),
    .X(_00586_));
 sky130_fd_sc_hd__o21a_1 _08389_ (.A1(_07364_),
    .A2(_00586_),
    .B1(_07362_),
    .X(_00587_));
 sky130_fd_sc_hd__o21a_1 _08390_ (.A1(_00587_),
    .A2(_07361_),
    .B1(_07359_),
    .X(_00588_));
 sky130_fd_sc_hd__o21a_1 _08391_ (.A1(_07358_),
    .A2(_00588_),
    .B1(_07356_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_4 _08392_ (.A(_00589_),
    .B(_07355_),
    .Y(_00590_));
 sky130_fd_sc_hd__inv_2 _08393_ (.A(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__a21oi_4 _08394_ (.A1(_00591_),
    .A2(_07353_),
    .B1(_07352_),
    .Y(_00592_));
 sky130_fd_sc_hd__buf_6 _08395_ (.A(_07690_),
    .X(_00593_));
 sky130_fd_sc_hd__buf_6 _08396_ (.A(_00593_),
    .X(_00594_));
 sky130_fd_sc_hd__o21ai_4 _08397_ (.A1(_00592_),
    .A2(_00567_),
    .B1(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__buf_4 _08398_ (.A(_00564_),
    .X(_00596_));
 sky130_fd_sc_hd__clkbuf_4 _08399_ (.A(_00596_),
    .X(_00597_));
 sky130_fd_sc_hd__buf_4 _08400_ (.A(_00597_),
    .X(_00598_));
 sky130_fd_sc_hd__buf_4 _08401_ (.A(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__nor2_2 _08402_ (.A(_00599_),
    .B(_00592_),
    .Y(_00600_));
 sky130_fd_sc_hd__o21a_1 _08403_ (.A1(_07250_),
    .A2(_07249_),
    .B1(_07248_),
    .X(_00601_));
 sky130_fd_sc_hd__o21ai_2 _08404_ (.A1(_07247_),
    .A2(_00601_),
    .B1(_07245_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2b_1 _08405_ (.A_N(_07244_),
    .B(_00602_),
    .Y(_00603_));
 sky130_fd_sc_hd__and2_0 _08406_ (.A(_07242_),
    .B(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__o21a_1 _08407_ (.A1(_07241_),
    .A2(_00604_),
    .B1(_07239_),
    .X(_00605_));
 sky130_fd_sc_hd__or3b_4 _08408_ (.A(\butterfly_count[2] ),
    .B(_07690_),
    .C_N(_07799_),
    .X(_00606_));
 sky130_fd_sc_hd__nand3_2 _08409_ (.A(_07172_),
    .B(_07175_),
    .C(_07178_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand4_2 _08410_ (.A(_07169_),
    .B(_07186_),
    .C(_07181_),
    .D(_07184_),
    .Y(_00608_));
 sky130_fd_sc_hd__o31ai_1 _08411_ (.A1(_00606_),
    .A2(_00607_),
    .A3(_00608_),
    .B1(_00596_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3b_1 _08412_ (.A_N(_07169_),
    .B(_07168_),
    .C(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2b_1 _08413_ (.A_N(_00564_),
    .B(_07168_),
    .Y(_00611_));
 sky130_fd_sc_hd__o31ai_4 _08414_ (.A1(_00606_),
    .A2(_00608_),
    .A3(_00607_),
    .B1(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _08415_ (.A(_07169_),
    .B(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__and2_4 _08416_ (.A(_07172_),
    .B(_07175_),
    .X(_00614_));
 sky130_fd_sc_hd__o211ai_4 _08417_ (.A1(_07186_),
    .A2(_07185_),
    .B1(_07184_),
    .C1(_07181_),
    .Y(_00615_));
 sky130_fd_sc_hd__a21oi_2 _08418_ (.A1(_07181_),
    .A2(_07183_),
    .B1(_07180_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_2 _08419_ (.A(_00615_),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__a221o_2 _08420_ (.A1(_07172_),
    .A2(_07174_),
    .B1(_00614_),
    .B2(_07177_),
    .C1(_07171_),
    .X(_00618_));
 sky130_fd_sc_hd__a31oi_4 _08421_ (.A1(_07178_),
    .A2(_00614_),
    .A3(_00617_),
    .B1(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__mux2i_4 _08422_ (.A0(_00610_),
    .A1(_00613_),
    .S(_00619_),
    .Y(_00620_));
 sky130_fd_sc_hd__o31a_1 _08423_ (.A1(_07805_),
    .A2(_00563_),
    .A3(_07811_),
    .B1(_00562_),
    .X(_00621_));
 sky130_fd_sc_hd__nor2_2 _08424_ (.A(_00564_),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__o21a_1 _08425_ (.A1(_07132_),
    .A2(_07131_),
    .B1(_07130_),
    .X(_00623_));
 sky130_fd_sc_hd__o21a_1 _08426_ (.A1(_07129_),
    .A2(_00623_),
    .B1(_07127_),
    .X(_00624_));
 sky130_fd_sc_hd__o21ai_1 _08427_ (.A1(_07126_),
    .A2(_00624_),
    .B1(_07124_),
    .Y(_00625_));
 sky130_fd_sc_hd__or3_1 _08428_ (.A(_07124_),
    .B(_07126_),
    .C(_00624_),
    .X(_00626_));
 sky130_fd_sc_hd__nand4_4 _08429_ (.A(_07123_),
    .B(_00622_),
    .C(_00625_),
    .D(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__and2_0 _08430_ (.A(_00570_),
    .B(_00572_),
    .X(_00628_));
 sky130_fd_sc_hd__o211ai_2 _08431_ (.A1(_07110_),
    .A2(_07106_),
    .B1(_00570_),
    .C1(_00572_),
    .Y(_00629_));
 sky130_fd_sc_hd__nor2_1 _08432_ (.A(_07111_),
    .B(_07110_),
    .Y(_00630_));
 sky130_fd_sc_hd__nor2b_4 _08433_ (.A(_07107_),
    .B_N(_07111_),
    .Y(_00631_));
 sky130_fd_sc_hd__and3b_1 _08434_ (.A_N(_07111_),
    .B(_07110_),
    .C(_07107_),
    .X(_00632_));
 sky130_fd_sc_hd__a311oi_2 _08435_ (.A1(_07108_),
    .A2(_00578_),
    .A3(_00630_),
    .B1(_00632_),
    .C1(_00631_),
    .Y(_00633_));
 sky130_fd_sc_hd__o32ai_4 _08436_ (.A1(_00579_),
    .A2(_00628_),
    .A3(_00577_),
    .B1(_00633_),
    .B2(_00629_),
    .Y(_07113_));
 sky130_fd_sc_hd__o211a_1 _08437_ (.A1(_07120_),
    .A2(_07119_),
    .B1(_07115_),
    .C1(_07118_),
    .X(_00634_));
 sky130_fd_sc_hd__a21o_1 _08438_ (.A1(_07117_),
    .A2(_07115_),
    .B1(_07114_),
    .X(_00635_));
 sky130_fd_sc_hd__o31ai_4 _08439_ (.A1(_07805_),
    .A2(_00563_),
    .A3(_07811_),
    .B1(_00562_),
    .Y(_00636_));
 sky130_fd_sc_hd__o211a_4 _08440_ (.A1(_00634_),
    .A2(_00635_),
    .B1(_00565_),
    .C1(_00636_),
    .X(_00637_));
 sky130_fd_sc_hd__nand3_4 _08441_ (.A(_07118_),
    .B(_07120_),
    .C(_07115_),
    .Y(_00638_));
 sky130_fd_sc_hd__nor4b_4 _08442_ (.A(_00638_),
    .B(_00606_),
    .C(_07702_),
    .D_N(_00575_),
    .Y(_00639_));
 sky130_fd_sc_hd__o21a_1 _08443_ (.A1(_00639_),
    .A2(_00637_),
    .B1(_07121_),
    .X(_00640_));
 sky130_fd_sc_hd__o21a_1 _08444_ (.A1(_07120_),
    .A2(_07119_),
    .B1(_07118_),
    .X(_00641_));
 sky130_fd_sc_hd__nor3_1 _08445_ (.A(_07117_),
    .B(_07115_),
    .C(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__o21a_1 _08446_ (.A1(_07117_),
    .A2(_00641_),
    .B1(_07115_),
    .X(_00643_));
 sky130_fd_sc_hd__o221ai_4 _08447_ (.A1(_00639_),
    .A2(_00637_),
    .B1(_00642_),
    .B2(_00643_),
    .C1(_07121_),
    .Y(_00644_));
 sky130_fd_sc_hd__or3_1 _08448_ (.A(_07129_),
    .B(_07126_),
    .C(_07123_),
    .X(_00645_));
 sky130_fd_sc_hd__or3_1 _08449_ (.A(_07127_),
    .B(_07123_),
    .C(_07126_),
    .X(_00646_));
 sky130_fd_sc_hd__o221a_4 _08450_ (.A1(_07124_),
    .A2(_07123_),
    .B1(_00623_),
    .B2(_00645_),
    .C1(_00646_),
    .X(_00647_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_00622_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__o211ai_4 _08452_ (.A1(_07113_),
    .A2(_00640_),
    .B1(_00644_),
    .C1(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__o2111ai_1 _08453_ (.A1(_07169_),
    .A2(_07168_),
    .B1(_07178_),
    .C1(_07175_),
    .D1(_07172_),
    .Y(_00650_));
 sky130_fd_sc_hd__a211oi_2 _08454_ (.A1(_00615_),
    .A2(_00616_),
    .B1(_00564_),
    .C1(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__a311o_4 _08455_ (.A1(_07169_),
    .A2(_00565_),
    .A3(_00618_),
    .B1(_00612_),
    .C1(_00651_),
    .X(_00652_));
 sky130_fd_sc_hd__a21oi_4 _08456_ (.A1(_00561_),
    .A2(_00563_),
    .B1(_00564_),
    .Y(_00653_));
 sky130_fd_sc_hd__o21a_1 _08457_ (.A1(_07165_),
    .A2(_07164_),
    .B1(_07162_),
    .X(_00654_));
 sky130_fd_sc_hd__or3_1 _08458_ (.A(_07149_),
    .B(_07161_),
    .C(_07164_),
    .X(_00655_));
 sky130_fd_sc_hd__o21a_1 _08459_ (.A1(_07152_),
    .A2(_07151_),
    .B1(_07150_),
    .X(_00656_));
 sky130_fd_sc_hd__o22a_4 _08460_ (.A1(_07161_),
    .A2(_00654_),
    .B1(_00656_),
    .B2(_00655_),
    .X(_00657_));
 sky130_fd_sc_hd__a21oi_2 _08461_ (.A1(_07158_),
    .A2(_07156_),
    .B1(_07155_),
    .Y(_00658_));
 sky130_fd_sc_hd__and2b_2 _08462_ (.A_N(_00658_),
    .B(_00653_),
    .X(_00659_));
 sky130_fd_sc_hd__a41o_4 _08463_ (.A1(_00657_),
    .A2(_07159_),
    .A3(_00653_),
    .A4(_07156_),
    .B1(_00659_),
    .X(_00660_));
 sky130_fd_sc_hd__a41o_1 clone36 (.A1(_00657_),
    .A2(_07159_),
    .A3(_00653_),
    .A4(_07156_),
    .B1(_00659_),
    .X(net36));
 sky130_fd_sc_hd__o21a_1 _08465_ (.A1(_07141_),
    .A2(_07142_),
    .B1(_07139_),
    .X(_00662_));
 sky130_fd_sc_hd__o21a_1 _08466_ (.A1(_07147_),
    .A2(_07146_),
    .B1(_07145_),
    .X(_00663_));
 sky130_fd_sc_hd__or3_1 _08467_ (.A(_07138_),
    .B(_07144_),
    .C(_07141_),
    .X(_00664_));
 sky130_fd_sc_hd__o22ai_2 _08468_ (.A1(_07138_),
    .A2(_00662_),
    .B1(_00664_),
    .B2(_00663_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand3_1 _08469_ (.A(_07136_),
    .B(_00565_),
    .C(_00575_),
    .Y(_00666_));
 sky130_fd_sc_hd__and4_1 _08470_ (.A(_07147_),
    .B(_07136_),
    .C(_07139_),
    .D(_07142_),
    .X(_00667_));
 sky130_fd_sc_hd__nand4_1 _08471_ (.A(_07145_),
    .B(_00574_),
    .C(_00575_),
    .D(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand3_1 _08472_ (.A(_07135_),
    .B(_00565_),
    .C(_00575_),
    .Y(_00669_));
 sky130_fd_sc_hd__o211ai_2 _08473_ (.A1(_00666_),
    .A2(_00665_),
    .B1(_00668_),
    .C1(_00669_),
    .Y(_00670_));
 sky130_fd_sc_hd__nor3_1 _08474_ (.A(_00652_),
    .B(net36),
    .C(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__a21boi_4 _08475_ (.A1(_00627_),
    .A2(_00649_),
    .B1_N(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__a41oi_4 _08476_ (.A1(_07156_),
    .A2(_07159_),
    .A3(_00653_),
    .A4(_00657_),
    .B1(_00659_),
    .Y(_00673_));
 sky130_fd_sc_hd__xnor2_1 _08477_ (.A(_07136_),
    .B(_00665_),
    .Y(_00674_));
 sky130_fd_sc_hd__buf_6 _08478_ (.A(_00670_),
    .X(_00675_));
 sky130_fd_sc_hd__nand3_2 _08479_ (.A(_00673_),
    .B(_00674_),
    .C(net6),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _08480_ (.A(_07155_),
    .B(_00653_),
    .Y(_00677_));
 sky130_fd_sc_hd__nor2_1 _08481_ (.A(_07156_),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__and3_1 _08482_ (.A(_07156_),
    .B(_07155_),
    .C(_00653_),
    .X(_00679_));
 sky130_fd_sc_hd__a21oi_2 _08483_ (.A1(_00657_),
    .A2(_07159_),
    .B1(_07158_),
    .Y(_00680_));
 sky130_fd_sc_hd__mux2i_4 _08484_ (.A0(_00678_),
    .A1(_00679_),
    .S(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21oi_4 _08485_ (.A1(_00676_),
    .A2(_00681_),
    .B1(_00652_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor3_4 _08486_ (.A(_00620_),
    .B(_00672_),
    .C(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__o211ai_4 _08487_ (.A1(_00634_),
    .A2(_00635_),
    .B1(_00565_),
    .C1(_00636_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand4_1 _08488_ (.A(_07121_),
    .B(_07133_),
    .C(_00574_),
    .D(_00575_),
    .Y(_00685_));
 sky130_fd_sc_hd__o221ai_4 _08489_ (.A1(_07706_),
    .A2(_00684_),
    .B1(_00638_),
    .B2(_00685_),
    .C1(_07116_),
    .Y(_00686_));
 sky130_fd_sc_hd__nor3_1 _08490_ (.A(_07118_),
    .B(_07120_),
    .C(_07119_),
    .Y(_00687_));
 sky130_fd_sc_hd__nor3_1 _08491_ (.A(_07706_),
    .B(_00641_),
    .C(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__o21ai_2 _08492_ (.A1(_00637_),
    .A2(_00639_),
    .B1(_00688_),
    .Y(_00689_));
 sky130_fd_sc_hd__a221oi_2 _08493_ (.A1(_00622_),
    .A2(_00647_),
    .B1(_00686_),
    .B2(_00689_),
    .C1(_00675_),
    .Y(_00690_));
 sky130_fd_sc_hd__a21oi_1 _08494_ (.A1(_07124_),
    .A2(_07126_),
    .B1(_07123_),
    .Y(_00691_));
 sky130_fd_sc_hd__nor3_1 _08495_ (.A(_07127_),
    .B(_07129_),
    .C(_00623_),
    .Y(_00692_));
 sky130_fd_sc_hd__or4b_1 _08496_ (.A(_00624_),
    .B(_00691_),
    .C(_00692_),
    .D_N(_00622_),
    .X(_00693_));
 sky130_fd_sc_hd__or2_0 _08497_ (.A(_07141_),
    .B(_07144_),
    .X(_00694_));
 sky130_fd_sc_hd__o22ai_1 _08498_ (.A1(_07142_),
    .A2(_07141_),
    .B1(_00663_),
    .B2(_00694_),
    .Y(_00695_));
 sky130_fd_sc_hd__xor2_1 _08499_ (.A(_07139_),
    .B(_00695_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2i_4 _08500_ (.A0(_00693_),
    .A1(_00696_),
    .S(net6),
    .Y(_00697_));
 sky130_fd_sc_hd__buf_6 _08501_ (.A(_00652_),
    .X(_00698_));
 sky130_fd_sc_hd__o211ai_2 _08502_ (.A1(_07206_),
    .A2(_07205_),
    .B1(_07204_),
    .C1(_07201_),
    .Y(_00699_));
 sky130_fd_sc_hd__a21oi_2 _08503_ (.A1(_07201_),
    .A2(_07203_),
    .B1(_07200_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand4_4 _08504_ (.A(_07195_),
    .B(_07192_),
    .C(_07198_),
    .D(_07189_),
    .Y(_00701_));
 sky130_fd_sc_hd__a21o_1 _08505_ (.A1(_00699_),
    .A2(_00700_),
    .B1(_00701_),
    .X(_00702_));
 sky130_fd_sc_hd__nand3_1 _08506_ (.A(_07189_),
    .B(_07192_),
    .C(_07194_),
    .Y(_00703_));
 sky130_fd_sc_hd__a21oi_2 _08507_ (.A1(_07189_),
    .A2(_07191_),
    .B1(_07188_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand4_4 _08508_ (.A(_07189_),
    .B(_07192_),
    .C(_07195_),
    .D(_07197_),
    .Y(_00705_));
 sky130_fd_sc_hd__and3_4 _08509_ (.A(_00703_),
    .B(_00704_),
    .C(_00705_),
    .X(_00706_));
 sky130_fd_sc_hd__a21oi_4 _08510_ (.A1(_00702_),
    .A2(_00706_),
    .B1(_07690_),
    .Y(_00707_));
 sky130_fd_sc_hd__nor3_1 _08511_ (.A(net26),
    .B(net36),
    .C(_00707_),
    .Y(_00708_));
 sky130_fd_sc_hd__o21ai_1 _08512_ (.A1(_00690_),
    .A2(_00697_),
    .B1(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__a311oi_4 _08513_ (.A1(_00618_),
    .A2(_00565_),
    .A3(_07169_),
    .B1(_00612_),
    .C1(_00651_),
    .Y(_00710_));
 sky130_fd_sc_hd__and2_0 _08514_ (.A(_07175_),
    .B(_07177_),
    .X(_00711_));
 sky130_fd_sc_hd__nand2_1 _08515_ (.A(_07175_),
    .B(_07178_),
    .Y(_00712_));
 sky130_fd_sc_hd__a21oi_1 _08516_ (.A1(_00615_),
    .A2(_00616_),
    .B1(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__o31a_1 _08517_ (.A1(_07174_),
    .A2(_00711_),
    .A3(_00713_),
    .B1(_07172_),
    .X(_00714_));
 sky130_fd_sc_hd__nor4_1 _08518_ (.A(_07172_),
    .B(_07174_),
    .C(_00711_),
    .D(_00713_),
    .Y(_00715_));
 sky130_fd_sc_hd__nor3_2 _08519_ (.A(_00710_),
    .B(_00714_),
    .C(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__xor2_1 _08520_ (.A(_07159_),
    .B(_00657_),
    .X(_00717_));
 sky130_fd_sc_hd__and3_1 _08521_ (.A(_00710_),
    .B(net36),
    .C(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__nand3_1 _08522_ (.A(_07192_),
    .B(_07195_),
    .C(_07198_),
    .Y(_00719_));
 sky130_fd_sc_hd__a21oi_1 _08523_ (.A1(_00699_),
    .A2(_00700_),
    .B1(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__a21oi_1 _08524_ (.A1(_07195_),
    .A2(_07197_),
    .B1(_07194_),
    .Y(_00721_));
 sky130_fd_sc_hd__nor2b_1 _08525_ (.A(_00721_),
    .B_N(_07192_),
    .Y(_00722_));
 sky130_fd_sc_hd__o31a_1 _08526_ (.A1(_07191_),
    .A2(_00720_),
    .A3(_00722_),
    .B1(_07189_),
    .X(_00723_));
 sky130_fd_sc_hd__nor4_1 _08527_ (.A(_07189_),
    .B(_07191_),
    .C(_00720_),
    .D(_00722_),
    .Y(_00724_));
 sky130_fd_sc_hd__o21ai_0 _08528_ (.A1(_00723_),
    .A2(_00724_),
    .B1(_00707_),
    .Y(_00725_));
 sky130_fd_sc_hd__o31ai_1 _08529_ (.A1(_00707_),
    .A2(_00716_),
    .A3(_00718_),
    .B1(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__o21ai_2 _08530_ (.A1(_07230_),
    .A2(_07229_),
    .B1(_07228_),
    .Y(_00727_));
 sky130_fd_sc_hd__nor2_1 _08531_ (.A(_07224_),
    .B(_07227_),
    .Y(_00728_));
 sky130_fd_sc_hd__nor2_2 _08532_ (.A(_07225_),
    .B(_07224_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand3_1 _08533_ (.A(_07216_),
    .B(_07219_),
    .C(_07222_),
    .Y(_00730_));
 sky130_fd_sc_hd__a211oi_4 _08534_ (.A1(_00727_),
    .A2(_00728_),
    .B1(_00729_),
    .C1(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__a21o_1 _08535_ (.A1(_07219_),
    .A2(_07221_),
    .B1(_07218_),
    .X(_00732_));
 sky130_fd_sc_hd__a21o_1 _08536_ (.A1(_00732_),
    .A2(_07216_),
    .B1(_07215_),
    .X(_00733_));
 sky130_fd_sc_hd__o21ai_0 _08537_ (.A1(_07213_),
    .A2(_07212_),
    .B1(_07210_),
    .Y(_00734_));
 sky130_fd_sc_hd__or2b_1 _08538_ (.A(_07209_),
    .B_N(_00734_),
    .X(_00735_));
 sky130_fd_sc_hd__o41ai_4 _08539_ (.A1(_07209_),
    .A2(_07212_),
    .A3(_00733_),
    .A4(_00731_),
    .B1(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__a21boi_1 _08540_ (.A1(_00709_),
    .A2(_00726_),
    .B1_N(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__mux2_2 _08541_ (.A0(_00610_),
    .A1(_00613_),
    .S(_00619_),
    .X(_00738_));
 sky130_fd_sc_hd__or2_4 _08542_ (.A(_00670_),
    .B(_00660_),
    .X(_00739_));
 sky130_fd_sc_hd__a211o_2 _08543_ (.A1(_00627_),
    .A2(_00649_),
    .B1(_00739_),
    .C1(_00698_),
    .X(_00740_));
 sky130_fd_sc_hd__a21o_1 _08544_ (.A1(_00676_),
    .A2(_00681_),
    .B1(_00698_),
    .X(_00741_));
 sky130_fd_sc_hd__and4_1 _08545_ (.A(_07213_),
    .B(_07216_),
    .C(_07219_),
    .D(_07222_),
    .X(_00742_));
 sky130_fd_sc_hd__a21oi_2 _08546_ (.A1(_00727_),
    .A2(_00728_),
    .B1(_00729_),
    .Y(_00743_));
 sky130_fd_sc_hd__a221oi_1 _08547_ (.A1(_07213_),
    .A2(_00733_),
    .B1(_00742_),
    .B2(_00743_),
    .C1(_07212_),
    .Y(_00744_));
 sky130_fd_sc_hd__xor2_1 _08548_ (.A(_07210_),
    .B(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__clkinv_8 _08549_ (.A(_07690_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_2 _08550_ (.A1(_00702_),
    .A2(_00706_),
    .B1(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__nor2_4 _08551_ (.A(_07690_),
    .B(_00596_),
    .Y(_00748_));
 sky130_fd_sc_hd__and3_1 _08552_ (.A(_00702_),
    .B(_00706_),
    .C(_00748_),
    .X(_00749_));
 sky130_fd_sc_hd__or2_1 _08553_ (.A(_00747_),
    .B(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__o21a_1 _08554_ (.A1(_00747_),
    .A2(_00749_),
    .B1(_00736_),
    .X(_00751_));
 sky130_fd_sc_hd__nor2_1 _08555_ (.A(_00723_),
    .B(_00724_),
    .Y(_00752_));
 sky130_fd_sc_hd__a2bb2oi_1 _08556_ (.A1_N(_00745_),
    .A2_N(_00750_),
    .B1(_00751_),
    .B2(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__a31oi_2 _08557_ (.A1(_00738_),
    .A2(_00740_),
    .A3(_00741_),
    .B1(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__nor2_1 _08558_ (.A(_00736_),
    .B(_00745_),
    .Y(_00755_));
 sky130_fd_sc_hd__a211oi_4 _08559_ (.A1(_00683_),
    .A2(_00737_),
    .B1(_00754_),
    .C1(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__and4_4 _08560_ (.A(_00603_),
    .B(_07236_),
    .C(_07239_),
    .D(_07242_),
    .X(_00757_));
 sky130_fd_sc_hd__nand3_1 _08561_ (.A(_07236_),
    .B(_07239_),
    .C(_07241_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand2_1 _08562_ (.A(_07236_),
    .B(_07238_),
    .Y(_00759_));
 sky130_fd_sc_hd__nand2_1 _08563_ (.A(_00758_),
    .B(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__or3_4 _08564_ (.A(_07235_),
    .B(_00760_),
    .C(_00757_),
    .X(_00761_));
 sky130_fd_sc_hd__a21oi_4 _08565_ (.A1(_00761_),
    .A2(_07233_),
    .B1(_07232_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_2 _08566_ (.A(_00596_),
    .B(_00762_),
    .Y(_00763_));
 sky130_fd_sc_hd__o21ai_2 _08567_ (.A1(_00565_),
    .A2(_00762_),
    .B1(_07690_),
    .Y(_00764_));
 sky130_fd_sc_hd__nor3_4 _08568_ (.A(_07706_),
    .B(_07120_),
    .C(_00684_),
    .Y(_07128_));
 sky130_fd_sc_hd__nor3_1 _08569_ (.A(_07132_),
    .B(_07130_),
    .C(_07131_),
    .Y(_00765_));
 sky130_fd_sc_hd__nor4_1 _08570_ (.A(_00564_),
    .B(_00621_),
    .C(_00623_),
    .D(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__mux2i_4 _08571_ (.A0(_07128_),
    .A1(_00766_),
    .S(_00647_),
    .Y(_00767_));
 sky130_fd_sc_hd__o21ai_1 _08572_ (.A1(_07149_),
    .A2(_00656_),
    .B1(_07165_),
    .Y(_00768_));
 sky130_fd_sc_hd__or2b_1 _08573_ (.A(_07164_),
    .B_N(_00768_),
    .X(_00769_));
 sky130_fd_sc_hd__xnor2_1 _08574_ (.A(_07162_),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__nor2_1 _08575_ (.A(_07144_),
    .B(_00663_),
    .Y(_00771_));
 sky130_fd_sc_hd__xnor2_1 _08576_ (.A(_07142_),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand3_1 _08577_ (.A(_00673_),
    .B(net6),
    .C(_00772_),
    .Y(_00773_));
 sky130_fd_sc_hd__o221ai_4 _08578_ (.A1(_00767_),
    .A2(_00739_),
    .B1(_00770_),
    .B2(_00673_),
    .C1(_00773_),
    .Y(_07173_));
 sky130_fd_sc_hd__a211oi_1 _08579_ (.A1(_07178_),
    .A2(_00617_),
    .B1(_07177_),
    .C1(_07175_),
    .Y(_00774_));
 sky130_fd_sc_hd__o31a_1 _08580_ (.A1(_00711_),
    .A2(_00713_),
    .A3(_00774_),
    .B1(_00652_),
    .X(_00775_));
 sky130_fd_sc_hd__nor2_1 _08581_ (.A(_00707_),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__a21oi_4 _08582_ (.A1(_00699_),
    .A2(_00700_),
    .B1(_00701_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand3_2 _08583_ (.A(_00703_),
    .B(_00704_),
    .C(_00705_),
    .Y(_00778_));
 sky130_fd_sc_hd__o21ai_4 _08584_ (.A1(_00778_),
    .A2(_00777_),
    .B1(_00746_),
    .Y(_00779_));
 sky130_fd_sc_hd__o211a_1 _08585_ (.A1(_07206_),
    .A2(_07205_),
    .B1(_07204_),
    .C1(_07201_),
    .X(_00780_));
 sky130_fd_sc_hd__a21o_1 _08586_ (.A1(_07201_),
    .A2(_07203_),
    .B1(_07200_),
    .X(_00781_));
 sky130_fd_sc_hd__o21ai_0 _08587_ (.A1(_00780_),
    .A2(_00781_),
    .B1(_07198_),
    .Y(_00782_));
 sky130_fd_sc_hd__nor3_1 _08588_ (.A(_07192_),
    .B(_07194_),
    .C(_07197_),
    .Y(_00783_));
 sky130_fd_sc_hd__a211oi_2 _08589_ (.A1(_00782_),
    .A2(_00783_),
    .B1(_00722_),
    .C1(_00720_),
    .Y(_00784_));
 sky130_fd_sc_hd__or3_1 _08590_ (.A(_07192_),
    .B(_07195_),
    .C(_07194_),
    .X(_00785_));
 sky130_fd_sc_hd__nand2_2 _08591_ (.A(_00784_),
    .B(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__nor2_2 _08592_ (.A(_00779_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__o32ai_4 _08593_ (.A1(net26),
    .A2(_00707_),
    .A3(_07173_),
    .B1(_00776_),
    .B2(_00787_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor2_1 _08594_ (.A(_00731_),
    .B(_00733_),
    .Y(_00789_));
 sky130_fd_sc_hd__xnor2_2 _08595_ (.A(_07213_),
    .B(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__o211ai_1 _08596_ (.A1(_00565_),
    .A2(_00747_),
    .B1(_00784_),
    .C1(_00785_),
    .Y(_00791_));
 sky130_fd_sc_hd__a2bb2oi_1 _08597_ (.A1_N(_00750_),
    .A2_N(_00790_),
    .B1(_00791_),
    .B2(_00751_),
    .Y(_00792_));
 sky130_fd_sc_hd__a31oi_2 _08598_ (.A1(_00738_),
    .A2(_00740_),
    .A3(_00741_),
    .B1(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_1 _08599_ (.A(_00736_),
    .B(_00790_),
    .Y(_00794_));
 sky130_fd_sc_hd__a311oi_4 _08600_ (.A1(_00736_),
    .A2(_00683_),
    .A3(_00788_),
    .B1(_00793_),
    .C1(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__mux2i_4 _08601_ (.A0(_00763_),
    .A1(_00764_),
    .S(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_2 _08602_ (.A(_00738_),
    .B(_00740_),
    .C(_00741_),
    .Y(_00797_));
 sky130_fd_sc_hd__a2111oi_0 _08603_ (.A1(_00627_),
    .A2(_00649_),
    .B1(_00739_),
    .C1(_00786_),
    .D1(net26),
    .Y(_00798_));
 sky130_fd_sc_hd__a211oi_1 _08604_ (.A1(_00676_),
    .A2(_00681_),
    .B1(_00786_),
    .C1(net26),
    .Y(_00799_));
 sky130_fd_sc_hd__nor2_1 _08605_ (.A(_00738_),
    .B(_00786_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor4_1 _08606_ (.A(_00596_),
    .B(_00798_),
    .C(_00799_),
    .D(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__o21ai_0 _08607_ (.A1(_00797_),
    .A2(_00788_),
    .B1(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor2_1 _08608_ (.A(_00736_),
    .B(_00750_),
    .Y(_00803_));
 sky130_fd_sc_hd__o31a_1 _08609_ (.A1(_00620_),
    .A2(_00672_),
    .A3(_00682_),
    .B1(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__buf_4 _08610_ (.A(_00804_),
    .X(_00805_));
 sky130_fd_sc_hd__a31oi_1 _08611_ (.A1(_00596_),
    .A2(_00683_),
    .A3(_00787_),
    .B1(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__a21o_1 _08612_ (.A1(_00738_),
    .A2(net26),
    .B1(_00750_),
    .X(_00807_));
 sky130_fd_sc_hd__nand4_1 _08613_ (.A(_00738_),
    .B(_00736_),
    .C(_00676_),
    .D(_00681_),
    .Y(_00808_));
 sky130_fd_sc_hd__a21oi_1 _08614_ (.A1(_00627_),
    .A2(_00649_),
    .B1(_00739_),
    .Y(_00809_));
 sky130_fd_sc_hd__o2bb2ai_4 _08615_ (.A1_N(_00736_),
    .A2_N(_00807_),
    .B1(_00809_),
    .B2(_00808_),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_1 _08616_ (.A(\butterfly_count[2] ),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_4 _08617_ (.A(_00811_),
    .B(_07799_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand4_1 _08618_ (.A(_07242_),
    .B(_07236_),
    .C(_07239_),
    .D(_07245_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand3_1 _08619_ (.A(_07248_),
    .B(_07250_),
    .C(_07233_),
    .Y(_00814_));
 sky130_fd_sc_hd__nor3_2 _08620_ (.A(_00812_),
    .B(_00813_),
    .C(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__a21oi_1 _08621_ (.A1(_00810_),
    .A2(_00815_),
    .B1(_00805_),
    .Y(_00816_));
 sky130_fd_sc_hd__a21o_2 _08622_ (.A1(_00802_),
    .A2(_00806_),
    .B1(_00816_),
    .X(_00817_));
 sky130_fd_sc_hd__and3_4 _08623_ (.A(_00756_),
    .B(_00817_),
    .C(_00796_),
    .X(_00818_));
 sky130_fd_sc_hd__buf_8 _08624_ (.A(_00818_),
    .X(_00819_));
 sky130_fd_sc_hd__buf_8 _08625_ (.A(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__nor3_1 _08626_ (.A(_07239_),
    .B(_07241_),
    .C(_00604_),
    .Y(_00821_));
 sky130_fd_sc_hd__buf_6 _08627_ (.A(_00810_),
    .X(_00822_));
 sky130_fd_sc_hd__xnor2_1 _08628_ (.A(_07222_),
    .B(_00743_),
    .Y(_00823_));
 sky130_fd_sc_hd__o31ai_2 _08629_ (.A1(_00620_),
    .A2(_00672_),
    .A3(_00682_),
    .B1(_00565_),
    .Y(_00824_));
 sky130_fd_sc_hd__o21ai_2 _08630_ (.A1(_00797_),
    .A2(_00779_),
    .B1(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__o21a_1 _08631_ (.A1(_07206_),
    .A2(_07205_),
    .B1(_07204_),
    .X(_00826_));
 sky130_fd_sc_hd__nor2_1 _08632_ (.A(_07203_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__xor2_1 _08633_ (.A(_07201_),
    .B(_00827_),
    .X(_00828_));
 sky130_fd_sc_hd__o21a_1 _08634_ (.A1(_07186_),
    .A2(_07185_),
    .B1(_07184_),
    .X(_00829_));
 sky130_fd_sc_hd__nor3_1 _08635_ (.A(_07186_),
    .B(_07184_),
    .C(_07185_),
    .Y(_00830_));
 sky130_fd_sc_hd__nor2_1 _08636_ (.A(_07152_),
    .B(_00673_),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_1 _08637_ (.A(_00710_),
    .B(_07182_),
    .Y(_00831_));
 sky130_fd_sc_hd__o31ai_1 _08638_ (.A1(_00829_),
    .A2(_00710_),
    .A3(_00830_),
    .B1(_00831_),
    .Y(_07199_));
 sky130_fd_sc_hd__nor2_1 _08639_ (.A(_00825_),
    .B(_07199_),
    .Y(_00832_));
 sky130_fd_sc_hd__a21oi_1 _08640_ (.A1(_00825_),
    .A2(_00828_),
    .B1(_00832_),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_1 _08641_ (.A(_00822_),
    .B(_07220_),
    .Y(_00833_));
 sky130_fd_sc_hd__o21ai_1 _08642_ (.A1(_00822_),
    .A2(_00823_),
    .B1(_00833_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_2 _08643_ (.A(net30),
    .B(_07237_),
    .Y(_00834_));
 sky130_fd_sc_hd__o31ai_4 _08644_ (.A1(_00605_),
    .A2(_00820_),
    .A3(_00821_),
    .B1(_00834_),
    .Y(_07254_));
 sky130_fd_sc_hd__clkbuf_2 clone8 (.A(_02255_),
    .X(net8));
 sky130_fd_sc_hd__a21o_1 _08646_ (.A1(_07259_),
    .A2(_07269_),
    .B1(_07258_),
    .X(_00836_));
 sky130_fd_sc_hd__nor2_1 _08647_ (.A(_07247_),
    .B(_00601_),
    .Y(_00837_));
 sky130_fd_sc_hd__xnor2_1 _08648_ (.A(_07245_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__o21a_1 _08649_ (.A1(_07230_),
    .A2(_07229_),
    .B1(_07228_),
    .X(_00839_));
 sky130_fd_sc_hd__nor3_1 _08650_ (.A(_07228_),
    .B(_07230_),
    .C(_07229_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_1 _08651_ (.A(_00839_),
    .B(_00840_),
    .Y(_00841_));
 sky130_fd_sc_hd__a31oi_2 _08652_ (.A1(_00738_),
    .A2(_00740_),
    .A3(_00741_),
    .B1(_00596_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor4_4 _08653_ (.A(_00620_),
    .B(_00672_),
    .C(_00779_),
    .D(_00682_),
    .Y(_00843_));
 sky130_fd_sc_hd__nor2_4 _08654_ (.A(_00843_),
    .B(_00842_),
    .Y(_00844_));
 sky130_fd_sc_hd__nor2_1 _08655_ (.A(_07206_),
    .B(_00844_),
    .Y(_07226_));
 sky130_fd_sc_hd__mux2_4 _08656_ (.A0(_00841_),
    .A1(_07226_),
    .S(_00822_),
    .X(_07243_));
 sky130_fd_sc_hd__mux2_4 _08657_ (.A0(_00838_),
    .A1(_07243_),
    .S(_00820_),
    .X(_07268_));
 sky130_fd_sc_hd__xor2_1 _08658_ (.A(_07821_),
    .B(_07268_),
    .X(_00845_));
 sky130_fd_sc_hd__o21a_1 _08659_ (.A1(_07267_),
    .A2(_07266_),
    .B1(_07265_),
    .X(_00846_));
 sky130_fd_sc_hd__o21ai_4 _08660_ (.A1(_07264_),
    .A2(_00846_),
    .B1(_07262_),
    .Y(_00847_));
 sky130_fd_sc_hd__nand2b_1 _08661_ (.A_N(_07261_),
    .B(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand2_1 _08662_ (.A(_07259_),
    .B(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__nor2_1 _08663_ (.A(_00845_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__o21a_1 _08664_ (.A1(_07269_),
    .A2(_00848_),
    .B1(_07259_),
    .X(_00851_));
 sky130_fd_sc_hd__o21ai_0 _08665_ (.A1(_07258_),
    .A2(_00851_),
    .B1(_07256_),
    .Y(_00852_));
 sky130_fd_sc_hd__nor3b_1 _08666_ (.A(_07258_),
    .B(_07269_),
    .C_N(_00845_),
    .Y(_00853_));
 sky130_fd_sc_hd__o32a_1 _08667_ (.A1(_07256_),
    .A2(_00836_),
    .A3(_00850_),
    .B1(_00852_),
    .B2(_00853_),
    .X(_00854_));
 sky130_fd_sc_hd__buf_6 _08668_ (.A(_07253_),
    .X(_00855_));
 sky130_fd_sc_hd__nor2_1 _08669_ (.A(_00855_),
    .B(_07252_),
    .Y(_00856_));
 sky130_fd_sc_hd__nor3_1 _08670_ (.A(_07235_),
    .B(_00757_),
    .C(_00760_),
    .Y(_00857_));
 sky130_fd_sc_hd__xnor2_2 _08671_ (.A(_07233_),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__or3_1 _08672_ (.A(_00597_),
    .B(_00856_),
    .C(_00858_),
    .X(_00859_));
 sky130_fd_sc_hd__nand3b_1 _08673_ (.A_N(_00856_),
    .B(_00858_),
    .C(_00597_),
    .Y(_00860_));
 sky130_fd_sc_hd__a21o_1 _08674_ (.A1(_00859_),
    .A2(_00860_),
    .B1(net31),
    .X(_00861_));
 sky130_fd_sc_hd__a21o_1 _08675_ (.A1(_07222_),
    .A2(_00743_),
    .B1(_07221_),
    .X(_00862_));
 sky130_fd_sc_hd__a21oi_1 _08676_ (.A1(_07219_),
    .A2(_00862_),
    .B1(_07218_),
    .Y(_00863_));
 sky130_fd_sc_hd__xnor2_1 _08677_ (.A(_07216_),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _08678_ (.A(net9),
    .B(_00864_),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_1 _08679_ (.A(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__a21boi_2 _08680_ (.A1(_00699_),
    .A2(_00700_),
    .B1_N(_07198_),
    .Y(_00867_));
 sky130_fd_sc_hd__nor2_1 _08681_ (.A(_07197_),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__xnor2_2 _08682_ (.A(_07195_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__nand3b_4 _08683_ (.A_N(_07132_),
    .B(_00622_),
    .C(_00647_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor3_1 _08684_ (.A(_07147_),
    .B(_07145_),
    .C(_07146_),
    .Y(_00871_));
 sky130_fd_sc_hd__or2_0 _08685_ (.A(_00663_),
    .B(_00871_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2i_4 _08686_ (.A0(_00870_),
    .A1(_00872_),
    .S(_00675_),
    .Y(_07163_));
 sky130_fd_sc_hd__xnor2_1 _08687_ (.A(_07178_),
    .B(_00617_),
    .Y(_00873_));
 sky130_fd_sc_hd__nor2_1 _08688_ (.A(_00873_),
    .B(_00710_),
    .Y(_00874_));
 sky130_fd_sc_hd__or3_1 _08689_ (.A(_07165_),
    .B(_07149_),
    .C(_00656_),
    .X(_00875_));
 sky130_fd_sc_hd__nand2_1 _08690_ (.A(_00768_),
    .B(_00875_),
    .Y(_00876_));
 sky130_fd_sc_hd__nor3_2 _08691_ (.A(_00698_),
    .B(_00673_),
    .C(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__a311o_1 _08692_ (.A1(_00710_),
    .A2(_00673_),
    .A3(_07163_),
    .B1(_00877_),
    .C1(_00874_),
    .X(_07193_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_00593_),
    .B(_07193_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _08694_ (.A(_00747_),
    .B(_00869_),
    .Y(_00879_));
 sky130_fd_sc_hd__mux2i_2 _08695_ (.A0(_00878_),
    .A1(_00879_),
    .S(_00797_),
    .Y(_00880_));
 sky130_fd_sc_hd__nor2_1 _08696_ (.A(_00777_),
    .B(_00778_),
    .Y(_00881_));
 sky130_fd_sc_hd__and3_1 _08697_ (.A(_00881_),
    .B(_00824_),
    .C(_07193_),
    .X(_00882_));
 sky130_fd_sc_hd__inv_2 _08698_ (.A(_00822_),
    .Y(_00883_));
 sky130_fd_sc_hd__a2111o_1 _08699_ (.A1(_00869_),
    .A2(_00825_),
    .B1(_00880_),
    .C1(_00882_),
    .D1(_00883_),
    .X(_00884_));
 sky130_fd_sc_hd__a211oi_1 _08700_ (.A1(_00866_),
    .A2(_00884_),
    .B1(_00597_),
    .C1(_00856_),
    .Y(_00885_));
 sky130_fd_sc_hd__nor4b_1 _08701_ (.A(_00566_),
    .B(_00856_),
    .C(_00865_),
    .D_N(_00884_),
    .Y(_00886_));
 sky130_fd_sc_hd__o21ai_1 _08702_ (.A1(_00885_),
    .A2(_00886_),
    .B1(net31),
    .Y(_00887_));
 sky130_fd_sc_hd__nand2_4 _08703_ (.A(_00861_),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_4 _08704_ (.A(_07256_),
    .B(_07259_),
    .Y(_00889_));
 sky130_fd_sc_hd__nor3b_2 _08705_ (.A(_00889_),
    .B(_07206_),
    .C_N(_07821_),
    .Y(_00890_));
 sky130_fd_sc_hd__o211ai_2 _08706_ (.A1(_00842_),
    .A2(_00843_),
    .B1(_00890_),
    .C1(_00810_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2_4 _08707_ (.A(_07821_),
    .B(_00889_),
    .Y(_00892_));
 sky130_fd_sc_hd__o2111ai_1 _08708_ (.A1(_00797_),
    .A2(_00779_),
    .B1(_00810_),
    .C1(_00824_),
    .D1(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__xnor2_1 _08709_ (.A(_07821_),
    .B(_00841_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3_1 _08710_ (.A(_07256_),
    .B(_07259_),
    .C(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_07206_),
    .B(_00892_),
    .Y(_00896_));
 sky130_fd_sc_hd__mux2_4 _08712_ (.A0(_00895_),
    .A1(_00896_),
    .S(_00810_),
    .X(_00897_));
 sky130_fd_sc_hd__nand3_4 _08713_ (.A(_00891_),
    .B(_00893_),
    .C(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand4_4 _08714_ (.A(_00756_),
    .B(_00796_),
    .C(_00898_),
    .D(_00817_),
    .Y(_00899_));
 sky130_fd_sc_hd__xor2_1 _08715_ (.A(_07821_),
    .B(_00838_),
    .X(_00900_));
 sky130_fd_sc_hd__or3_1 _08716_ (.A(_00847_),
    .B(_00889_),
    .C(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__a21o_1 _08717_ (.A1(_07270_),
    .A2(_07261_),
    .B1(_07269_),
    .X(_00902_));
 sky130_fd_sc_hd__a21o_1 _08718_ (.A1(_07259_),
    .A2(_00902_),
    .B1(_07258_),
    .X(_00903_));
 sky130_fd_sc_hd__a21oi_2 _08719_ (.A1(_07256_),
    .A2(_00903_),
    .B1(_07255_),
    .Y(_00904_));
 sky130_fd_sc_hd__o221ai_4 _08720_ (.A1(_00899_),
    .A2(_00847_),
    .B1(_00901_),
    .B2(_00819_),
    .C1(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__or2_4 _08721_ (.A(_00905_),
    .B(_07252_),
    .X(_00906_));
 sky130_fd_sc_hd__a22oi_4 clone10 (.A1(_01172_),
    .A2(_01231_),
    .B1(_01245_),
    .B2(_01237_),
    .Y(net10));
 sky130_fd_sc_hd__and2_1 _08723_ (.A(_00866_),
    .B(_00884_),
    .X(_07231_));
 sky130_fd_sc_hd__mux2i_4 _08724_ (.A0(_00858_),
    .A1(_07231_),
    .S(_00819_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand2_1 _08725_ (.A(_00855_),
    .B(_07262_),
    .Y(_00909_));
 sky130_fd_sc_hd__nor2_1 _08726_ (.A(_00812_),
    .B(_00909_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_2 _08727_ (.A(_07265_),
    .B(_07267_),
    .C(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__nor2_1 _08728_ (.A(_00882_),
    .B(_00880_),
    .Y(_00912_));
 sky130_fd_sc_hd__nor2_1 _08729_ (.A(_00597_),
    .B(_00883_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand3_1 _08730_ (.A(_00596_),
    .B(net9),
    .C(_00869_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _08731_ (.A(_00597_),
    .B(_00864_),
    .Y(_00915_));
 sky130_fd_sc_hd__or3_1 _08732_ (.A(_00596_),
    .B(_00810_),
    .C(_00864_),
    .X(_00916_));
 sky130_fd_sc_hd__o221ai_1 _08733_ (.A1(_00844_),
    .A2(_00914_),
    .B1(_00915_),
    .B2(net9),
    .C1(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_1 _08734_ (.A(_00596_),
    .B(_00869_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_1 _08735_ (.A(net9),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__nor3_1 _08736_ (.A(_00882_),
    .B(_00880_),
    .C(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__a311oi_2 _08737_ (.A1(_00844_),
    .A2(_00912_),
    .A3(_00913_),
    .B1(_00917_),
    .C1(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__or3_4 _08738_ (.A(_00911_),
    .B(_00899_),
    .C(_00921_),
    .X(_00922_));
 sky130_fd_sc_hd__nor2_1 _08739_ (.A(_00889_),
    .B(_00900_),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_1 _08740_ (.A(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__xnor2_1 _08741_ (.A(_00566_),
    .B(_00858_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(_00597_),
    .B(_00762_),
    .Y(_00926_));
 sky130_fd_sc_hd__nor2_1 _08743_ (.A(_00566_),
    .B(_00762_),
    .Y(_00927_));
 sky130_fd_sc_hd__a2bb2oi_1 _08744_ (.A1_N(_00795_),
    .A2_N(_00926_),
    .B1(_00756_),
    .B2(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_00748_),
    .B(_00762_),
    .Y(_00929_));
 sky130_fd_sc_hd__a21bo_1 _08746_ (.A1(_00795_),
    .A2(_00929_),
    .B1_N(_00756_),
    .X(_00930_));
 sky130_fd_sc_hd__nor2_2 _08747_ (.A(_00746_),
    .B(_00597_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand4b_1 _08748_ (.A_N(_00756_),
    .B(_00762_),
    .C(_00931_),
    .D(_00795_),
    .Y(_00932_));
 sky130_fd_sc_hd__a31oi_1 _08749_ (.A1(_00928_),
    .A2(_00930_),
    .A3(_00932_),
    .B1(_00805_),
    .Y(_00933_));
 sky130_fd_sc_hd__o41a_1 _08750_ (.A1(_00819_),
    .A2(_00924_),
    .A3(_00911_),
    .A4(_00925_),
    .B1(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__o211ai_4 _08751_ (.A1(_00593_),
    .A2(_00908_),
    .B1(_00922_),
    .C1(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__a21o_1 _08752_ (.A1(_00888_),
    .A2(_00906_),
    .B1(_00935_),
    .X(_00936_));
 sky130_fd_sc_hd__buf_6 _08753_ (.A(_00936_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_2 _08754_ (.A0(_07254_),
    .A1(_00854_),
    .S(_00937_),
    .X(_07271_));
 sky130_fd_sc_hd__o21a_1 _08755_ (.A1(_07290_),
    .A2(_07289_),
    .B1(_07288_),
    .X(_00938_));
 sky130_fd_sc_hd__o21a_1 _08756_ (.A1(_07287_),
    .A2(_00938_),
    .B1(_07285_),
    .X(_00939_));
 sky130_fd_sc_hd__o21a_1 _08757_ (.A1(_07284_),
    .A2(_00939_),
    .B1(_07282_),
    .X(_00940_));
 sky130_fd_sc_hd__o21a_1 _08758_ (.A1(_07281_),
    .A2(_00940_),
    .B1(_07279_),
    .X(_00941_));
 sky130_fd_sc_hd__o21a_1 _08759_ (.A1(_07278_),
    .A2(_00941_),
    .B1(_07276_),
    .X(_00942_));
 sky130_fd_sc_hd__nor2_4 _08760_ (.A(_00942_),
    .B(_07275_),
    .Y(_00943_));
 sky130_fd_sc_hd__xnor2_2 _08761_ (.A(_07273_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__and2_2 _08762_ (.A(_00922_),
    .B(_00934_),
    .X(_00945_));
 sky130_fd_sc_hd__a21boi_2 _08763_ (.A1(_00888_),
    .A2(_00906_),
    .B1_N(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__nor2b_1 _08764_ (.A(_07261_),
    .B_N(_00847_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_00923_),
    .B(_00848_),
    .Y(_00948_));
 sky130_fd_sc_hd__a21oi_2 _08766_ (.A1(_07256_),
    .A2(_00836_),
    .B1(_07255_),
    .Y(_00949_));
 sky130_fd_sc_hd__o221a_1 _08767_ (.A1(_00899_),
    .A2(_00947_),
    .B1(_00948_),
    .B2(net31),
    .C1(_00949_),
    .X(_00950_));
 sky130_fd_sc_hd__nand2b_1 _08768_ (.A_N(_07252_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__xnor2_1 _08769_ (.A(_00597_),
    .B(_00762_),
    .Y(_00952_));
 sky130_fd_sc_hd__a31oi_4 _08770_ (.A1(_00756_),
    .A2(_00796_),
    .A3(_00817_),
    .B1(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hd__xor2_4 _08771_ (.A(_00795_),
    .B(_00953_),
    .X(_00954_));
 sky130_fd_sc_hd__o21bai_2 _08772_ (.A1(_00593_),
    .A2(_00908_),
    .B1_N(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__a21o_1 _08773_ (.A1(_00888_),
    .A2(_00951_),
    .B1(_00955_),
    .X(_00956_));
 sky130_fd_sc_hd__and2_1 _08774_ (.A(_00756_),
    .B(_00796_),
    .X(_00957_));
 sky130_fd_sc_hd__xnor2_1 _08775_ (.A(_00598_),
    .B(_00790_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _08776_ (.A(_00815_),
    .B(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__o21ai_0 _08777_ (.A1(net9),
    .A2(_00959_),
    .B1(_00817_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_00957_),
    .B(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__o21ai_0 _08779_ (.A1(_00946_),
    .A2(_00956_),
    .B1(net30),
    .Y(_00962_));
 sky130_fd_sc_hd__o31a_2 _08780_ (.A1(_00946_),
    .A2(_00956_),
    .A3(_00961_),
    .B1(_00962_),
    .X(_00963_));
 sky130_fd_sc_hd__or2_2 _08781_ (.A(_00756_),
    .B(_00796_),
    .X(_00964_));
 sky130_fd_sc_hd__nor3b_1 _08782_ (.A(_00957_),
    .B(_00805_),
    .C_N(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__nor2_1 _08783_ (.A(_00805_),
    .B(_00964_),
    .Y(_00966_));
 sky130_fd_sc_hd__nor2_1 _08784_ (.A(_00946_),
    .B(_00956_),
    .Y(_00967_));
 sky130_fd_sc_hd__mux2i_4 _08785_ (.A0(_00965_),
    .A1(_00966_),
    .S(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__o221ai_4 _08786_ (.A1(_00899_),
    .A2(_00947_),
    .B1(_00948_),
    .B2(net31),
    .C1(_00949_),
    .Y(_00969_));
 sky130_fd_sc_hd__a211o_1 _08787_ (.A1(_00855_),
    .A2(_00969_),
    .B1(_00598_),
    .C1(_07252_),
    .X(_00970_));
 sky130_fd_sc_hd__nand3_1 _08788_ (.A(_00855_),
    .B(_00598_),
    .C(_00969_),
    .Y(_00971_));
 sky130_fd_sc_hd__a22oi_2 _08789_ (.A1(_00593_),
    .A2(_00945_),
    .B1(_00970_),
    .B2(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__a31oi_1 _08790_ (.A1(_00855_),
    .A2(_00905_),
    .A3(_00969_),
    .B1(_07252_),
    .Y(_00973_));
 sky130_fd_sc_hd__nor2_1 _08791_ (.A(_00566_),
    .B(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(_00855_),
    .B(_00598_),
    .Y(_00975_));
 sky130_fd_sc_hd__a211oi_1 _08793_ (.A1(_00922_),
    .A2(_00934_),
    .B1(_00950_),
    .C1(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__nor2b_1 _08794_ (.A(_07252_),
    .B_N(_00855_),
    .Y(_00977_));
 sky130_fd_sc_hd__and4_1 _08795_ (.A(_00566_),
    .B(_00905_),
    .C(_00950_),
    .D(_00977_),
    .X(_00978_));
 sky130_fd_sc_hd__xor2_1 _08796_ (.A(_07252_),
    .B(_00598_),
    .X(_00979_));
 sky130_fd_sc_hd__a221oi_1 _08797_ (.A1(_00922_),
    .A2(_00934_),
    .B1(_00969_),
    .B2(_00977_),
    .C1(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__o31ai_2 _08798_ (.A1(_00976_),
    .A2(_00978_),
    .A3(_00980_),
    .B1(_00908_),
    .Y(_00981_));
 sky130_fd_sc_hd__o31ai_4 _08799_ (.A1(_00908_),
    .A2(_00972_),
    .A3(_00974_),
    .B1(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__o2bb2ai_1 _08800_ (.A1_N(_00888_),
    .A2_N(_00906_),
    .B1(_00593_),
    .B2(_00908_),
    .Y(_00983_));
 sky130_fd_sc_hd__a211oi_4 _08801_ (.A1(_00888_),
    .A2(_00906_),
    .B1(_00945_),
    .C1(_00955_),
    .Y(_00984_));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(_00954_),
    .A2(_00983_),
    .B1(_00984_),
    .X(_00985_));
 sky130_fd_sc_hd__inv_2 _08803_ (.A(_00943_),
    .Y(_00986_));
 sky130_fd_sc_hd__a21oi_4 _08804_ (.A1(_00986_),
    .A2(_07273_),
    .B1(_07272_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _08805_ (.A(_00598_),
    .B(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2b_4 _08806_ (.A_N(_00987_),
    .B(_00597_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_4 _08807_ (.A(_00989_),
    .B(_00593_),
    .Y(_00990_));
 sky130_fd_sc_hd__xor2_2 _08808_ (.A(_00855_),
    .B(_00905_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2i_4 _08809_ (.A0(_00988_),
    .A1(_00990_),
    .S(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__nor3_1 _08810_ (.A(_07236_),
    .B(_07238_),
    .C(_00605_),
    .Y(_00993_));
 sky130_fd_sc_hd__nor3_1 _08811_ (.A(_00757_),
    .B(_00760_),
    .C(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__nor3_1 _08812_ (.A(_07198_),
    .B(_00780_),
    .C(_00781_),
    .Y(_00995_));
 sky130_fd_sc_hd__nor2b_4 _08813_ (.A(_07147_),
    .B_N(_00675_),
    .Y(_07148_));
 sky130_fd_sc_hd__nor3_1 _08814_ (.A(_07150_),
    .B(_07152_),
    .C(_07151_),
    .Y(_00996_));
 sky130_fd_sc_hd__o21ai_0 _08815_ (.A1(_00656_),
    .A2(_00996_),
    .B1(net36),
    .Y(_00997_));
 sky130_fd_sc_hd__o21a_1 _08816_ (.A1(_00660_),
    .A2(_07148_),
    .B1(_00997_),
    .X(_07179_));
 sky130_fd_sc_hd__nor2_1 _08817_ (.A(_07183_),
    .B(_00829_),
    .Y(_00998_));
 sky130_fd_sc_hd__xnor2_1 _08818_ (.A(_07181_),
    .B(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hd__mux2_2 _08819_ (.A0(_07179_),
    .A1(_00999_),
    .S(_00698_),
    .X(_07196_));
 sky130_fd_sc_hd__nand2_2 _08820_ (.A(_07196_),
    .B(_00844_),
    .Y(_01000_));
 sky130_fd_sc_hd__o31ai_4 _08821_ (.A1(_00867_),
    .A2(_00995_),
    .A3(_00844_),
    .B1(_01000_),
    .Y(_07217_));
 sky130_fd_sc_hd__xor2_1 _08822_ (.A(_07219_),
    .B(_00862_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_2 _08823_ (.A0(_07217_),
    .A1(_01001_),
    .S(_00883_),
    .X(_07234_));
 sky130_fd_sc_hd__mux2i_4 _08824_ (.A0(_00994_),
    .A1(_07234_),
    .S(net30),
    .Y(_01002_));
 sky130_fd_sc_hd__inv_2 _08825_ (.A(_01002_),
    .Y(_07251_));
 sky130_fd_sc_hd__mux2i_4 _08826_ (.A0(_00988_),
    .A1(_00990_),
    .S(_07251_),
    .Y(_01003_));
 sky130_fd_sc_hd__a21oi_4 _08827_ (.A1(_00888_),
    .A2(_00906_),
    .B1(_00935_),
    .Y(_01004_));
 sky130_fd_sc_hd__mux2i_4 _08828_ (.A0(_00992_),
    .A1(_01003_),
    .S(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__or3_4 _08829_ (.A(_00982_),
    .B(_01005_),
    .C(_00985_),
    .X(_01006_));
 sky130_fd_sc_hd__buf_6 _08830_ (.A(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__a21o_4 _08831_ (.A1(_00963_),
    .A2(_00968_),
    .B1(_01007_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_4 _08832_ (.A0(_07271_),
    .A1(_00944_),
    .S(_01008_),
    .X(_01009_));
 sky130_fd_sc_hd__o21a_1 _08833_ (.A1(_07304_),
    .A2(_07303_),
    .B1(_07296_),
    .X(_01010_));
 sky130_fd_sc_hd__o21a_1 _08834_ (.A1(_07295_),
    .A2(_01010_),
    .B1(_07293_),
    .X(_01011_));
 sky130_fd_sc_hd__o21a_1 _08835_ (.A1(_07292_),
    .A2(_01011_),
    .B1(_07302_),
    .X(_01012_));
 sky130_fd_sc_hd__o21a_1 _08836_ (.A1(_07301_),
    .A2(_01012_),
    .B1(_07299_),
    .X(_01013_));
 sky130_fd_sc_hd__o21ai_1 _08837_ (.A1(_01013_),
    .A2(_07298_),
    .B1(_07310_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2b_2 _08838_ (.A_N(_07309_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__a21oi_4 _08839_ (.A1(_01015_),
    .A2(_07307_),
    .B1(_07306_),
    .Y(_01016_));
 sky130_fd_sc_hd__xnor2_2 _08840_ (.A(_00855_),
    .B(_00905_),
    .Y(_01017_));
 sky130_fd_sc_hd__a211oi_2 _08841_ (.A1(_00888_),
    .A2(_00906_),
    .B1(_00935_),
    .C1(_07251_),
    .Y(_01018_));
 sky130_fd_sc_hd__a21oi_2 _08842_ (.A1(_00937_),
    .A2(_01017_),
    .B1(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__nor2_2 _08843_ (.A(_00982_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand4_1 _08844_ (.A(_07290_),
    .B(_07273_),
    .C(_07285_),
    .D(_07288_),
    .Y(_01021_));
 sky130_fd_sc_hd__nor2_1 _08845_ (.A(_00812_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand4_1 _08846_ (.A(_07276_),
    .B(_07279_),
    .C(_07282_),
    .D(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__a211oi_1 _08847_ (.A1(_00936_),
    .A2(_01017_),
    .B1(_01018_),
    .C1(_00598_),
    .Y(_01024_));
 sky130_fd_sc_hd__a211oi_2 _08848_ (.A1(_00888_),
    .A2(_00906_),
    .B1(_00935_),
    .C1(_01002_),
    .Y(_01025_));
 sky130_fd_sc_hd__a211oi_1 _08849_ (.A1(_00936_),
    .A2(_00991_),
    .B1(_01025_),
    .C1(_00566_),
    .Y(_01026_));
 sky130_fd_sc_hd__a21oi_4 _08850_ (.A1(_00954_),
    .A2(_00983_),
    .B1(_00984_),
    .Y(_01027_));
 sky130_fd_sc_hd__o31ai_2 _08851_ (.A1(_01023_),
    .A2(_01024_),
    .A3(_01026_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__a21oi_4 _08852_ (.A1(_00963_),
    .A2(_00968_),
    .B1(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__xnor2_1 _08853_ (.A(_00566_),
    .B(_00987_),
    .Y(_01030_));
 sky130_fd_sc_hd__and2_0 _08854_ (.A(_01019_),
    .B(_01030_),
    .X(_01031_));
 sky130_fd_sc_hd__nor2_1 _08855_ (.A(_01019_),
    .B(_01030_),
    .Y(_01032_));
 sky130_fd_sc_hd__a221oi_4 _08856_ (.A1(_01020_),
    .A2(_01029_),
    .B1(_01031_),
    .B2(_01008_),
    .C1(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(_00961_),
    .B(_00964_),
    .Y(_01034_));
 sky130_fd_sc_hd__o21bai_1 _08858_ (.A1(_00946_),
    .A2(_00956_),
    .B1_N(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__or3b_1 _08859_ (.A(_00946_),
    .B(_00956_),
    .C_N(_01034_),
    .X(_01036_));
 sky130_fd_sc_hd__o21ai_2 _08860_ (.A1(_00957_),
    .A2(_00984_),
    .B1(_00964_),
    .Y(_01037_));
 sky130_fd_sc_hd__a22oi_2 _08861_ (.A1(_01035_),
    .A2(_01036_),
    .B1(_01037_),
    .B2(_00805_),
    .Y(_01038_));
 sky130_fd_sc_hd__o31a_1 _08862_ (.A1(_00908_),
    .A2(_00972_),
    .A3(_00974_),
    .B1(_00981_),
    .X(_01039_));
 sky130_fd_sc_hd__buf_2 _08863_ (.A(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__or2_0 _08864_ (.A(_00598_),
    .B(_00987_),
    .X(_01041_));
 sky130_fd_sc_hd__a211oi_1 _08865_ (.A1(_00937_),
    .A2(_00991_),
    .B1(_01041_),
    .C1(_01025_),
    .Y(_01042_));
 sky130_fd_sc_hd__and2_0 _08866_ (.A(_01040_),
    .B(_01042_),
    .X(_01043_));
 sky130_fd_sc_hd__a31oi_4 _08867_ (.A1(_01027_),
    .A2(_01020_),
    .A3(_01038_),
    .B1(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_00746_),
    .B(_01040_),
    .Y(_01045_));
 sky130_fd_sc_hd__and3_1 _08869_ (.A(_00566_),
    .B(_00987_),
    .C(_01019_),
    .X(_01046_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_00599_),
    .B(_00987_),
    .Y(_01047_));
 sky130_fd_sc_hd__a211oi_1 _08871_ (.A1(_00937_),
    .A2(_00991_),
    .B1(_01025_),
    .C1(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__a211oi_1 _08872_ (.A1(_00937_),
    .A2(_01017_),
    .B1(_00989_),
    .C1(_01018_),
    .Y(_01049_));
 sky130_fd_sc_hd__mux2i_1 _08873_ (.A0(_01048_),
    .A1(_01049_),
    .S(_01040_),
    .Y(_01050_));
 sky130_fd_sc_hd__a21boi_2 _08874_ (.A1(_01045_),
    .A2(_01046_),
    .B1_N(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__and2_1 _08875_ (.A(_01035_),
    .B(_01036_),
    .X(_01052_));
 sky130_fd_sc_hd__o211ai_1 _08876_ (.A1(_00982_),
    .A2(_01005_),
    .B1(_01035_),
    .C1(_01036_),
    .Y(_01053_));
 sky130_fd_sc_hd__a21oi_1 _08877_ (.A1(_00805_),
    .A2(_01037_),
    .B1(_00985_),
    .Y(_01054_));
 sky130_fd_sc_hd__a2bb2oi_1 _08878_ (.A1_N(_01007_),
    .A2_N(_01052_),
    .B1(_01053_),
    .B2(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__a21oi_2 _08879_ (.A1(_01044_),
    .A2(_01051_),
    .B1(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__buf_4 _08880_ (.A(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__a21oi_1 _08881_ (.A1(_01016_),
    .A2(_01033_),
    .B1(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__buf_6 _08882_ (.A(_01008_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2i_1 _08883_ (.A0(_07271_),
    .A1(_00944_),
    .S(net22),
    .Y(_01060_));
 sky130_fd_sc_hd__nand3_1 _08884_ (.A(_01016_),
    .B(_01060_),
    .C(_01057_),
    .Y(_01061_));
 sky130_fd_sc_hd__o31a_1 _08885_ (.A1(_00567_),
    .A2(_01009_),
    .A3(_01058_),
    .B1(_01061_),
    .X(_01062_));
 sky130_fd_sc_hd__and4_1 _08886_ (.A(_01016_),
    .B(_00931_),
    .C(_01009_),
    .D(_01033_),
    .X(_01063_));
 sky130_fd_sc_hd__nand2b_4 _08887_ (.A_N(_01016_),
    .B(_00598_),
    .Y(_01064_));
 sky130_fd_sc_hd__nor3_1 _08888_ (.A(_01064_),
    .B(_01060_),
    .C(_01033_),
    .Y(_01065_));
 sky130_fd_sc_hd__or2_2 _08889_ (.A(_00599_),
    .B(_01016_),
    .X(_01066_));
 sky130_fd_sc_hd__a21oi_4 clone5 (.A1(_01173_),
    .A2(_01187_),
    .B1(_01200_),
    .Y(net5));
 sky130_fd_sc_hd__nor2_2 _08891_ (.A(_00944_),
    .B(_01066_),
    .Y(_01068_));
 sky130_fd_sc_hd__and3_1 _08892_ (.A(_01016_),
    .B(_00748_),
    .C(_00944_),
    .X(_01069_));
 sky130_fd_sc_hd__o21ai_0 _08893_ (.A1(_01068_),
    .A2(_01069_),
    .B1(net22),
    .Y(_01070_));
 sky130_fd_sc_hd__nor2_2 _08894_ (.A(_07271_),
    .B(_01066_),
    .Y(_01071_));
 sky130_fd_sc_hd__and3_1 _08895_ (.A(_01016_),
    .B(_00748_),
    .C(_07271_),
    .X(_01072_));
 sky130_fd_sc_hd__a21oi_4 _08896_ (.A1(_00963_),
    .A2(_00968_),
    .B1(_01007_),
    .Y(_01073_));
 sky130_fd_sc_hd__o21ai_0 _08897_ (.A1(_01071_),
    .A2(_01072_),
    .B1(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21oi_1 _08898_ (.A1(_01070_),
    .A2(_01074_),
    .B1(_01033_),
    .Y(_01075_));
 sky130_fd_sc_hd__nor3_1 _08899_ (.A(_01063_),
    .B(_01065_),
    .C(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__o21a_1 _08900_ (.A1(_07330_),
    .A2(_07329_),
    .B1(_07328_),
    .X(_01077_));
 sky130_fd_sc_hd__o21a_1 _08901_ (.A1(_07327_),
    .A2(_01077_),
    .B1(_07325_),
    .X(_01078_));
 sky130_fd_sc_hd__o21a_1 _08902_ (.A1(_07324_),
    .A2(_01078_),
    .B1(_07322_),
    .X(_01079_));
 sky130_fd_sc_hd__o21a_1 _08903_ (.A1(_07321_),
    .A2(_01079_),
    .B1(_07319_),
    .X(_01080_));
 sky130_fd_sc_hd__o21a_1 _08904_ (.A1(_07318_),
    .A2(_01080_),
    .B1(_07316_),
    .X(_01081_));
 sky130_fd_sc_hd__nor2_4 _08905_ (.A(_01081_),
    .B(_07315_),
    .Y(_01082_));
 sky130_fd_sc_hd__inv_2 _08906_ (.A(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_4 _08907_ (.A1(_01083_),
    .A2(_07313_),
    .B1(_07312_),
    .Y(_01084_));
 sky130_fd_sc_hd__o21ai_2 _08908_ (.A1(_00566_),
    .A2(_01084_),
    .B1(_00593_),
    .Y(_01085_));
 sky130_fd_sc_hd__nor2_1 _08909_ (.A(_00599_),
    .B(_01084_),
    .Y(_01086_));
 sky130_fd_sc_hd__o21bai_1 _08910_ (.A1(_00847_),
    .A2(_00845_),
    .B1_N(_00902_),
    .Y(_01087_));
 sky130_fd_sc_hd__xnor2_1 _08911_ (.A(_07259_),
    .B(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__nor2_1 _08912_ (.A(_07242_),
    .B(_00603_),
    .Y(_01089_));
 sky130_fd_sc_hd__nor3_1 _08913_ (.A(_07206_),
    .B(_07204_),
    .C(_07205_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _08914_ (.A(_07186_),
    .B(_00710_),
    .Y(_07202_));
 sky130_fd_sc_hd__nand2_1 _08915_ (.A(_00844_),
    .B(_07202_),
    .Y(_01091_));
 sky130_fd_sc_hd__o31ai_2 _08916_ (.A1(_00826_),
    .A2(_00844_),
    .A3(_01090_),
    .B1(_01091_),
    .Y(_07223_));
 sky130_fd_sc_hd__nor2_1 _08917_ (.A(_07227_),
    .B(_00839_),
    .Y(_01092_));
 sky130_fd_sc_hd__xnor2_1 _08918_ (.A(_07225_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__mux2_1 _08919_ (.A0(_07223_),
    .A1(_01093_),
    .S(_00883_),
    .X(_07240_));
 sky130_fd_sc_hd__nand2_2 _08920_ (.A(_00820_),
    .B(_07240_),
    .Y(_01094_));
 sky130_fd_sc_hd__o31ai_4 _08921_ (.A1(_00604_),
    .A2(_01089_),
    .A3(_00820_),
    .B1(_01094_),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_00937_),
    .B(_07257_),
    .Y(_01095_));
 sky130_fd_sc_hd__a21oi_2 _08923_ (.A1(_00937_),
    .A2(_01088_),
    .B1(_01095_),
    .Y(_07274_));
 sky130_fd_sc_hd__nor3_1 _08924_ (.A(_07276_),
    .B(_07278_),
    .C(_00941_),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_1 _08925_ (.A(_00942_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__mux2i_4 _08926_ (.A0(_07274_),
    .A1(_01097_),
    .S(net22),
    .Y(_01098_));
 sky130_fd_sc_hd__mux2i_2 _08927_ (.A0(_01085_),
    .A1(_01086_),
    .S(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__xor2_4 _08928_ (.A(_07307_),
    .B(_01015_),
    .X(_01100_));
 sky130_fd_sc_hd__nor3_1 _08929_ (.A(_00599_),
    .B(_01100_),
    .C(_01084_),
    .Y(_01101_));
 sky130_fd_sc_hd__a21oi_2 _08930_ (.A1(_01085_),
    .A2(_01100_),
    .B1(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_2 _08931_ (.A(_01064_),
    .B(_00593_),
    .Y(_01103_));
 sky130_fd_sc_hd__and2_4 _08932_ (.A(_01103_),
    .B(_00944_),
    .X(_01104_));
 sky130_fd_sc_hd__o21ai_4 _08933_ (.A1(_01068_),
    .A2(_01104_),
    .B1(net22),
    .Y(_01105_));
 sky130_fd_sc_hd__and2_4 _08934_ (.A(_01103_),
    .B(_07271_),
    .X(_01106_));
 sky130_fd_sc_hd__o21ai_4 _08935_ (.A1(_01106_),
    .A2(_01071_),
    .B1(_01073_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand3_4 _08936_ (.A(_01107_),
    .B(_01105_),
    .C(_01056_),
    .Y(_01108_));
 sky130_fd_sc_hd__mux2i_4 _08937_ (.A0(_01099_),
    .A1(_01102_),
    .S(net4),
    .Y(_01109_));
 sky130_fd_sc_hd__a21o_4 _08938_ (.A1(_01062_),
    .A2(_01076_),
    .B1(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__o21a_1 _08939_ (.A1(_01068_),
    .A2(_01104_),
    .B1(net22),
    .X(_01111_));
 sky130_fd_sc_hd__o21a_1 _08940_ (.A1(_01071_),
    .A2(_01106_),
    .B1(_01073_),
    .X(_01112_));
 sky130_fd_sc_hd__nor2_4 _08941_ (.A(_01112_),
    .B(_01111_),
    .Y(_01113_));
 sky130_fd_sc_hd__buf_6 _08942_ (.A(_00812_),
    .X(_01114_));
 sky130_fd_sc_hd__nand4_1 _08943_ (.A(_07330_),
    .B(_07322_),
    .C(_07325_),
    .D(_07328_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand3_1 _08944_ (.A(_07313_),
    .B(_07316_),
    .C(_07319_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor3_2 _08945_ (.A(_01114_),
    .B(_01115_),
    .C(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__xnor2_1 _08946_ (.A(_00567_),
    .B(_01098_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand4_2 _08947_ (.A(_01113_),
    .B(_01057_),
    .C(_01117_),
    .D(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__xnor2_1 _08948_ (.A(_00599_),
    .B(_01100_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _08949_ (.A(_00805_),
    .B(_01037_),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _08950_ (.A(_01007_),
    .B(_01052_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_2 _08951_ (.A(_01121_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__mux2i_4 _08952_ (.A0(_01104_),
    .A1(_01106_),
    .S(_01073_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _08953_ (.A(_01027_),
    .B(_01053_),
    .Y(_01125_));
 sky130_fd_sc_hd__a21oi_1 _08954_ (.A1(_01044_),
    .A2(_01051_),
    .B1(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hd__o211ai_4 _08955_ (.A1(_01009_),
    .A2(_01066_),
    .B1(_01124_),
    .C1(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__a32oi_4 _08956_ (.A1(net4),
    .A2(_01117_),
    .A3(_01120_),
    .B1(_01123_),
    .B2(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__and3_1 _08957_ (.A(_00805_),
    .B(_01052_),
    .C(_01037_),
    .X(_01129_));
 sky130_fd_sc_hd__a21oi_1 _08958_ (.A1(_01027_),
    .A2(_01121_),
    .B1(_01052_),
    .Y(_01130_));
 sky130_fd_sc_hd__mux2i_1 _08959_ (.A0(_01129_),
    .A1(_01130_),
    .S(net32),
    .Y(_01131_));
 sky130_fd_sc_hd__nor3_1 _08960_ (.A(_01007_),
    .B(_01052_),
    .C(_01029_),
    .Y(_01132_));
 sky130_fd_sc_hd__a21oi_1 _08961_ (.A1(net32),
    .A2(_01052_),
    .B1(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand3_1 _08962_ (.A(_01027_),
    .B(_01020_),
    .C(_01038_),
    .Y(_01134_));
 sky130_fd_sc_hd__nand2_1 _08963_ (.A(_01040_),
    .B(_01042_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand4_1 _08964_ (.A(_00931_),
    .B(_00982_),
    .C(_00987_),
    .D(_01019_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand4_1 _08965_ (.A(_00748_),
    .B(_01040_),
    .C(_00987_),
    .D(_01019_),
    .Y(_01137_));
 sky130_fd_sc_hd__a41o_1 _08966_ (.A1(_01135_),
    .A2(_01050_),
    .A3(_01136_),
    .A4(_01137_),
    .B1(_00985_),
    .X(_01138_));
 sky130_fd_sc_hd__o21ai_1 _08967_ (.A1(_01005_),
    .A2(_01134_),
    .B1(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__o211ai_1 _08968_ (.A1(_01009_),
    .A2(_01066_),
    .B1(_01124_),
    .C1(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__mux2_4 _08969_ (.A0(_01131_),
    .A1(_01133_),
    .S(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__nand3_4 _08970_ (.A(_01119_),
    .B(_01128_),
    .C(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2b_1 _08971_ (.A_N(_01005_),
    .B(_01040_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand2_1 _08972_ (.A(_00985_),
    .B(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__o21a_1 _08973_ (.A1(net32),
    .A2(_01029_),
    .B1(_01144_),
    .X(_01145_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_00982_),
    .B(_01005_),
    .Y(_01146_));
 sky130_fd_sc_hd__o21ai_0 _08975_ (.A1(_01143_),
    .A2(_01029_),
    .B1(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__o31ai_1 _08976_ (.A1(_01111_),
    .A2(_01112_),
    .A3(_01033_),
    .B1(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__a21boi_0 _08977_ (.A1(_01044_),
    .A2(_01051_),
    .B1_N(_01055_),
    .Y(_01149_));
 sky130_fd_sc_hd__o211ai_1 _08978_ (.A1(_01009_),
    .A2(_01066_),
    .B1(_01124_),
    .C1(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hd__and2_1 _08979_ (.A(_01148_),
    .B(_01150_),
    .X(_01151_));
 sky130_fd_sc_hd__nand2_4 _08980_ (.A(_01145_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor3_1 _08981_ (.A(_07316_),
    .B(_07318_),
    .C(_01080_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _08982_ (.A(_01081_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__o31ai_1 _08983_ (.A1(_01110_),
    .A2(_01142_),
    .A3(_01152_),
    .B1(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__a21oi_2 _08984_ (.A1(_01062_),
    .A2(_01076_),
    .B1(_01109_),
    .Y(_01156_));
 sky130_fd_sc_hd__buf_4 _08985_ (.A(_01156_),
    .X(_01157_));
 sky130_fd_sc_hd__and3_2 _08986_ (.A(_01119_),
    .B(_01128_),
    .C(_01141_),
    .X(_01158_));
 sky130_fd_sc_hd__and3_1 _08987_ (.A(_01145_),
    .B(_01148_),
    .C(_01150_),
    .X(_01159_));
 sky130_fd_sc_hd__buf_2 _08988_ (.A(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__nor3_1 _08989_ (.A(_07282_),
    .B(_07284_),
    .C(_00939_),
    .Y(_01161_));
 sky130_fd_sc_hd__nor3_1 _08990_ (.A(_07248_),
    .B(_07250_),
    .C(_07249_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_4 _08991_ (.A(_07230_),
    .B(_00822_),
    .Y(_07246_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(net30),
    .B(_07246_),
    .Y(_01163_));
 sky130_fd_sc_hd__o31ai_2 _08993_ (.A1(_00601_),
    .A2(net30),
    .A3(_01162_),
    .B1(_01163_),
    .Y(_07260_));
 sky130_fd_sc_hd__nor2_1 _08994_ (.A(_00937_),
    .B(_07260_),
    .Y(_01164_));
 sky130_fd_sc_hd__or3_1 _08995_ (.A(_07262_),
    .B(_07264_),
    .C(_00846_),
    .X(_01165_));
 sky130_fd_sc_hd__a21oi_1 _08996_ (.A1(_00847_),
    .A2(_01165_),
    .B1(_01004_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _08997_ (.A(_01166_),
    .B(_01164_),
    .Y(_07280_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(_01073_),
    .B(_07280_),
    .Y(_01167_));
 sky130_fd_sc_hd__o31ai_2 _08999_ (.A1(_00940_),
    .A2(_01073_),
    .A3(_01161_),
    .B1(_01167_),
    .Y(_07297_));
 sky130_fd_sc_hd__nor3_1 _09000_ (.A(_07299_),
    .B(_07301_),
    .C(_01012_),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_1 _09001_ (.A(_01013_),
    .B(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__mux2_2 _09002_ (.A0(_07297_),
    .A1(_01169_),
    .S(net4),
    .X(_07314_));
 sky130_fd_sc_hd__nand4_2 _09003_ (.A(_01157_),
    .B(_01158_),
    .C(_01160_),
    .D(_07314_),
    .Y(_01170_));
 sky130_fd_sc_hd__and2_1 _09004_ (.A(_01155_),
    .B(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2i_4 _09005_ (.A0(_00595_),
    .A1(_00600_),
    .S(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand3_4 _09006_ (.A(_01156_),
    .B(_01158_),
    .C(_01160_),
    .Y(_01173_));
 sky130_fd_sc_hd__xor2_2 _09007_ (.A(_07313_),
    .B(_01082_),
    .X(_01174_));
 sky130_fd_sc_hd__xnor2_1 _09008_ (.A(_00599_),
    .B(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__o21a_4 _09009_ (.A1(_07350_),
    .A2(_07349_),
    .B1(_07348_),
    .X(_01176_));
 sky130_fd_sc_hd__o21a_1 _09010_ (.A1(_07347_),
    .A2(_01176_),
    .B1(_07345_),
    .X(_01177_));
 sky130_fd_sc_hd__o21a_1 _09011_ (.A1(_01177_),
    .A2(_07344_),
    .B1(_07342_),
    .X(_01178_));
 sky130_fd_sc_hd__o21a_1 _09012_ (.A1(_07341_),
    .A2(_01178_),
    .B1(_07339_),
    .X(_01179_));
 sky130_fd_sc_hd__o21a_1 _09013_ (.A1(_01179_),
    .A2(_07338_),
    .B1(_07336_),
    .X(_01180_));
 sky130_fd_sc_hd__o21a_1 _09014_ (.A1(_07335_),
    .A2(_01180_),
    .B1(_07333_),
    .X(_01181_));
 sky130_fd_sc_hd__nor2_4 _09015_ (.A(_01181_),
    .B(_07332_),
    .Y(_01182_));
 sky130_fd_sc_hd__o22ai_1 _09016_ (.A1(_00594_),
    .A2(_01174_),
    .B1(_01175_),
    .B2(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__inv_1 _09017_ (.A(_01098_),
    .Y(_07305_));
 sky130_fd_sc_hd__mux2i_4 _09018_ (.A0(_07305_),
    .A1(_01100_),
    .S(net4),
    .Y(_01184_));
 sky130_fd_sc_hd__xnor2_1 _09019_ (.A(_00567_),
    .B(_01084_),
    .Y(_01185_));
 sky130_fd_sc_hd__xnor2_1 _09020_ (.A(_01184_),
    .B(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_2 _09021_ (.A(_01183_),
    .B(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__xnor2_1 _09022_ (.A(_07270_),
    .B(_00848_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_1 _09023_ (.A(_00937_),
    .B(_07268_),
    .Y(_01189_));
 sky130_fd_sc_hd__a21oi_1 _09024_ (.A1(_00937_),
    .A2(_01188_),
    .B1(_01189_),
    .Y(_07277_));
 sky130_fd_sc_hd__nor3_1 _09025_ (.A(_07279_),
    .B(_07281_),
    .C(_00940_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _09026_ (.A(_00941_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__mux2_1 _09027_ (.A0(_07277_),
    .A1(_01191_),
    .S(_01059_),
    .X(_07308_));
 sky130_fd_sc_hd__o2111a_1 _09028_ (.A1(_01009_),
    .A2(_01066_),
    .B1(_01124_),
    .C1(_01057_),
    .D1(_07308_),
    .X(_01192_));
 sky130_fd_sc_hd__nor2_1 _09029_ (.A(_07298_),
    .B(_01013_),
    .Y(_01193_));
 sky130_fd_sc_hd__xor2_1 _09030_ (.A(_07310_),
    .B(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a31oi_2 _09031_ (.A1(_01105_),
    .A2(_01107_),
    .A3(_01057_),
    .B1(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__o21ai_1 _09032_ (.A1(_00567_),
    .A2(_01182_),
    .B1(_00593_),
    .Y(_01196_));
 sky130_fd_sc_hd__o21ai_1 _09033_ (.A1(_01192_),
    .A2(_01195_),
    .B1(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__or4_1 _09034_ (.A(_00599_),
    .B(_01182_),
    .C(_01192_),
    .D(_01195_),
    .X(_01198_));
 sky130_fd_sc_hd__nand3_1 _09035_ (.A(_01184_),
    .B(_01198_),
    .C(_01197_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor4_4 _09036_ (.A(_01152_),
    .B(_01142_),
    .C(_01110_),
    .D(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__a21oi_4 _09037_ (.A1(_01173_),
    .A2(_01187_),
    .B1(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__o21ai_2 _09038_ (.A1(net32),
    .A2(_01029_),
    .B1(_01144_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor3_1 _09039_ (.A(_01110_),
    .B(_01202_),
    .C(_01142_),
    .Y(_01203_));
 sky130_fd_sc_hd__or3_2 _09040_ (.A(_01111_),
    .B(_01112_),
    .C(_01057_),
    .X(_01204_));
 sky130_fd_sc_hd__xnor2_2 _09041_ (.A(_01033_),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_00567_),
    .B(_01016_),
    .Y(_01206_));
 sky130_fd_sc_hd__nor3_1 _09043_ (.A(_01064_),
    .B(_01009_),
    .C(_01057_),
    .Y(_01207_));
 sky130_fd_sc_hd__a31o_1 _09044_ (.A1(_01064_),
    .A2(_01009_),
    .A3(_01206_),
    .B1(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__nand3_1 _09045_ (.A(_00931_),
    .B(_01009_),
    .C(_01057_),
    .Y(_01209_));
 sky130_fd_sc_hd__o31ai_4 _09046_ (.A1(_01009_),
    .A2(_01057_),
    .A3(_01206_),
    .B1(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor3_4 _09047_ (.A(_01208_),
    .B(_01210_),
    .C(_01109_),
    .Y(_01211_));
 sky130_fd_sc_hd__o21ai_1 _09048_ (.A1(_01208_),
    .A2(_01210_),
    .B1(_01109_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor3b_1 _09049_ (.A(_01205_),
    .B(_01211_),
    .C_N(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__nor2_2 _09050_ (.A(_01203_),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor3_4 _09051_ (.A(_01152_),
    .B(_01142_),
    .C(_01110_),
    .Y(_01215_));
 sky130_fd_sc_hd__xnor2_1 _09052_ (.A(_01040_),
    .B(_01005_),
    .Y(_01216_));
 sky130_fd_sc_hd__nand2_1 _09053_ (.A(_00985_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__a21oi_1 _09054_ (.A1(_01105_),
    .A2(_01107_),
    .B1(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__and3_1 _09055_ (.A(_01044_),
    .B(_01051_),
    .C(_01202_),
    .X(_01219_));
 sky130_fd_sc_hd__a311o_2 _09056_ (.A1(_01113_),
    .A2(_01055_),
    .A3(_01139_),
    .B1(_01218_),
    .C1(_01219_),
    .X(_01220_));
 sky130_fd_sc_hd__nand2b_1 _09057_ (.A_N(_01220_),
    .B(_01141_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _09058_ (.A(_01127_),
    .B(_01123_),
    .Y(_01222_));
 sky130_fd_sc_hd__buf_2 _09059_ (.A(_01151_),
    .X(_01223_));
 sky130_fd_sc_hd__nand2_1 _09060_ (.A(_01222_),
    .B(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor3_1 _09061_ (.A(_01157_),
    .B(_01221_),
    .C(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__nor2_1 _09062_ (.A(_01215_),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _09063_ (.A(_01192_),
    .B(_01195_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor4_2 _09064_ (.A(_01110_),
    .B(_01142_),
    .C(_01152_),
    .D(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__a31oi_2 _09065_ (.A1(_01157_),
    .A2(_01158_),
    .A3(_01160_),
    .B1(_01174_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_2 _09066_ (.A(_01228_),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor4b_4 _09067_ (.A(_01201_),
    .B(_01214_),
    .C(_01226_),
    .D_N(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__a21o_2 _09068_ (.A1(_01173_),
    .A2(_01187_),
    .B1(_01200_),
    .X(_01232_));
 sky130_fd_sc_hd__nor2_1 _09069_ (.A(_01157_),
    .B(_01221_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor4b_1 _09070_ (.A(_01205_),
    .B(_01224_),
    .C(_01211_),
    .D_N(_01212_),
    .Y(_01234_));
 sky130_fd_sc_hd__buf_6 _09071_ (.A(_01215_),
    .X(_01235_));
 sky130_fd_sc_hd__a21o_4 _09072_ (.A1(_01233_),
    .A2(_01234_),
    .B1(net15),
    .X(_01236_));
 sky130_fd_sc_hd__nand2_8 _09073_ (.A(_01232_),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__xnor2_2 _09074_ (.A(_00599_),
    .B(_01182_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor3_1 _09075_ (.A(_01228_),
    .B(_01229_),
    .C(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor3_1 _09076_ (.A(_07333_),
    .B(_07335_),
    .C(_01180_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_2 _09077_ (.A(_01181_),
    .B(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__mux2i_2 _09078_ (.A0(_00600_),
    .A1(_00595_),
    .S(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__inv_2 _09079_ (.A(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o21ai_0 _09080_ (.A1(_01228_),
    .A2(_01229_),
    .B1(_01238_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor3b_4 _09081_ (.A(_01243_),
    .B(_01239_),
    .C_N(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__a22o_1 _09082_ (.A1(_01172_),
    .A2(_01231_),
    .B1(_01237_),
    .B2(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__buf_4 _09083_ (.A(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__buf_6 _09084_ (.A(_00599_),
    .X(_01248_));
 sky130_fd_sc_hd__nand4_1 _09085_ (.A(_07368_),
    .B(_07359_),
    .C(_07362_),
    .D(_07365_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand3_1 _09086_ (.A(_07370_),
    .B(_07353_),
    .C(_07356_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor3_1 _09087_ (.A(_01114_),
    .B(_01249_),
    .C(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__and3_1 _09088_ (.A(_01248_),
    .B(_01241_),
    .C(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__nand3_1 _09089_ (.A(_01157_),
    .B(_01141_),
    .C(_01160_),
    .Y(_01253_));
 sky130_fd_sc_hd__a211oi_1 _09090_ (.A1(_01173_),
    .A2(_01187_),
    .B1(_01200_),
    .C1(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(_01183_),
    .B(_01186_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21o_1 _09092_ (.A1(_01197_),
    .A2(_01198_),
    .B1(_01184_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_2 _09093_ (.A0(_01255_),
    .A1(_01256_),
    .S(_01215_),
    .X(_01257_));
 sky130_fd_sc_hd__or2_0 _09094_ (.A(_01208_),
    .B(_01210_),
    .X(_01258_));
 sky130_fd_sc_hd__o41ai_1 _09095_ (.A1(_01205_),
    .A2(_01258_),
    .A3(_01142_),
    .A4(_01152_),
    .B1(_01211_),
    .Y(_01259_));
 sky130_fd_sc_hd__and2_2 _09096_ (.A(_01212_),
    .B(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__o211ai_4 _09097_ (.A1(_01222_),
    .A2(_01254_),
    .B1(_01257_),
    .C1(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__xor2_2 _09098_ (.A(_01033_),
    .B(_01204_),
    .X(_01262_));
 sky130_fd_sc_hd__o22ai_2 _09099_ (.A1(_01262_),
    .A2(_01211_),
    .B1(_01225_),
    .B2(net15),
    .Y(_01263_));
 sky130_fd_sc_hd__o221ai_1 _09100_ (.A1(_01203_),
    .A2(_01233_),
    .B1(_01211_),
    .B2(_01262_),
    .C1(_01223_),
    .Y(_01264_));
 sky130_fd_sc_hd__a31o_1 _09101_ (.A1(_01232_),
    .A2(_01263_),
    .A3(_01260_),
    .B1(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__a211o_4 _09102_ (.A1(_01237_),
    .A2(_01252_),
    .B1(_01261_),
    .C1(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__xnor2_1 _09103_ (.A(_01230_),
    .B(_01238_),
    .Y(_01267_));
 sky130_fd_sc_hd__a21oi_1 _09104_ (.A1(_01233_),
    .A2(_01234_),
    .B1(net15),
    .Y(_01268_));
 sky130_fd_sc_hd__clkbuf_4 _09105_ (.A(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__o21ai_2 _09106_ (.A1(_01201_),
    .A2(_01269_),
    .B1(_01243_),
    .Y(_01270_));
 sky130_fd_sc_hd__o32ai_4 _09107_ (.A1(_01172_),
    .A2(_01230_),
    .A3(_01237_),
    .B1(_01267_),
    .B2(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__a21oi_4 _09108_ (.A1(_01247_),
    .A2(_01266_),
    .B1(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__a211oi_1 _09109_ (.A1(_01237_),
    .A2(_01252_),
    .B1(_01261_),
    .C1(_01265_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor3_1 _09110_ (.A(_07336_),
    .B(_07338_),
    .C(_01179_),
    .Y(_01274_));
 sky130_fd_sc_hd__o22ai_2 _09111_ (.A1(_01201_),
    .A2(_01269_),
    .B1(_01274_),
    .B2(_01180_),
    .Y(_01275_));
 sky130_fd_sc_hd__nor3_1 _09112_ (.A(_07302_),
    .B(_07292_),
    .C(_01011_),
    .Y(_01276_));
 sky130_fd_sc_hd__or2_0 _09113_ (.A(_01012_),
    .B(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__nor3_1 _09114_ (.A(_07265_),
    .B(_07267_),
    .C(_07266_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _09115_ (.A(_07250_),
    .B(_00820_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand2_2 _09116_ (.A(_01004_),
    .B(_07263_),
    .Y(_01279_));
 sky130_fd_sc_hd__o31ai_4 _09117_ (.A1(_00846_),
    .A2(_01278_),
    .A3(_01004_),
    .B1(_01279_),
    .Y(_07283_));
 sky130_fd_sc_hd__nor3_1 _09118_ (.A(_07285_),
    .B(_07287_),
    .C(_00938_),
    .Y(_01280_));
 sky130_fd_sc_hd__o21ai_0 _09119_ (.A1(_00939_),
    .A2(_01280_),
    .B1(_01059_),
    .Y(_01281_));
 sky130_fd_sc_hd__o21a_1 _09120_ (.A1(_01059_),
    .A2(_07283_),
    .B1(_01281_),
    .X(_07300_));
 sky130_fd_sc_hd__nor2_1 _09121_ (.A(_01108_),
    .B(_07300_),
    .Y(_01282_));
 sky130_fd_sc_hd__a21oi_2 _09122_ (.A1(_01108_),
    .A2(_01277_),
    .B1(_01282_),
    .Y(_07317_));
 sky130_fd_sc_hd__nor3_1 _09123_ (.A(_07319_),
    .B(_07321_),
    .C(_01079_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _09124_ (.A(_01080_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(_07317_),
    .A1(_01284_),
    .S(_01173_),
    .X(_07334_));
 sky130_fd_sc_hd__or3_1 _09126_ (.A(_01201_),
    .B(_01268_),
    .C(_07334_),
    .X(_01285_));
 sky130_fd_sc_hd__and2_0 _09127_ (.A(_01275_),
    .B(_01285_),
    .X(_07351_));
 sky130_fd_sc_hd__and3_1 _09128_ (.A(_01247_),
    .B(_01273_),
    .C(_07351_),
    .X(_01286_));
 sky130_fd_sc_hd__buf_4 _09129_ (.A(_01273_),
    .X(_01287_));
 sky130_fd_sc_hd__xor2_4 _09130_ (.A(_07353_),
    .B(_00590_),
    .X(_01288_));
 sky130_fd_sc_hd__a21oi_2 _09131_ (.A1(_01247_),
    .A2(_01287_),
    .B1(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__nor2_2 _09132_ (.A(_01286_),
    .B(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(_01157_),
    .B(_01223_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor3_2 _09134_ (.A(_01205_),
    .B(_01202_),
    .C(_01142_),
    .Y(_01292_));
 sky130_fd_sc_hd__or2_1 _09135_ (.A(_01157_),
    .B(_01223_),
    .X(_01293_));
 sky130_fd_sc_hd__o21ai_4 _09136_ (.A1(_01291_),
    .A2(_01292_),
    .B1(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__buf_6 _09137_ (.A(_01201_),
    .X(_01295_));
 sky130_fd_sc_hd__o22a_1 _09138_ (.A1(_01262_),
    .A2(_01211_),
    .B1(_01225_),
    .B2(net15),
    .X(_01296_));
 sky130_fd_sc_hd__nand2_2 _09139_ (.A(_01212_),
    .B(_01259_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor3_1 _09140_ (.A(_01295_),
    .B(_01296_),
    .C(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _09141_ (.A(_01262_),
    .B(_01211_),
    .Y(_01299_));
 sky130_fd_sc_hd__a2111oi_2 _09142_ (.A1(_01158_),
    .A2(_01160_),
    .B1(_01205_),
    .C1(_01258_),
    .D1(_01109_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_2 _09143_ (.A(_01299_),
    .B(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__o21ai_0 _09144_ (.A1(_01247_),
    .A2(_01298_),
    .B1(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__clkbuf_4 _09145_ (.A(_01232_),
    .X(_01303_));
 sky130_fd_sc_hd__inv_1 _09146_ (.A(_01171_),
    .Y(_07331_));
 sky130_fd_sc_hd__nand3_1 _09147_ (.A(_01303_),
    .B(_07331_),
    .C(_01236_),
    .Y(_01304_));
 sky130_fd_sc_hd__o21ai_1 _09148_ (.A1(net5),
    .A2(_01269_),
    .B1(_01241_),
    .Y(_01305_));
 sky130_fd_sc_hd__xnor2_2 _09149_ (.A(_01248_),
    .B(_00592_),
    .Y(_01306_));
 sky130_fd_sc_hd__a21oi_2 _09150_ (.A1(_01304_),
    .A2(_01305_),
    .B1(_01306_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor3_1 _09151_ (.A(net5),
    .B(_01171_),
    .C(_01269_),
    .Y(_01308_));
 sky130_fd_sc_hd__a21boi_1 _09152_ (.A1(_01232_),
    .A2(_01236_),
    .B1_N(_01241_),
    .Y(_01309_));
 sky130_fd_sc_hd__xnor2_1 _09153_ (.A(_00567_),
    .B(_00592_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor3_1 _09154_ (.A(_01308_),
    .B(_01309_),
    .C(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__xor2_1 _09155_ (.A(_01242_),
    .B(_01238_),
    .X(_01312_));
 sky130_fd_sc_hd__o21ai_0 _09156_ (.A1(net21),
    .A2(_01269_),
    .B1(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__o211ai_1 _09157_ (.A1(_01172_),
    .A2(_01237_),
    .B1(_01313_),
    .C1(_01230_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_8 _09158_ (.A(_01269_),
    .B(_01295_),
    .Y(_01315_));
 sky130_fd_sc_hd__a21oi_1 _09159_ (.A1(_01303_),
    .A2(_01236_),
    .B1(_01312_),
    .Y(_01316_));
 sky130_fd_sc_hd__a211o_1 _09160_ (.A1(_01172_),
    .A2(_01315_),
    .B1(_01316_),
    .C1(_01230_),
    .X(_01317_));
 sky130_fd_sc_hd__o211ai_1 _09161_ (.A1(_01307_),
    .A2(_01311_),
    .B1(_01314_),
    .C1(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_1 _09162_ (.A(_01308_),
    .B(_01309_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand3_2 _09163_ (.A(_01247_),
    .B(_01287_),
    .C(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__and2_1 _09164_ (.A(_01127_),
    .B(_01123_),
    .X(_01321_));
 sky130_fd_sc_hd__o211a_1 _09165_ (.A1(_01321_),
    .A2(_01221_),
    .B1(_01213_),
    .C1(_01223_),
    .X(_01322_));
 sky130_fd_sc_hd__nand3_1 _09166_ (.A(_01157_),
    .B(_01223_),
    .C(_01142_),
    .Y(_01323_));
 sky130_fd_sc_hd__and2_0 _09167_ (.A(_01157_),
    .B(_01223_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2i_2 _09168_ (.A0(_01323_),
    .A1(_01324_),
    .S(_01220_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21oi_2 _09169_ (.A1(_01303_),
    .A2(_01322_),
    .B1(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__mux2i_4 _09170_ (.A0(_01255_),
    .A1(_01256_),
    .S(net15),
    .Y(_01327_));
 sky130_fd_sc_hd__a211oi_2 _09171_ (.A1(_01232_),
    .A2(_01269_),
    .B1(_01297_),
    .C1(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _09172_ (.A(_01326_),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__a221oi_1 _09173_ (.A1(_01294_),
    .A2(_01302_),
    .B1(_01318_),
    .B2(_01320_),
    .C1(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__a211oi_1 _09174_ (.A1(_01303_),
    .A2(_01236_),
    .B1(_01241_),
    .C1(_01248_),
    .Y(_01331_));
 sky130_fd_sc_hd__a21oi_1 _09175_ (.A1(_01155_),
    .A2(_01170_),
    .B1(_01248_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand3_1 _09176_ (.A(_01248_),
    .B(_01155_),
    .C(_01170_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor4b_1 _09177_ (.A(net5),
    .B(_01269_),
    .C(_01332_),
    .D_N(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__o21ai_2 _09178_ (.A1(_01331_),
    .A2(_01334_),
    .B1(_01251_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_2 _09179_ (.A(_01287_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__a21o_1 _09180_ (.A1(_01246_),
    .A2(_01328_),
    .B1(_01298_),
    .X(_01337_));
 sky130_fd_sc_hd__or2_2 _09181_ (.A(_01299_),
    .B(_01300_),
    .X(_01338_));
 sky130_fd_sc_hd__o31ai_2 _09182_ (.A1(_01295_),
    .A2(_01296_),
    .A3(_01297_),
    .B1(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__a21oi_2 _09183_ (.A1(_01247_),
    .A2(_01328_),
    .B1(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__a31oi_4 _09184_ (.A1(_01301_),
    .A2(_01336_),
    .A3(_01337_),
    .B1(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o211a_1 _09185_ (.A1(_00594_),
    .A2(_01290_),
    .B1(_01330_),
    .C1(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__or2_1 _09186_ (.A(_01286_),
    .B(_01289_),
    .X(_01343_));
 sky130_fd_sc_hd__o21a_1 _09187_ (.A1(_07372_),
    .A2(_07371_),
    .B1(_07390_),
    .X(_01344_));
 sky130_fd_sc_hd__o21a_1 _09188_ (.A1(_07389_),
    .A2(_01344_),
    .B1(_07387_),
    .X(_01345_));
 sky130_fd_sc_hd__o21a_1 _09189_ (.A1(_07386_),
    .A2(_01345_),
    .B1(_07384_),
    .X(_01346_));
 sky130_fd_sc_hd__o21a_1 _09190_ (.A1(_07383_),
    .A2(_01346_),
    .B1(_07381_),
    .X(_01347_));
 sky130_fd_sc_hd__o21a_1 _09191_ (.A1(_07380_),
    .A2(_01347_),
    .B1(_07378_),
    .X(_01348_));
 sky130_fd_sc_hd__o21a_1 _09192_ (.A1(_01348_),
    .A2(_07377_),
    .B1(_07375_),
    .X(_01349_));
 sky130_fd_sc_hd__nor2_4 _09193_ (.A(_01349_),
    .B(_07374_),
    .Y(_01350_));
 sky130_fd_sc_hd__o21ai_1 _09194_ (.A1(net21),
    .A2(_01236_),
    .B1(_01257_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _09195_ (.A(_01350_),
    .B(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand3_1 _09196_ (.A(_00568_),
    .B(_01272_),
    .C(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__o2111ai_1 _09197_ (.A1(_01286_),
    .A2(_01289_),
    .B1(_01352_),
    .C1(_01272_),
    .D1(_01248_),
    .Y(_01354_));
 sky130_fd_sc_hd__o21a_1 _09198_ (.A1(_01343_),
    .A2(_01353_),
    .B1(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__a22oi_4 _09199_ (.A1(_01172_),
    .A2(_01231_),
    .B1(_01245_),
    .B2(_01237_),
    .Y(_01356_));
 sky130_fd_sc_hd__o211ai_4 _09200_ (.A1(net21),
    .A2(_01236_),
    .B1(_01260_),
    .C1(_01257_),
    .Y(_01357_));
 sky130_fd_sc_hd__a311oi_2 _09201_ (.A1(_01303_),
    .A2(_01263_),
    .A3(_01260_),
    .B1(_01338_),
    .C1(_01294_),
    .Y(_01358_));
 sky130_fd_sc_hd__o221ai_1 _09202_ (.A1(_01299_),
    .A2(_01300_),
    .B1(_01292_),
    .B2(_01291_),
    .C1(_01293_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor4_1 _09203_ (.A(_01295_),
    .B(_01296_),
    .C(_01297_),
    .D(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(_01323_),
    .A1(_01324_),
    .S(_01220_),
    .X(_01361_));
 sky130_fd_sc_hd__nor2_1 _09205_ (.A(_01110_),
    .B(_01152_),
    .Y(_01362_));
 sky130_fd_sc_hd__nand2_1 _09206_ (.A(_01119_),
    .B(_01128_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand4_1 _09207_ (.A(_01363_),
    .B(_01157_),
    .C(_01141_),
    .D(_01160_),
    .Y(_01364_));
 sky130_fd_sc_hd__o21ai_4 _09208_ (.A1(_01141_),
    .A2(_01362_),
    .B1(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__a211oi_2 _09209_ (.A1(_01303_),
    .A2(_01322_),
    .B1(_01361_),
    .C1(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__and4_1 _09210_ (.A(_01303_),
    .B(_01322_),
    .C(_01361_),
    .D(_01365_),
    .X(_01367_));
 sky130_fd_sc_hd__o21ai_1 _09211_ (.A1(_01203_),
    .A2(_01233_),
    .B1(_01223_),
    .Y(_01368_));
 sky130_fd_sc_hd__o311ai_4 _09212_ (.A1(_01368_),
    .A2(net5),
    .A3(_01214_),
    .B1(_01253_),
    .C1(_01321_),
    .Y(_01369_));
 sky130_fd_sc_hd__o221ai_4 _09213_ (.A1(_01358_),
    .A2(_01360_),
    .B1(_01366_),
    .B2(_01367_),
    .C1(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__o211ai_1 _09214_ (.A1(_01321_),
    .A2(_01221_),
    .B1(_01213_),
    .C1(_01223_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor3_1 _09215_ (.A(_01295_),
    .B(_01371_),
    .C(_01361_),
    .Y(_01372_));
 sky130_fd_sc_hd__inv_1 _09216_ (.A(_01365_),
    .Y(_01373_));
 sky130_fd_sc_hd__o211ai_2 _09217_ (.A1(_01326_),
    .A2(_01372_),
    .B1(_01369_),
    .C1(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__o31ai_4 _09218_ (.A1(_01356_),
    .A2(_01357_),
    .A3(_01370_),
    .B1(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_8 _09219_ (.A(_01266_),
    .B(_01356_),
    .Y(_01376_));
 sky130_fd_sc_hd__a211o_1 _09220_ (.A1(_01275_),
    .A2(_01285_),
    .B1(_01350_),
    .C1(_01248_),
    .X(_01377_));
 sky130_fd_sc_hd__o21ai_0 _09221_ (.A1(_00567_),
    .A2(_01350_),
    .B1(_00594_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand3_2 _09222_ (.A(_01275_),
    .B(_01285_),
    .C(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__and3_1 _09223_ (.A(_01377_),
    .B(_01319_),
    .C(_01379_),
    .X(_01380_));
 sky130_fd_sc_hd__o21ai_2 _09224_ (.A1(_01308_),
    .A2(_01309_),
    .B1(_01310_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand3_1 _09225_ (.A(_01304_),
    .B(_01305_),
    .C(_01306_),
    .Y(_01382_));
 sky130_fd_sc_hd__xnor2_1 _09226_ (.A(_01248_),
    .B(_01288_),
    .Y(_01383_));
 sky130_fd_sc_hd__o22ai_4 _09227_ (.A1(_00594_),
    .A2(_01288_),
    .B1(_01383_),
    .B2(_01350_),
    .Y(_01384_));
 sky130_fd_sc_hd__a221o_1 _09228_ (.A1(_01172_),
    .A2(_01231_),
    .B1(_01237_),
    .B2(_01245_),
    .C1(_01384_),
    .X(_01385_));
 sky130_fd_sc_hd__o21a_1 _09229_ (.A1(_01291_),
    .A2(_01292_),
    .B1(_01293_),
    .X(_01386_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_01386_),
    .B(_01328_),
    .Y(_01387_));
 sky130_fd_sc_hd__a2111oi_4 _09231_ (.A1(_01381_),
    .A2(_01382_),
    .B1(_01387_),
    .C1(_01271_),
    .D1(_01385_),
    .Y(_01388_));
 sky130_fd_sc_hd__a21o_1 _09232_ (.A1(_01376_),
    .A2(_01380_),
    .B1(_01388_),
    .X(_01389_));
 sky130_fd_sc_hd__nand3_4 _09233_ (.A(_01375_),
    .B(_01341_),
    .C(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor3_1 _09234_ (.A(net21),
    .B(_01371_),
    .C(_01325_),
    .Y(_01391_));
 sky130_fd_sc_hd__xnor2_2 _09235_ (.A(_01365_),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand4_1 _09236_ (.A(_01303_),
    .B(_01263_),
    .C(_01260_),
    .D(_01301_),
    .Y(_01393_));
 sky130_fd_sc_hd__a2111oi_2 _09237_ (.A1(_01303_),
    .A2(_01269_),
    .B1(_01297_),
    .C1(_01327_),
    .D1(_01294_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand3_1 _09238_ (.A(_01339_),
    .B(_01393_),
    .C(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__a211oi_1 _09239_ (.A1(_01287_),
    .A2(_01335_),
    .B1(_01356_),
    .C1(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__o21ai_1 _09240_ (.A1(_01326_),
    .A2(_01372_),
    .B1(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__xor2_2 _09241_ (.A(_01392_),
    .B(_01397_),
    .X(_01398_));
 sky130_fd_sc_hd__a31oi_4 _09242_ (.A1(_01342_),
    .A2(_01355_),
    .A3(_01390_),
    .B1(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__and4_1 _09243_ (.A(_01398_),
    .B(_01342_),
    .C(_01355_),
    .D(_01390_),
    .X(_01400_));
 sky130_fd_sc_hd__buf_6 _09244_ (.A(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__nor2_4 _09245_ (.A(_01004_),
    .B(_07267_),
    .Y(_07286_));
 sky130_fd_sc_hd__nor3_1 _09246_ (.A(_07290_),
    .B(_07288_),
    .C(_07289_),
    .Y(_01402_));
 sky130_fd_sc_hd__o21ai_0 _09247_ (.A1(_00938_),
    .A2(_01402_),
    .B1(_01059_),
    .Y(_01403_));
 sky130_fd_sc_hd__o21a_1 _09248_ (.A1(_07286_),
    .A2(_01059_),
    .B1(_01403_),
    .X(_07291_));
 sky130_fd_sc_hd__nor3_1 _09249_ (.A(_07293_),
    .B(_07295_),
    .C(_01010_),
    .Y(_01404_));
 sky130_fd_sc_hd__o21ai_0 _09250_ (.A1(_01011_),
    .A2(_01404_),
    .B1(_01108_),
    .Y(_01405_));
 sky130_fd_sc_hd__o21a_1 _09251_ (.A1(_01108_),
    .A2(_07291_),
    .B1(_01405_),
    .X(_07320_));
 sky130_fd_sc_hd__nand2_1 _09252_ (.A(_01235_),
    .B(_07320_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor3_1 _09253_ (.A(_07322_),
    .B(_07324_),
    .C(_01078_),
    .Y(_01407_));
 sky130_fd_sc_hd__or3_1 _09254_ (.A(_01079_),
    .B(_01235_),
    .C(_01407_),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_01406_),
    .B(_01408_),
    .Y(_07337_));
 sky130_fd_sc_hd__nor3_1 _09256_ (.A(_07339_),
    .B(_07341_),
    .C(_01178_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _09257_ (.A(_01179_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__mux2_1 _09258_ (.A0(_07337_),
    .A1(_01410_),
    .S(_01237_),
    .X(_07354_));
 sky130_fd_sc_hd__nand3_1 _09259_ (.A(_01247_),
    .B(_01287_),
    .C(_07354_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor3_1 _09260_ (.A(_07356_),
    .B(_07358_),
    .C(_00588_),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _09261_ (.A(_00589_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__o21ai_1 _09262_ (.A1(_01356_),
    .A2(_01266_),
    .B1(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__a21oi_1 _09263_ (.A1(_01411_),
    .A2(_01414_),
    .B1(_00568_),
    .Y(_01415_));
 sky130_fd_sc_hd__and3_1 _09264_ (.A(_00568_),
    .B(_01411_),
    .C(_01414_),
    .X(_01416_));
 sky130_fd_sc_hd__nand4_1 _09265_ (.A(_07393_),
    .B(_07404_),
    .C(_07407_),
    .D(_07410_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand3_1 _09266_ (.A(_07395_),
    .B(_07398_),
    .C(_07401_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor3_1 _09267_ (.A(_01114_),
    .B(_01417_),
    .C(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__o21ai_1 _09268_ (.A1(_01415_),
    .A2(_01416_),
    .B1(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hd__buf_4 _09269_ (.A(_01248_),
    .X(_01421_));
 sky130_fd_sc_hd__nor3_1 _09270_ (.A(_07375_),
    .B(_07377_),
    .C(_01348_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_2 _09271_ (.A(_01349_),
    .B(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__xnor2_1 _09272_ (.A(_01421_),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _09273_ (.A(_01419_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__buf_8 _09274_ (.A(_01390_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_4 _09275_ (.A0(_01420_),
    .A1(_01425_),
    .S(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(_01339_),
    .B(_01393_),
    .Y(_01428_));
 sky130_fd_sc_hd__o31a_1 _09277_ (.A1(_01110_),
    .A2(_01223_),
    .A3(_01221_),
    .B1(_01368_),
    .X(_01429_));
 sky130_fd_sc_hd__nor4_1 _09278_ (.A(net10),
    .B(_01428_),
    .C(_01357_),
    .D(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__a21oi_1 _09279_ (.A1(_01336_),
    .A2(_01430_),
    .B1(_01369_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _09280_ (.A(_01326_),
    .B(_01372_),
    .Y(_01432_));
 sky130_fd_sc_hd__xnor2_1 _09281_ (.A(_01432_),
    .B(_01396_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand4_1 _09282_ (.A(_01392_),
    .B(_01341_),
    .C(_01389_),
    .D(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_4 _09283_ (.A(_01431_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__a2111oi_1 _09284_ (.A1(_01381_),
    .A2(_01382_),
    .B1(_01385_),
    .C1(_01271_),
    .D1(_01357_),
    .Y(_01436_));
 sky130_fd_sc_hd__a21oi_2 _09285_ (.A1(_01376_),
    .A2(_01380_),
    .B1(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__nor2_1 _09286_ (.A(_01338_),
    .B(_01294_),
    .Y(_01438_));
 sky130_fd_sc_hd__o31a_2 _09287_ (.A1(_01356_),
    .A2(_01357_),
    .A3(_01370_),
    .B1(_01374_),
    .X(_01439_));
 sky130_fd_sc_hd__nand2_1 _09288_ (.A(_01438_),
    .B(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__o21a_1 _09289_ (.A1(_01437_),
    .A2(_01440_),
    .B1(_01433_),
    .X(_01441_));
 sky130_fd_sc_hd__nor3_1 _09290_ (.A(_01437_),
    .B(_01440_),
    .C(_01433_),
    .Y(_01442_));
 sky130_fd_sc_hd__o32a_1 _09291_ (.A1(_01172_),
    .A2(_01230_),
    .A3(_01237_),
    .B1(_01267_),
    .B2(_01270_),
    .X(_01443_));
 sky130_fd_sc_hd__o21ai_1 _09292_ (.A1(net10),
    .A2(_01287_),
    .B1(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor3_1 _09293_ (.A(_01387_),
    .B(_01439_),
    .C(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__and2_0 _09294_ (.A(_01341_),
    .B(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__clkbuf_2 _09295_ (.A(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__a21oi_1 _09296_ (.A1(_01381_),
    .A2(_01382_),
    .B1(_01385_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21oi_1 _09297_ (.A1(_01376_),
    .A2(_01380_),
    .B1(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand4_2 _09298_ (.A(_01394_),
    .B(_01443_),
    .C(_01377_),
    .D(_01379_),
    .Y(_01450_));
 sky130_fd_sc_hd__o22a_1 _09299_ (.A1(_00594_),
    .A2(_01288_),
    .B1(_01383_),
    .B2(_01350_),
    .X(_01451_));
 sky130_fd_sc_hd__o21ai_2 _09300_ (.A1(_01307_),
    .A2(_01311_),
    .B1(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__o221ai_4 _09301_ (.A1(_01320_),
    .A2(_01450_),
    .B1(_01452_),
    .B2(_01376_),
    .C1(_01444_),
    .Y(_01453_));
 sky130_fd_sc_hd__a21oi_1 _09302_ (.A1(_01303_),
    .A2(_01269_),
    .B1(_01327_),
    .Y(_01454_));
 sky130_fd_sc_hd__o21ai_1 _09303_ (.A1(net10),
    .A2(_01287_),
    .B1(_01454_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand3_1 _09304_ (.A(_01247_),
    .B(_01266_),
    .C(_01351_),
    .Y(_01456_));
 sky130_fd_sc_hd__a21oi_1 _09305_ (.A1(net21),
    .A2(_01297_),
    .B1(_01298_),
    .Y(_01457_));
 sky130_fd_sc_hd__a21boi_1 _09306_ (.A1(_01455_),
    .A2(_01456_),
    .B1_N(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__a311oi_1 _09307_ (.A1(_01301_),
    .A2(_01336_),
    .A3(_01337_),
    .B1(_01340_),
    .C1(_01294_),
    .Y(_01459_));
 sky130_fd_sc_hd__o2111a_1 _09308_ (.A1(_01271_),
    .A2(_01449_),
    .B1(_01453_),
    .C1(_01458_),
    .D1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__o22a_2 _09309_ (.A1(_01441_),
    .A2(_01442_),
    .B1(_01447_),
    .B2(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__o2111ai_4 _09310_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01427_),
    .C1(_01435_),
    .D1(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand4_1 _09311_ (.A(_01247_),
    .B(_01287_),
    .C(_01377_),
    .D(_01379_),
    .Y(_01463_));
 sky130_fd_sc_hd__xnor2_1 _09312_ (.A(_01306_),
    .B(_01451_),
    .Y(_01464_));
 sky130_fd_sc_hd__o21ai_0 _09313_ (.A1(net10),
    .A2(_01266_),
    .B1(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _09314_ (.A(_01304_),
    .B(_01305_),
    .Y(_01466_));
 sky130_fd_sc_hd__a21oi_1 _09315_ (.A1(_01463_),
    .A2(_01465_),
    .B1(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__and3_1 _09316_ (.A(_01466_),
    .B(_01463_),
    .C(_01465_),
    .X(_01468_));
 sky130_fd_sc_hd__xnor2_1 _09317_ (.A(_01248_),
    .B(_01350_),
    .Y(_01469_));
 sky130_fd_sc_hd__nor3_1 _09318_ (.A(_01286_),
    .B(_01289_),
    .C(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__o21ai_0 _09319_ (.A1(_01286_),
    .A2(_01289_),
    .B1(_01469_),
    .Y(_01471_));
 sky130_fd_sc_hd__nor4b_4 _09320_ (.A(_01467_),
    .B(_01468_),
    .C(_01470_),
    .D_N(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__a31o_2 _09321_ (.A1(_01301_),
    .A2(_01336_),
    .A3(_01337_),
    .B1(_01340_),
    .X(_01473_));
 sky130_fd_sc_hd__a21oi_4 _09322_ (.A1(_01376_),
    .A2(_01380_),
    .B1(_01388_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor4_2 _09323_ (.A(_01439_),
    .B(_01473_),
    .C(_01474_),
    .D(_01343_),
    .Y(_01475_));
 sky130_fd_sc_hd__o21a_1 _09324_ (.A1(_07395_),
    .A2(_07394_),
    .B1(_07393_),
    .X(_01476_));
 sky130_fd_sc_hd__o21a_1 _09325_ (.A1(_07392_),
    .A2(_01476_),
    .B1(_07410_),
    .X(_01477_));
 sky130_fd_sc_hd__o21a_1 _09326_ (.A1(_07409_),
    .A2(_01477_),
    .B1(_07407_),
    .X(_01478_));
 sky130_fd_sc_hd__o21a_1 _09327_ (.A1(_07406_),
    .A2(_01478_),
    .B1(_07404_),
    .X(_01479_));
 sky130_fd_sc_hd__o21a_1 _09328_ (.A1(_07403_),
    .A2(_01479_),
    .B1(_07401_),
    .X(_01480_));
 sky130_fd_sc_hd__nor2_4 _09329_ (.A(_01480_),
    .B(_07400_),
    .Y(_01481_));
 sky130_fd_sc_hd__inv_2 _09330_ (.A(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__a21oi_4 _09331_ (.A1(_01482_),
    .A2(_07398_),
    .B1(_07397_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _09332_ (.A(_01421_),
    .B(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__o21ai_4 _09333_ (.A1(_00567_),
    .A2(_01483_),
    .B1(_00594_),
    .Y(_01485_));
 sky130_fd_sc_hd__nand2_2 _09334_ (.A(_01411_),
    .B(_01414_),
    .Y(_07373_));
 sky130_fd_sc_hd__mux2i_4 _09335_ (.A0(_01484_),
    .A1(_01485_),
    .S(_07373_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor3_1 _09336_ (.A(_01421_),
    .B(_01423_),
    .C(_01483_),
    .Y(_01487_));
 sky130_fd_sc_hd__and2_4 _09337_ (.A(_01423_),
    .B(_01485_),
    .X(_01488_));
 sky130_fd_sc_hd__o32ai_4 _09338_ (.A1(_01439_),
    .A2(_01473_),
    .A3(_01474_),
    .B1(_01487_),
    .B2(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__o221a_4 _09339_ (.A1(_01472_),
    .A2(_01475_),
    .B1(_01486_),
    .B2(_01390_),
    .C1(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__o221a_1 clone27 (.A1(_01472_),
    .A2(_01475_),
    .B1(_01486_),
    .B2(_01390_),
    .C1(_01489_),
    .X(net27));
 sky130_fd_sc_hd__buf_6 _09341_ (.A(_01376_),
    .X(_01492_));
 sky130_fd_sc_hd__o22a_1 _09342_ (.A1(_01320_),
    .A2(_01450_),
    .B1(_01452_),
    .B2(net17),
    .X(_01493_));
 sky130_fd_sc_hd__nor2_2 _09343_ (.A(_01493_),
    .B(_01447_),
    .Y(_01494_));
 sky130_fd_sc_hd__o2bb2ai_1 _09344_ (.A1_N(_01272_),
    .A2_N(_01494_),
    .B1(_01490_),
    .B2(_01453_),
    .Y(_01495_));
 sky130_fd_sc_hd__a31oi_4 _09345_ (.A1(_01272_),
    .A2(_01462_),
    .A3(_01490_),
    .B1(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__o2111ai_4 _09346_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01461_),
    .C1(_01435_),
    .D1(_01490_),
    .Y(_01497_));
 sky130_fd_sc_hd__a31oi_2 _09347_ (.A1(_01375_),
    .A2(_01341_),
    .A3(_01389_),
    .B1(_01469_),
    .Y(_01498_));
 sky130_fd_sc_hd__xnor2_2 _09348_ (.A(_01290_),
    .B(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__xor2_2 _09349_ (.A(_01485_),
    .B(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__xnor2_2 _09350_ (.A(_00568_),
    .B(_01483_),
    .Y(_01501_));
 sky130_fd_sc_hd__mux2i_4 _09351_ (.A0(_07373_),
    .A1(_01423_),
    .S(_01426_),
    .Y(_01502_));
 sky130_fd_sc_hd__a31o_1 _09352_ (.A1(_01497_),
    .A2(_01500_),
    .A3(_01501_),
    .B1(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__and2_0 _09353_ (.A(_01421_),
    .B(_01483_),
    .X(_01504_));
 sky130_fd_sc_hd__xnor2_1 _09354_ (.A(_01350_),
    .B(_01343_),
    .Y(_01505_));
 sky130_fd_sc_hd__o211ai_1 _09355_ (.A1(_01484_),
    .A2(_01504_),
    .B1(_01505_),
    .C1(net401),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_01343_),
    .B(_01504_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand2_1 _09357_ (.A(_01290_),
    .B(_01484_),
    .Y(_01508_));
 sky130_fd_sc_hd__a21o_1 _09358_ (.A1(_01507_),
    .A2(_01508_),
    .B1(net401),
    .X(_01509_));
 sky130_fd_sc_hd__and3_1 _09359_ (.A(_01502_),
    .B(_01506_),
    .C(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_01247_),
    .B(_01287_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _09361_ (.A(_01307_),
    .B(_01311_),
    .Y(_01512_));
 sky130_fd_sc_hd__a211oi_2 _09362_ (.A1(_01377_),
    .A2(_01379_),
    .B1(_01319_),
    .C1(_01511_),
    .Y(_01513_));
 sky130_fd_sc_hd__a311o_2 _09363_ (.A1(_01511_),
    .A2(_01512_),
    .A3(_01384_),
    .B1(_01494_),
    .C1(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__a21oi_1 _09364_ (.A1(_01497_),
    .A2(_01510_),
    .B1(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__and3_1 _09365_ (.A(_01496_),
    .B(_01503_),
    .C(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_07420_),
    .B(_01421_),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _09367_ (.A(_07420_),
    .B(_00568_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor3_1 _09368_ (.A(_07359_),
    .B(_07361_),
    .C(_00587_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor3_1 _09369_ (.A(_07342_),
    .B(_07344_),
    .C(_01177_),
    .Y(_01520_));
 sky130_fd_sc_hd__nor2_2 _09370_ (.A(_01073_),
    .B(_07290_),
    .Y(_07294_));
 sky130_fd_sc_hd__nor3_1 _09371_ (.A(_07296_),
    .B(_07304_),
    .C(_07303_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(_01010_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__mux2_4 _09373_ (.A0(_07294_),
    .A1(_01522_),
    .S(_01108_),
    .X(_07323_));
 sky130_fd_sc_hd__nor3_1 _09374_ (.A(_07325_),
    .B(_07327_),
    .C(_01077_),
    .Y(_01523_));
 sky130_fd_sc_hd__nor3_1 _09375_ (.A(_01078_),
    .B(_01235_),
    .C(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__a21o_1 _09376_ (.A1(_01235_),
    .A2(_07323_),
    .B1(_01524_),
    .X(_07340_));
 sky130_fd_sc_hd__nand2_1 _09377_ (.A(_01315_),
    .B(_07340_),
    .Y(_01525_));
 sky130_fd_sc_hd__o31ai_2 _09378_ (.A1(_01178_),
    .A2(_01315_),
    .A3(_01520_),
    .B1(_01525_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand2_1 _09379_ (.A(net17),
    .B(_07357_),
    .Y(_01526_));
 sky130_fd_sc_hd__o31ai_2 _09380_ (.A1(_00588_),
    .A2(net17),
    .A3(_01519_),
    .B1(_01526_),
    .Y(_07376_));
 sky130_fd_sc_hd__nor3_1 _09381_ (.A(_07378_),
    .B(_07380_),
    .C(_01347_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _09382_ (.A(_01348_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__mux2i_4 _09383_ (.A0(_07376_),
    .A1(_01528_),
    .S(_01390_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_2 _09384_ (.A(_01427_),
    .B(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__xnor2_4 _09385_ (.A(_07398_),
    .B(_01481_),
    .Y(_01531_));
 sky130_fd_sc_hd__mux2i_4 _09386_ (.A0(_01530_),
    .A1(_01531_),
    .S(_01497_),
    .Y(_01532_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(_01517_),
    .A1(_01518_),
    .S(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__or2_1 _09388_ (.A(_00594_),
    .B(_01532_),
    .X(_01534_));
 sky130_fd_sc_hd__and3_1 _09389_ (.A(_01516_),
    .B(_01533_),
    .C(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__buf_4 _09390_ (.A(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__o211ai_1 _09391_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01461_),
    .C1(_01435_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _09392_ (.A(_01472_),
    .B(_01475_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _09393_ (.A(_01427_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_2 _09394_ (.A(_01537_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__o21a_1 _09395_ (.A1(_01271_),
    .A2(_01449_),
    .B1(_01453_),
    .X(_01541_));
 sky130_fd_sc_hd__a21o_1 _09396_ (.A1(_01541_),
    .A2(_01458_),
    .B1(_01447_),
    .X(_01542_));
 sky130_fd_sc_hd__a211oi_1 _09397_ (.A1(_01386_),
    .A2(_01375_),
    .B1(_01473_),
    .C1(_01437_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_1 _09398_ (.A1(_01473_),
    .A2(_01437_),
    .B1(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__a21o_1 _09399_ (.A1(net27),
    .A2(_01542_),
    .B1(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__nand3_1 _09400_ (.A(_01490_),
    .B(_01544_),
    .C(_01542_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(_01336_),
    .B(_01337_),
    .Y(_01547_));
 sky130_fd_sc_hd__o21ai_0 _09402_ (.A1(_01375_),
    .A2(_01437_),
    .B1(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__a21oi_1 _09403_ (.A1(_01547_),
    .A2(_01437_),
    .B1(_01338_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(_01386_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__a21oi_1 _09405_ (.A1(_01438_),
    .A2(_01548_),
    .B1(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__a21boi_2 _09406_ (.A1(_01545_),
    .A2(_01546_),
    .B1_N(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _09407_ (.A(_01455_),
    .B(_01456_),
    .Y(_01553_));
 sky130_fd_sc_hd__o21a_1 _09408_ (.A1(net27),
    .A2(_01494_),
    .B1(_01272_),
    .X(_01554_));
 sky130_fd_sc_hd__o221ai_4 _09409_ (.A1(_01472_),
    .A2(_01475_),
    .B1(_01486_),
    .B2(net401),
    .C1(_01489_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(_01272_),
    .B(_01553_),
    .Y(_01556_));
 sky130_fd_sc_hd__a211o_1 _09411_ (.A1(_01493_),
    .A2(_01555_),
    .B1(_01556_),
    .C1(_01447_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _09412_ (.A(net10),
    .B(_01287_),
    .Y(_01558_));
 sky130_fd_sc_hd__a211oi_1 _09413_ (.A1(_01341_),
    .A2(_01445_),
    .B1(_01493_),
    .C1(_01271_),
    .Y(_01559_));
 sky130_fd_sc_hd__o21ai_0 _09414_ (.A1(_01558_),
    .A2(_01559_),
    .B1(_01454_),
    .Y(_01560_));
 sky130_fd_sc_hd__xnor2_1 _09415_ (.A(_01457_),
    .B(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__o211a_2 _09416_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01557_),
    .C1(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__o21ai_4 _09417_ (.A1(_01540_),
    .A2(_01552_),
    .B1(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hd__or2_1 _09418_ (.A(_01399_),
    .B(_01401_),
    .X(_01564_));
 sky130_fd_sc_hd__o2bb2ai_1 _09419_ (.A1_N(_01435_),
    .A2_N(_01427_),
    .B1(_01401_),
    .B2(_01399_),
    .Y(_01565_));
 sky130_fd_sc_hd__o22ai_2 _09420_ (.A1(_01441_),
    .A2(_01442_),
    .B1(_01447_),
    .B2(_01460_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_2 _09421_ (.A(_01566_),
    .B(_01555_),
    .Y(_01567_));
 sky130_fd_sc_hd__mux2i_2 _09422_ (.A0(_01564_),
    .A1(_01565_),
    .S(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__o21a_1 _09423_ (.A1(_07418_),
    .A2(_07417_),
    .B1(_07416_),
    .X(_01569_));
 sky130_fd_sc_hd__o21a_1 _09424_ (.A1(_07415_),
    .A2(_01569_),
    .B1(_07413_),
    .X(_01570_));
 sky130_fd_sc_hd__o21a_1 _09425_ (.A1(_07412_),
    .A2(_01570_),
    .B1(_07430_),
    .X(_01571_));
 sky130_fd_sc_hd__o21a_1 _09426_ (.A1(_07429_),
    .A2(_01571_),
    .B1(_07427_),
    .X(_01572_));
 sky130_fd_sc_hd__o21a_2 _09427_ (.A1(_07426_),
    .A2(_01572_),
    .B1(_07424_),
    .X(_01573_));
 sky130_fd_sc_hd__o21ai_4 _09428_ (.A1(_01573_),
    .A2(_07423_),
    .B1(_07421_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor3_4 _09429_ (.A(_01421_),
    .B(_01531_),
    .C(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__xor2_2 _09430_ (.A(_07398_),
    .B(_01481_),
    .X(_01576_));
 sky130_fd_sc_hd__nor3_4 _09431_ (.A(_01574_),
    .B(_01576_),
    .C(_00568_),
    .Y(_01577_));
 sky130_fd_sc_hd__o21ai_4 _09432_ (.A1(_01577_),
    .A2(_01575_),
    .B1(_01497_),
    .Y(_01578_));
 sky130_fd_sc_hd__mux2i_2 _09433_ (.A0(_01420_),
    .A1(_01425_),
    .S(net401),
    .Y(_01579_));
 sky130_fd_sc_hd__inv_1 _09434_ (.A(_01529_),
    .Y(_07396_));
 sky130_fd_sc_hd__o21ai_0 _09435_ (.A1(_01579_),
    .A2(_07396_),
    .B1(_01421_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand3_1 _09436_ (.A(_00568_),
    .B(_01427_),
    .C(_01529_),
    .Y(_01581_));
 sky130_fd_sc_hd__a211o_2 _09437_ (.A1(_01580_),
    .A2(_01581_),
    .B1(_01497_),
    .C1(_01574_),
    .X(_01582_));
 sky130_fd_sc_hd__o211ai_1 _09438_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01427_),
    .C1(_01435_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _09439_ (.A(_01447_),
    .B(_01460_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _09440_ (.A(_01441_),
    .B(_01442_),
    .Y(_01585_));
 sky130_fd_sc_hd__o21a_1 _09441_ (.A1(_01584_),
    .A2(_01555_),
    .B1(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__a21oi_2 _09442_ (.A1(_01567_),
    .A2(_01583_),
    .B1(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand4b_2 _09443_ (.A_N(_01568_),
    .B(_01578_),
    .C(_01582_),
    .D(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _09444_ (.A(_01563_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__or3_1 _09445_ (.A(_07421_),
    .B(_07423_),
    .C(_01573_),
    .X(_01590_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_01574_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__a21boi_2 _09447_ (.A1(_01536_),
    .A2(_01589_),
    .B1_N(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__a21oi_4 _09448_ (.A1(_01564_),
    .A2(_01567_),
    .B1(_01435_),
    .Y(_01593_));
 sky130_fd_sc_hd__and2_0 _09449_ (.A(_01591_),
    .B(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__nand3_1 _09450_ (.A(_01496_),
    .B(_01503_),
    .C(_01515_),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(_01582_),
    .B(_01578_),
    .Y(_01596_));
 sky130_fd_sc_hd__o21ai_1 _09452_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01435_),
    .Y(_01597_));
 sky130_fd_sc_hd__or2_0 _09453_ (.A(_01597_),
    .B(_01586_),
    .X(_01598_));
 sky130_fd_sc_hd__nand4_1 _09454_ (.A(_07418_),
    .B(_07424_),
    .C(_07427_),
    .D(_07430_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand3_1 _09455_ (.A(_07413_),
    .B(_07416_),
    .C(_07421_),
    .Y(_01600_));
 sky130_fd_sc_hd__nor3_2 _09456_ (.A(_01114_),
    .B(_01599_),
    .C(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_1 _09457_ (.A(_07420_),
    .B(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__clkbuf_4 _09458_ (.A(_00594_),
    .X(_01603_));
 sky130_fd_sc_hd__o21ai_1 _09459_ (.A1(_00568_),
    .A2(_01602_),
    .B1(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _09460_ (.A(_01531_),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__o21ai_0 _09461_ (.A1(_01579_),
    .A2(_07396_),
    .B1(_01604_),
    .Y(_01606_));
 sky130_fd_sc_hd__o2111a_2 _09462_ (.A1(_01399_),
    .A2(_01401_),
    .B1(_01461_),
    .C1(_01435_),
    .D1(_01490_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2i_1 _09463_ (.A0(_01605_),
    .A1(_01606_),
    .S(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor3_1 _09464_ (.A(_07362_),
    .B(_07364_),
    .C(_00586_),
    .Y(_01609_));
 sky130_fd_sc_hd__nor3_1 _09465_ (.A(_07345_),
    .B(_07347_),
    .C(_01176_),
    .Y(_01610_));
 sky130_fd_sc_hd__a21oi_2 _09466_ (.A1(_01057_),
    .A2(_01113_),
    .B1(_07304_),
    .Y(_07326_));
 sky130_fd_sc_hd__nor3_1 _09467_ (.A(_07330_),
    .B(_07328_),
    .C(_07329_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _09468_ (.A(_01077_),
    .B(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(_07326_),
    .A1(_01612_),
    .S(_01173_),
    .X(_07343_));
 sky130_fd_sc_hd__nand2_1 _09470_ (.A(_01315_),
    .B(_07343_),
    .Y(_01613_));
 sky130_fd_sc_hd__o31ai_2 _09471_ (.A1(_01177_),
    .A2(_01315_),
    .A3(_01610_),
    .B1(_01613_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(net17),
    .B(_07360_),
    .Y(_01614_));
 sky130_fd_sc_hd__o31ai_1 _09473_ (.A1(_00587_),
    .A2(net17),
    .A3(_01609_),
    .B1(_01614_),
    .Y(_07379_));
 sky130_fd_sc_hd__nor3_1 _09474_ (.A(_07381_),
    .B(_07383_),
    .C(_01346_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _09475_ (.A(_01347_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__mux2_1 _09476_ (.A0(_07379_),
    .A1(_01616_),
    .S(_01426_),
    .X(_07399_));
 sky130_fd_sc_hd__nor3_1 _09477_ (.A(_07401_),
    .B(_07403_),
    .C(_01479_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_01480_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__buf_6 _09479_ (.A(_01497_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(_07399_),
    .A1(_01618_),
    .S(_01619_),
    .X(_07419_));
 sky130_fd_sc_hd__nor2_1 _09481_ (.A(_01421_),
    .B(_01602_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _09482_ (.A(_01576_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__nand3_1 _09483_ (.A(_01427_),
    .B(_01529_),
    .C(_01620_),
    .Y(_01622_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(_01621_),
    .A1(_01622_),
    .S(_01607_),
    .X(_01623_));
 sky130_fd_sc_hd__or4b_1 _09485_ (.A(_01598_),
    .B(_01608_),
    .C(_07419_),
    .D_N(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__nor4_1 _09486_ (.A(_01595_),
    .B(_01563_),
    .C(_01596_),
    .D(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__a31oi_4 _09487_ (.A1(_01619_),
    .A2(_01500_),
    .A3(_01501_),
    .B1(_01502_),
    .Y(_01626_));
 sky130_fd_sc_hd__a21o_1 _09488_ (.A1(_01619_),
    .A2(_01510_),
    .B1(_01514_),
    .X(_01627_));
 sky130_fd_sc_hd__o21ai_1 _09489_ (.A1(_01540_),
    .A2(_01552_),
    .B1(_01496_),
    .Y(_01628_));
 sky130_fd_sc_hd__clkbuf_4 _09490_ (.A(_01421_),
    .X(_01629_));
 sky130_fd_sc_hd__nor4_1 _09491_ (.A(_01629_),
    .B(_01114_),
    .C(_01599_),
    .D(_01600_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _09492_ (.A(_01576_),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand3_1 _09493_ (.A(_01629_),
    .B(_01531_),
    .C(_01601_),
    .Y(_01632_));
 sky130_fd_sc_hd__buf_6 _09494_ (.A(_01607_),
    .X(_01633_));
 sky130_fd_sc_hd__a21oi_1 _09495_ (.A1(_01631_),
    .A2(_01632_),
    .B1(net20),
    .Y(_01634_));
 sky130_fd_sc_hd__o211ai_1 _09496_ (.A1(_01579_),
    .A2(_07396_),
    .B1(_01601_),
    .C1(_01629_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_01427_),
    .B(_01529_),
    .C(_01630_),
    .Y(_01636_));
 sky130_fd_sc_hd__a21oi_1 _09498_ (.A1(_01635_),
    .A2(_01636_),
    .B1(net39),
    .Y(_01637_));
 sky130_fd_sc_hd__o21ai_0 _09499_ (.A1(_01634_),
    .A2(_01637_),
    .B1(_01562_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor4_2 _09500_ (.A(_01626_),
    .B(_01627_),
    .C(_01628_),
    .D(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__or3_2 _09501_ (.A(_01594_),
    .B(_01625_),
    .C(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__nand4_1 _09502_ (.A(_07433_),
    .B(_07441_),
    .C(_07447_),
    .D(_07450_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand3_1 _09503_ (.A(_07436_),
    .B(_07439_),
    .C(_07444_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor3_1 _09504_ (.A(_01114_),
    .B(_01641_),
    .C(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__o211a_1 _09505_ (.A1(_01592_),
    .A2(_01640_),
    .B1(_00569_),
    .C1(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__nand3_4 _09506_ (.A(_01516_),
    .B(_01533_),
    .C(_01534_),
    .Y(_01645_));
 sky130_fd_sc_hd__o31ai_4 _09507_ (.A1(_01563_),
    .A2(_01588_),
    .A3(_01645_),
    .B1(_01591_),
    .Y(_01646_));
 sky130_fd_sc_hd__nor3_2 _09508_ (.A(_01594_),
    .B(_01625_),
    .C(_01639_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand4_2 _09509_ (.A(_01629_),
    .B(_01643_),
    .C(_01646_),
    .D(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__o21ai_1 _09510_ (.A1(net401),
    .A2(_01486_),
    .B1(_01489_),
    .Y(_01649_));
 sky130_fd_sc_hd__xor2_1 _09511_ (.A(_01649_),
    .B(_01499_),
    .X(_01650_));
 sky130_fd_sc_hd__nor2_4 _09512_ (.A(net20),
    .B(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__nor2_2 _09513_ (.A(_01514_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand3b_4 _09514_ (.A_N(_01644_),
    .B(_01648_),
    .C(_01652_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _09515_ (.A(_01568_),
    .B(_01593_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _09516_ (.A(_01597_),
    .B(_01586_),
    .Y(_01655_));
 sky130_fd_sc_hd__o21a_1 _09517_ (.A1(_01540_),
    .A2(_01552_),
    .B1(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__and3_4 _09518_ (.A(_01578_),
    .B(_01582_),
    .C(_01562_),
    .X(_01657_));
 sky130_fd_sc_hd__and2_4 _09519_ (.A(_01656_),
    .B(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__clkbuf_2 clone7 (.A(_02624_),
    .X(net7));
 sky130_fd_sc_hd__o21a_1 _09521_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01557_),
    .X(_01660_));
 sky130_fd_sc_hd__and2_0 _09522_ (.A(_01496_),
    .B(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__nor2b_1 _09523_ (.A(_01496_),
    .B_N(_01660_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2b_1 _09524_ (.A(_07420_),
    .B_N(_01574_),
    .Y(_01663_));
 sky130_fd_sc_hd__or2_0 _09525_ (.A(_01421_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__o21ai_0 _09526_ (.A1(_00568_),
    .A2(_01663_),
    .B1(_00594_),
    .Y(_01665_));
 sky130_fd_sc_hd__o21ai_0 _09527_ (.A1(_01579_),
    .A2(_07396_),
    .B1(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__o211ai_2 _09528_ (.A1(_01530_),
    .A2(_01664_),
    .B1(_01666_),
    .C1(_01607_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _09529_ (.A(_01531_),
    .B(_01665_),
    .Y(_01668_));
 sky130_fd_sc_hd__o211ai_2 _09530_ (.A1(_01531_),
    .A2(_01664_),
    .B1(_01668_),
    .C1(net39),
    .Y(_01669_));
 sky130_fd_sc_hd__a211oi_2 _09531_ (.A1(_01667_),
    .A2(_01669_),
    .B1(_01626_),
    .C1(_01627_),
    .Y(_01670_));
 sky130_fd_sc_hd__mux2_1 _09532_ (.A0(_01661_),
    .A1(_01662_),
    .S(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__o22a_1 _09533_ (.A1(_01589_),
    .A2(_01654_),
    .B1(_01658_),
    .B2(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__a21o_1 _09534_ (.A1(_01654_),
    .A2(_01671_),
    .B1(_01536_),
    .X(_01673_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_01672_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__a21oi_1 _09536_ (.A1(_01541_),
    .A2(_01458_),
    .B1(_01447_),
    .Y(_01675_));
 sky130_fd_sc_hd__nor4_1 _09537_ (.A(_01555_),
    .B(_01544_),
    .C(_01540_),
    .D(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__o21ai_0 _09538_ (.A1(_01555_),
    .A2(_01675_),
    .B1(_01544_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand2b_1 _09539_ (.A_N(_01676_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__clkbuf_4 _09540_ (.A(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__nor2_2 _09541_ (.A(_01563_),
    .B(_01596_),
    .Y(_01680_));
 sky130_fd_sc_hd__xnor2_1 _09542_ (.A(_00569_),
    .B(_01532_),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_01681_),
    .B(_01601_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _09544_ (.A(_01682_),
    .B(_01655_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_01561_),
    .B(_01660_),
    .Y(_01684_));
 sky130_fd_sc_hd__a221oi_4 _09546_ (.A1(net39),
    .A2(_01510_),
    .B1(_01582_),
    .B2(_01578_),
    .C1(_01626_),
    .Y(_01685_));
 sky130_fd_sc_hd__xnor2_1 _09547_ (.A(_01551_),
    .B(_01676_),
    .Y(_01686_));
 sky130_fd_sc_hd__o41a_1 _09548_ (.A1(_01684_),
    .A2(_01645_),
    .A3(_01685_),
    .A4(_01679_),
    .B1(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__a31o_1 _09549_ (.A1(_01680_),
    .A2(_01536_),
    .A3(_01683_),
    .B1(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__and2_0 _09550_ (.A(_01582_),
    .B(_01578_),
    .X(_01689_));
 sky130_fd_sc_hd__a211oi_1 _09551_ (.A1(_01689_),
    .A2(_01656_),
    .B1(_01685_),
    .C1(_01684_),
    .Y(_01690_));
 sky130_fd_sc_hd__o21ai_0 _09552_ (.A1(_01566_),
    .A2(_01555_),
    .B1(_01576_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand4_1 _09553_ (.A(_01461_),
    .B(_01427_),
    .C(net27),
    .D(_01529_),
    .Y(_01692_));
 sky130_fd_sc_hd__a311oi_1 _09554_ (.A1(_01604_),
    .A2(_01691_),
    .A3(_01692_),
    .B1(_01586_),
    .C1(_01597_),
    .Y(_01693_));
 sky130_fd_sc_hd__nand4_1 _09555_ (.A(_01623_),
    .B(_01582_),
    .C(_01578_),
    .D(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__o211ai_1 _09556_ (.A1(_01563_),
    .A2(_01694_),
    .B1(_01670_),
    .C1(_01661_),
    .Y(_01695_));
 sky130_fd_sc_hd__a41oi_1 _09557_ (.A1(_01272_),
    .A2(_01553_),
    .A3(_01537_),
    .A4(net27),
    .B1(_01561_),
    .Y(_01696_));
 sky130_fd_sc_hd__a21oi_1 _09558_ (.A1(net27),
    .A2(_01542_),
    .B1(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _09559_ (.A(_01540_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__a22o_1 _09560_ (.A1(_01536_),
    .A2(_01690_),
    .B1(_01695_),
    .B2(_01698_),
    .X(_01699_));
 sky130_fd_sc_hd__a21o_1 _09561_ (.A1(_01680_),
    .A2(_01536_),
    .B1(_01587_),
    .X(_01700_));
 sky130_fd_sc_hd__and4_1 _09562_ (.A(_01598_),
    .B(_01533_),
    .C(_01534_),
    .D(_01587_),
    .X(_01701_));
 sky130_fd_sc_hd__nand3_1 _09563_ (.A(_01516_),
    .B(_01680_),
    .C(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand3b_1 _09564_ (.A_N(_01699_),
    .B(_01700_),
    .C(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__or4_1 _09565_ (.A(_01674_),
    .B(_01679_),
    .C(_01688_),
    .D(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__buf_2 _09566_ (.A(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__or2_0 _09567_ (.A(_01653_),
    .B(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__buf_4 _09568_ (.A(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__o21a_1 _09569_ (.A1(_07441_),
    .A2(_07440_),
    .B1(_07439_),
    .X(_01708_));
 sky130_fd_sc_hd__o21a_1 _09570_ (.A1(_07438_),
    .A2(_01708_),
    .B1(_07436_),
    .X(_01709_));
 sky130_fd_sc_hd__o21a_1 _09571_ (.A1(_07435_),
    .A2(_01709_),
    .B1(_07433_),
    .X(_01710_));
 sky130_fd_sc_hd__o21a_1 _09572_ (.A1(_07432_),
    .A2(_01710_),
    .B1(_07450_),
    .X(_01711_));
 sky130_fd_sc_hd__o21a_1 _09573_ (.A1(_07449_),
    .A2(_01711_),
    .B1(_07447_),
    .X(_01712_));
 sky130_fd_sc_hd__o21ai_2 _09574_ (.A1(_01712_),
    .A2(_07446_),
    .B1(_07444_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2b_2 _09575_ (.A_N(_07443_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__o211ai_4 _09576_ (.A1(_01592_),
    .A2(_01640_),
    .B1(_01714_),
    .C1(_00569_),
    .Y(_01715_));
 sky130_fd_sc_hd__nor2b_4 _09577_ (.A(_07443_),
    .B_N(_01713_),
    .Y(_01716_));
 sky130_fd_sc_hd__o21ai_2 _09578_ (.A1(_00569_),
    .A2(_01716_),
    .B1(_01603_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand3_2 _09579_ (.A(_01646_),
    .B(_01647_),
    .C(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(_00569_),
    .B(_01663_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21boi_1 _09581_ (.A1(_01536_),
    .A2(_01658_),
    .B1_N(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__xor2_2 _09582_ (.A(_01532_),
    .B(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__nand2_1 _09583_ (.A(_01667_),
    .B(_01669_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(net39),
    .B(_01501_),
    .Y(_01723_));
 sky130_fd_sc_hd__xnor2_2 _09585_ (.A(_01502_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_2 _09586_ (.A(_01722_),
    .B(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__a21o_1 _09587_ (.A1(_01536_),
    .A2(_01658_),
    .B1(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__o21a_2 _09588_ (.A1(_01722_),
    .A2(_01724_),
    .B1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__nand4_4 _09589_ (.A(_01715_),
    .B(_01718_),
    .C(_01721_),
    .D(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__and2_0 _09590_ (.A(_01651_),
    .B(_01725_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_4 _09591_ (.A(_01536_),
    .X(_01730_));
 sky130_fd_sc_hd__a211o_1 _09592_ (.A1(_01730_),
    .A2(_01658_),
    .B1(_01651_),
    .C1(_01725_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2b_2 _09593_ (.A(_01729_),
    .B_N(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_4 _09594_ (.A(_01658_),
    .B(_01730_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand2b_1 _09595_ (.A_N(_01671_),
    .B(net33),
    .Y(_01734_));
 sky130_fd_sc_hd__a311oi_4 _09596_ (.A1(_01511_),
    .A2(_01512_),
    .A3(_01384_),
    .B1(_01494_),
    .C1(_01513_),
    .Y(_01735_));
 sky130_fd_sc_hd__nor2_1 _09597_ (.A(_01649_),
    .B(_01499_),
    .Y(_01736_));
 sky130_fd_sc_hd__o21ai_2 _09598_ (.A1(_01462_),
    .A2(_01538_),
    .B1(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand3_1 _09599_ (.A(_01735_),
    .B(_01651_),
    .C(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__o21ai_0 _09600_ (.A1(_01735_),
    .A2(_01737_),
    .B1(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__a31oi_2 _09601_ (.A1(_01735_),
    .A2(_01725_),
    .A3(_01737_),
    .B1(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__o311ai_4 _09602_ (.A1(_01735_),
    .A2(_01651_),
    .A3(_01725_),
    .B1(_01740_),
    .C1(net33),
    .Y(_01741_));
 sky130_fd_sc_hd__nand3_1 _09603_ (.A(_01732_),
    .B(_01734_),
    .C(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__or3_2 _09604_ (.A(_01699_),
    .B(_01728_),
    .C(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__nor3_1 _09605_ (.A(_07404_),
    .B(_07406_),
    .C(_01478_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor3_4 _09606_ (.A(_01439_),
    .B(_01474_),
    .C(_01473_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor3_1 _09607_ (.A(_07384_),
    .B(_07386_),
    .C(_01345_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor3_1 _09608_ (.A(_07365_),
    .B(_07367_),
    .C(_00585_),
    .Y(_01747_));
 sky130_fd_sc_hd__nor3_1 _09609_ (.A(_07350_),
    .B(_07348_),
    .C(_07349_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_8 _09610_ (.A(_07330_),
    .B(_01235_),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_2 _09611_ (.A(_01315_),
    .B(_07346_),
    .Y(_01749_));
 sky130_fd_sc_hd__o31ai_4 _09612_ (.A1(_01176_),
    .A2(_01315_),
    .A3(_01748_),
    .B1(_01749_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand2_1 _09613_ (.A(_01492_),
    .B(_07363_),
    .Y(_01750_));
 sky130_fd_sc_hd__o31ai_1 _09614_ (.A1(_00586_),
    .A2(_01492_),
    .A3(_01747_),
    .B1(_01750_),
    .Y(_07382_));
 sky130_fd_sc_hd__nand2_1 _09615_ (.A(_01745_),
    .B(_07382_),
    .Y(_01751_));
 sky130_fd_sc_hd__o31ai_1 _09616_ (.A1(_01346_),
    .A2(_01745_),
    .A3(_01746_),
    .B1(_01751_),
    .Y(_07402_));
 sky130_fd_sc_hd__nand2_1 _09617_ (.A(net20),
    .B(_07402_),
    .Y(_01752_));
 sky130_fd_sc_hd__o31ai_4 _09618_ (.A1(_01479_),
    .A2(net20),
    .A3(_01744_),
    .B1(_01752_),
    .Y(_07422_));
 sky130_fd_sc_hd__nor3_1 _09619_ (.A(_07424_),
    .B(_07426_),
    .C(_01572_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _09620_ (.A(_01573_),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__mux2i_4 _09621_ (.A0(_07422_),
    .A1(_01754_),
    .S(_01733_),
    .Y(_01755_));
 sky130_fd_sc_hd__o21ai_0 _09622_ (.A1(_01573_),
    .A2(_01753_),
    .B1(_00569_),
    .Y(_01756_));
 sky130_fd_sc_hd__nand2_1 _09623_ (.A(_01629_),
    .B(_01754_),
    .Y(_01757_));
 sky130_fd_sc_hd__o21a_1 _09624_ (.A1(_07464_),
    .A2(_07463_),
    .B1(_07462_),
    .X(_01758_));
 sky130_fd_sc_hd__o21a_1 _09625_ (.A1(_07461_),
    .A2(_01758_),
    .B1(_07459_),
    .X(_01759_));
 sky130_fd_sc_hd__o21a_1 _09626_ (.A1(_07458_),
    .A2(_01759_),
    .B1(_07456_),
    .X(_01760_));
 sky130_fd_sc_hd__o21a_1 _09627_ (.A1(_07455_),
    .A2(_01760_),
    .B1(_07453_),
    .X(_01761_));
 sky130_fd_sc_hd__o21a_1 _09628_ (.A1(_07452_),
    .A2(_01761_),
    .B1(_07470_),
    .X(_01762_));
 sky130_fd_sc_hd__o21ai_1 _09629_ (.A1(_01762_),
    .A2(_07469_),
    .B1(_07467_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2b_4 _09630_ (.A(_07466_),
    .B_N(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__clkbuf_2 clone18 (.A(_02749_),
    .X(net18));
 sky130_fd_sc_hd__a221oi_1 _09632_ (.A1(_01730_),
    .A2(_01658_),
    .B1(_01756_),
    .B2(_01757_),
    .C1(_01764_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand3b_4 _09633_ (.A_N(_01764_),
    .B(_07422_),
    .C(_01629_),
    .Y(_01767_));
 sky130_fd_sc_hd__or3_1 _09634_ (.A(_01629_),
    .B(_01764_),
    .C(_07422_),
    .X(_01768_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_01656_),
    .B(_01657_),
    .Y(_01769_));
 sky130_fd_sc_hd__a211oi_2 _09636_ (.A1(_01767_),
    .A2(_01768_),
    .B1(_01645_),
    .C1(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_2 _09637_ (.A(_01770_),
    .B(_01766_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand2_2 _09638_ (.A(_01646_),
    .B(_01647_),
    .Y(_01772_));
 sky130_fd_sc_hd__o211ai_4 _09639_ (.A1(_01603_),
    .A2(_01755_),
    .B1(_01771_),
    .C1(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__o21ai_1 _09640_ (.A1(_01722_),
    .A2(_01724_),
    .B1(_01726_),
    .Y(_01774_));
 sky130_fd_sc_hd__and3_1 _09641_ (.A(_01715_),
    .B(_01718_),
    .C(_01721_),
    .X(_01775_));
 sky130_fd_sc_hd__or3_1 _09642_ (.A(_01651_),
    .B(_01774_),
    .C(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__nor2_1 _09643_ (.A(_01592_),
    .B(_01640_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand3_1 _09644_ (.A(_01532_),
    .B(_01716_),
    .C(_01719_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _09645_ (.A(_01532_),
    .B(_01714_),
    .Y(_01779_));
 sky130_fd_sc_hd__nand4_1 _09646_ (.A(_01730_),
    .B(_01656_),
    .C(_01657_),
    .D(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _09647_ (.A(_01657_),
    .B(_01778_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _09648_ (.A(_01656_),
    .B(_01778_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor3_1 _09649_ (.A(_01532_),
    .B(_01714_),
    .C(_01719_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor3_1 _09650_ (.A(_01781_),
    .B(_01782_),
    .C(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o211ai_1 _09651_ (.A1(_01730_),
    .A2(_01778_),
    .B1(_01780_),
    .C1(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__buf_4 _09652_ (.A(_01629_),
    .X(_01786_));
 sky130_fd_sc_hd__a31oi_1 _09653_ (.A1(_01603_),
    .A2(_01777_),
    .A3(_01785_),
    .B1(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor4_1 _09654_ (.A(_01603_),
    .B(_01592_),
    .C(_01640_),
    .D(_01714_),
    .Y(_01788_));
 sky130_fd_sc_hd__a21oi_1 _09655_ (.A1(_01646_),
    .A2(_01647_),
    .B1(_01716_),
    .Y(_01789_));
 sky130_fd_sc_hd__o21ai_0 _09656_ (.A1(_01788_),
    .A2(_01789_),
    .B1(_01721_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _09657_ (.A(net20),
    .B(_01531_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _09658_ (.A(net39),
    .B(_01530_),
    .Y(_01792_));
 sky130_fd_sc_hd__o211ai_1 _09659_ (.A1(_01645_),
    .A2(_01769_),
    .B1(_01719_),
    .C1(_01532_),
    .Y(_01793_));
 sky130_fd_sc_hd__o311a_1 _09660_ (.A1(_01791_),
    .A2(_01792_),
    .A3(_01720_),
    .B1(_01793_),
    .C1(_01714_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2i_1 _09661_ (.A0(_01785_),
    .A1(_01794_),
    .S(_01777_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_2 _09662_ (.A(_07446_),
    .B(_01712_),
    .Y(_01796_));
 sky130_fd_sc_hd__xor2_2 _09663_ (.A(_07444_),
    .B(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__xnor2_4 _09664_ (.A(_07444_),
    .B(_01796_),
    .Y(_01798_));
 sky130_fd_sc_hd__xnor2_1 _09665_ (.A(_00569_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__o22ai_2 _09666_ (.A1(_01603_),
    .A2(_01797_),
    .B1(_01799_),
    .B2(_01764_),
    .Y(_01800_));
 sky130_fd_sc_hd__a221o_2 _09667_ (.A1(_01787_),
    .A2(_01790_),
    .B1(_01795_),
    .B2(_01786_),
    .C1(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__o32ai_4 _09668_ (.A1(_01707_),
    .A2(_01773_),
    .A3(_01743_),
    .B1(_01776_),
    .B2(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(_01496_),
    .B(_01652_),
    .Y(_01803_));
 sky130_fd_sc_hd__o22a_1 _09670_ (.A1(_01496_),
    .A2(_01670_),
    .B1(_01726_),
    .B2(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__nand2_1 _09671_ (.A(_01741_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2b_2 _09672_ (.A_N(_01729_),
    .B(_01731_),
    .Y(_01806_));
 sky130_fd_sc_hd__xnor2_1 _09673_ (.A(_01735_),
    .B(_01737_),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(_01496_),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__o21ai_0 _09675_ (.A1(_01806_),
    .A2(_01808_),
    .B1(_01804_),
    .Y(_01809_));
 sky130_fd_sc_hd__and4_4 _09676_ (.A(_01715_),
    .B(_01727_),
    .C(_01721_),
    .D(_01718_),
    .X(_01810_));
 sky130_fd_sc_hd__buf_4 _09677_ (.A(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2i_1 _09678_ (.A0(_01805_),
    .A1(_01809_),
    .S(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _09679_ (.A(_01806_),
    .B(_01808_),
    .Y(_01813_));
 sky130_fd_sc_hd__a211oi_1 _09680_ (.A1(_01705_),
    .A2(_01813_),
    .B1(_01653_),
    .C1(_01728_),
    .Y(_01814_));
 sky130_fd_sc_hd__and3b_1 _09681_ (.A_N(_01644_),
    .B(_01648_),
    .C(_01652_),
    .X(_01815_));
 sky130_fd_sc_hd__clkinvlp_4 _09682_ (.A(_01741_),
    .Y(_01816_));
 sky130_fd_sc_hd__a32oi_1 _09683_ (.A1(_01815_),
    .A2(_01811_),
    .A3(_01705_),
    .B1(_01806_),
    .B2(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__o21a_4 _09684_ (.A1(_01812_),
    .A2(_01814_),
    .B1(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__and2_4 _09685_ (.A(_01818_),
    .B(_01802_),
    .X(_01819_));
 sky130_fd_sc_hd__buf_8 _09686_ (.A(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__nor2_1 _09687_ (.A(_01645_),
    .B(_01685_),
    .Y(_01821_));
 sky130_fd_sc_hd__o21ai_1 _09688_ (.A1(_01660_),
    .A2(_01821_),
    .B1(_01695_),
    .Y(_01822_));
 sky130_fd_sc_hd__and2_0 _09689_ (.A(_01730_),
    .B(_01690_),
    .X(_01823_));
 sky130_fd_sc_hd__xor2_1 _09690_ (.A(_01679_),
    .B(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_1 _09691_ (.A(_01822_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__nor3_2 _09692_ (.A(_01699_),
    .B(_01728_),
    .C(_01742_),
    .Y(_01826_));
 sky130_fd_sc_hd__and3_1 _09693_ (.A(_01732_),
    .B(_01734_),
    .C(_01741_),
    .X(_01827_));
 sky130_fd_sc_hd__a21boi_2 _09694_ (.A1(_01811_),
    .A2(_01827_),
    .B1_N(_01699_),
    .Y(_01828_));
 sky130_fd_sc_hd__a21oi_4 _09695_ (.A1(_01707_),
    .A2(_01826_),
    .B1(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_2 _09696_ (.A(_01730_),
    .B(_01589_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _09697_ (.A(_01593_),
    .B(_01639_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand3_1 _09698_ (.A(_01680_),
    .B(_01587_),
    .C(_01730_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _09699_ (.A(_01568_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__o21ai_4 _09700_ (.A1(_01830_),
    .A2(_01831_),
    .B1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__nand3_1 _09701_ (.A(_01672_),
    .B(_01673_),
    .C(_01652_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor3b_1 _09702_ (.A(_01835_),
    .B(_01644_),
    .C_N(_01648_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor3_2 _09703_ (.A(_01679_),
    .B(_01688_),
    .C(_01703_),
    .Y(_01837_));
 sky130_fd_sc_hd__nand4b_4 _09704_ (.A_N(_01836_),
    .B(_01837_),
    .C(_01810_),
    .D(_01827_),
    .Y(_01838_));
 sky130_fd_sc_hd__o211ai_4 _09705_ (.A1(_01834_),
    .A2(_01838_),
    .B1(_01830_),
    .C1(_01593_),
    .Y(_01839_));
 sky130_fd_sc_hd__xor2_4 _09706_ (.A(_01834_),
    .B(_01838_),
    .X(_01840_));
 sky130_fd_sc_hd__a31oi_4 _09707_ (.A1(_01680_),
    .A2(_01730_),
    .A3(_01683_),
    .B1(_01687_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand4_1 _09708_ (.A(_01841_),
    .B(_01700_),
    .C(_01702_),
    .D(_01825_),
    .Y(_01842_));
 sky130_fd_sc_hd__a211oi_4 _09709_ (.A1(_01707_),
    .A2(_01826_),
    .B1(_01828_),
    .C1(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__and3_1 _09710_ (.A(_01839_),
    .B(_01840_),
    .C(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__buf_4 _09711_ (.A(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__clkinvlp_4 _09712_ (.A(_01755_),
    .Y(_07442_));
 sky130_fd_sc_hd__xnor2_1 _09713_ (.A(_00569_),
    .B(_07442_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor4_1 _09714_ (.A(_01653_),
    .B(_01728_),
    .C(_01705_),
    .D(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__a21oi_1 _09715_ (.A1(_01715_),
    .A2(_01718_),
    .B1(_01721_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor3_1 _09716_ (.A(_01775_),
    .B(_01799_),
    .C(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand4_1 _09717_ (.A(_07464_),
    .B(_07453_),
    .C(_07456_),
    .D(_07470_),
    .Y(_01850_));
 sky130_fd_sc_hd__nand3_1 _09718_ (.A(_07459_),
    .B(_07462_),
    .C(_07467_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor3_1 _09719_ (.A(_01114_),
    .B(_01850_),
    .C(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__o21ai_2 _09720_ (.A1(_01847_),
    .A2(_01849_),
    .B1(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__xnor2_1 _09721_ (.A(_01629_),
    .B(_01716_),
    .Y(_01854_));
 sky130_fd_sc_hd__a31oi_2 _09722_ (.A1(_01836_),
    .A2(_01837_),
    .A3(_01811_),
    .B1(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__xnor2_2 _09723_ (.A(_01772_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__or2_2 _09724_ (.A(_01853_),
    .B(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__nand3_1 _09725_ (.A(_01818_),
    .B(_01845_),
    .C(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand4_2 _09726_ (.A(net25),
    .B(_01825_),
    .C(_01829_),
    .D(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_2 _09727_ (.A(_01653_),
    .B(_01705_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor4_2 _09728_ (.A(_01679_),
    .B(_01688_),
    .C(_01860_),
    .D(_01743_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_01679_),
    .B(_01743_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _09730_ (.A(_01841_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_2 _09731_ (.A(_01861_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__xnor2_4 _09732_ (.A(_01859_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__inv_1 _09733_ (.A(_01822_),
    .Y(_01866_));
 sky130_fd_sc_hd__and3_1 _09734_ (.A(_01802_),
    .B(_01818_),
    .C(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__or2_0 _09735_ (.A(_01829_),
    .B(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__buf_2 _09736_ (.A(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__nand3_4 _09737_ (.A(_01839_),
    .B(_01840_),
    .C(_01843_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _09738_ (.A(_01853_),
    .B(_01856_),
    .Y(_01871_));
 sky130_fd_sc_hd__o211ai_4 _09739_ (.A1(_01870_),
    .A2(_01871_),
    .B1(_01867_),
    .C1(_01829_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_2 _09740_ (.A(_01869_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__o211a_1 _09741_ (.A1(_01834_),
    .A2(_01838_),
    .B1(_01830_),
    .C1(_01593_),
    .X(_01874_));
 sky130_fd_sc_hd__a31oi_2 _09742_ (.A1(_01802_),
    .A2(_01818_),
    .A3(_01843_),
    .B1(_01840_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21o_1 _09743_ (.A1(_01707_),
    .A2(_01826_),
    .B1(_01823_),
    .X(_01876_));
 sky130_fd_sc_hd__and3_4 _09744_ (.A(_01836_),
    .B(_01837_),
    .C(_01810_),
    .X(_01877_));
 sky130_fd_sc_hd__buf_6 _09745_ (.A(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__a21o_1 _09746_ (.A1(_01841_),
    .A2(_01743_),
    .B1(net29),
    .X(_01879_));
 sky130_fd_sc_hd__nor2_1 _09747_ (.A(_01679_),
    .B(_01823_),
    .Y(_01880_));
 sky130_fd_sc_hd__a32oi_4 _09748_ (.A1(_01679_),
    .A2(_01841_),
    .A3(_01876_),
    .B1(_01879_),
    .B2(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(_01700_),
    .B(_01702_),
    .Y(_01882_));
 sky130_fd_sc_hd__xor2_2 _09750_ (.A(_01882_),
    .B(_01861_),
    .X(_01883_));
 sky130_fd_sc_hd__nor4_2 _09751_ (.A(_01874_),
    .B(_01875_),
    .C(_01881_),
    .D(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__and3_2 _09752_ (.A(_01869_),
    .B(_01872_),
    .C(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__nand2_8 _09753_ (.A(_01802_),
    .B(_01818_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor3_1 _09754_ (.A(_07447_),
    .B(_07449_),
    .C(_01711_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _09755_ (.A(_01712_),
    .B(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor3_1 _09756_ (.A(_07407_),
    .B(_07409_),
    .C(_01477_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor3_1 _09757_ (.A(_07368_),
    .B(_07370_),
    .C(_07369_),
    .Y(_01890_));
 sky130_fd_sc_hd__nor2_4 _09758_ (.A(_01315_),
    .B(_07350_),
    .Y(_07366_));
 sky130_fd_sc_hd__nand2_2 _09759_ (.A(_01492_),
    .B(_07366_),
    .Y(_01891_));
 sky130_fd_sc_hd__o31ai_2 _09760_ (.A1(_00585_),
    .A2(_01492_),
    .A3(_01890_),
    .B1(_01891_),
    .Y(_07385_));
 sky130_fd_sc_hd__nor3_1 _09761_ (.A(_07387_),
    .B(_07389_),
    .C(_01344_),
    .Y(_01892_));
 sky130_fd_sc_hd__o21ai_2 _09762_ (.A1(_01345_),
    .A2(_01892_),
    .B1(_01426_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_1 _09763_ (.A1(_01426_),
    .A2(_07385_),
    .B1(_01893_),
    .X(_07405_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_01633_),
    .B(_07405_),
    .Y(_01894_));
 sky130_fd_sc_hd__o31ai_1 _09765_ (.A1(_01478_),
    .A2(_01633_),
    .A3(_01889_),
    .B1(_01894_),
    .Y(_07425_));
 sky130_fd_sc_hd__nor3_1 _09766_ (.A(_07427_),
    .B(_07429_),
    .C(_01571_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _09767_ (.A(_01572_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(_07425_),
    .A1(_01896_),
    .S(net33),
    .X(_07445_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(_01888_),
    .A1(_07445_),
    .S(_01878_),
    .X(_07465_));
 sky130_fd_sc_hd__or3_1 _09770_ (.A(_01886_),
    .B(_01870_),
    .C(_07465_),
    .X(_01897_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_07469_),
    .B(_01762_),
    .Y(_01898_));
 sky130_fd_sc_hd__xor2_1 _09772_ (.A(_07467_),
    .B(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__o21ai_2 _09773_ (.A1(_01886_),
    .A2(_01870_),
    .B1(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__o21a_1 _09774_ (.A1(_07487_),
    .A2(_07486_),
    .B1(_07485_),
    .X(_01901_));
 sky130_fd_sc_hd__o21a_1 _09775_ (.A1(_07484_),
    .A2(_01901_),
    .B1(_07482_),
    .X(_01902_));
 sky130_fd_sc_hd__o21a_1 _09776_ (.A1(_07481_),
    .A2(_01902_),
    .B1(_07479_),
    .X(_01903_));
 sky130_fd_sc_hd__o21a_1 _09777_ (.A1(_01903_),
    .A2(_07478_),
    .B1(_07476_),
    .X(_01904_));
 sky130_fd_sc_hd__o21a_1 _09778_ (.A1(_07475_),
    .A2(_01904_),
    .B1(_07473_),
    .X(_01905_));
 sky130_fd_sc_hd__o21ai_2 _09779_ (.A1(_01905_),
    .A2(_07472_),
    .B1(_07490_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2b_4 _09780_ (.A(_07489_),
    .B_N(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__nor2_4 _09781_ (.A(_01786_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__a21boi_4 _09782_ (.A1(_01897_),
    .A2(_01900_),
    .B1_N(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor3_4 _09783_ (.A(_01886_),
    .B(_01870_),
    .C(_07465_),
    .Y(_01910_));
 sky130_fd_sc_hd__xnor2_2 _09784_ (.A(_07467_),
    .B(_01898_),
    .Y(_01911_));
 sky130_fd_sc_hd__a21oi_4 _09785_ (.A1(_01820_),
    .A2(_01845_),
    .B1(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__nand2b_4 _09786_ (.A_N(_07489_),
    .B(_01906_),
    .Y(_01913_));
 sky130_fd_sc_hd__buf_6 clone6 (.A(_00670_),
    .X(net6));
 sky130_fd_sc_hd__a21oi_4 _09788_ (.A1(_01913_),
    .A2(_01786_),
    .B1(_00746_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor3_4 _09789_ (.A(_01910_),
    .B(_01912_),
    .C(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_1 _09790_ (.A(_01777_),
    .B(_01854_),
    .Y(_01917_));
 sky130_fd_sc_hd__xnor2_2 _09791_ (.A(_01629_),
    .B(_01764_),
    .Y(_01918_));
 sky130_fd_sc_hd__xnor2_1 _09792_ (.A(_01797_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__o21ai_0 _09793_ (.A1(_01800_),
    .A2(_01917_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2_1 _09794_ (.A(_01755_),
    .B(_01918_),
    .Y(_01921_));
 sky130_fd_sc_hd__xnor2_1 _09795_ (.A(_00569_),
    .B(_01764_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _09796_ (.A(_07442_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__o21ai_0 _09797_ (.A1(_01921_),
    .A2(_01923_),
    .B1(_01773_),
    .Y(_01924_));
 sky130_fd_sc_hd__mux2i_1 _09798_ (.A0(_01920_),
    .A1(_01924_),
    .S(net29),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_01800_),
    .B(_01917_),
    .Y(_01926_));
 sky130_fd_sc_hd__o21ai_0 _09800_ (.A1(_01603_),
    .A2(_01755_),
    .B1(_01771_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_1 _09801_ (.A(_01777_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(_01926_),
    .A1(_01928_),
    .S(_01878_),
    .X(_01929_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(_01925_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(_01727_),
    .B(_01860_),
    .Y(_01931_));
 sky130_fd_sc_hd__a21oi_2 _09805_ (.A1(_01775_),
    .A2(_01931_),
    .B1(_01848_),
    .Y(_01932_));
 sky130_fd_sc_hd__inv_1 _09806_ (.A(_01773_),
    .Y(_01933_));
 sky130_fd_sc_hd__o21ai_0 _09807_ (.A1(_01707_),
    .A2(_01933_),
    .B1(_01775_),
    .Y(_01934_));
 sky130_fd_sc_hd__inv_1 _09808_ (.A(_01775_),
    .Y(_01935_));
 sky130_fd_sc_hd__a21oi_1 _09809_ (.A1(_01935_),
    .A2(_01801_),
    .B1(_01727_),
    .Y(_01936_));
 sky130_fd_sc_hd__a31o_1 _09810_ (.A1(_01727_),
    .A2(_01801_),
    .A3(_01934_),
    .B1(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_01811_),
    .B(_01707_),
    .Y(_01938_));
 sky130_fd_sc_hd__xnor2_1 _09812_ (.A(_01732_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__and4b_1 _09813_ (.A_N(_01930_),
    .B(_01932_),
    .C(_01937_),
    .D(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__nor3_1 _09814_ (.A(_01728_),
    .B(_01806_),
    .C(_07442_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor3_1 _09815_ (.A(_01728_),
    .B(_01732_),
    .C(_01798_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor3_1 _09816_ (.A(_01811_),
    .B(_01806_),
    .C(_01798_),
    .Y(_01943_));
 sky130_fd_sc_hd__a211oi_2 _09817_ (.A1(_01860_),
    .A2(_01941_),
    .B1(_01942_),
    .C1(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor3_4 _09818_ (.A(_01886_),
    .B(_01870_),
    .C(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_2 _09819_ (.A(_01940_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__o211ai_2 _09820_ (.A1(_01853_),
    .A2(_01856_),
    .B1(_01840_),
    .C1(_01843_),
    .Y(_01947_));
 sky130_fd_sc_hd__a2bb2oi_2 _09821_ (.A1_N(_01801_),
    .A2_N(_01776_),
    .B1(_01933_),
    .B2(net29),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_01653_),
    .B(_01728_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand3_1 _09823_ (.A(_01811_),
    .B(_01705_),
    .C(_01813_),
    .Y(_01950_));
 sky130_fd_sc_hd__o21ai_1 _09824_ (.A1(_01804_),
    .A2(_01949_),
    .B1(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__o211ai_4 _09825_ (.A1(_01653_),
    .A2(_01705_),
    .B1(_01732_),
    .C1(_01811_),
    .Y(_01952_));
 sky130_fd_sc_hd__xnor2_4 _09826_ (.A(_01816_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__a31o_1 _09827_ (.A1(_01811_),
    .A2(_01705_),
    .A3(_01813_),
    .B1(_01866_),
    .X(_01954_));
 sky130_fd_sc_hd__nor2_1 _09828_ (.A(_01811_),
    .B(_01822_),
    .Y(_01955_));
 sky130_fd_sc_hd__a211oi_2 _09829_ (.A1(_01742_),
    .A2(_01954_),
    .B1(_01955_),
    .C1(_01860_),
    .Y(_01956_));
 sky130_fd_sc_hd__a211o_1 _09830_ (.A1(_01948_),
    .A2(_01951_),
    .B1(_01953_),
    .C1(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__nor3_1 _09831_ (.A(_01948_),
    .B(_01839_),
    .C(_01951_),
    .Y(_01958_));
 sky130_fd_sc_hd__a211o_1 _09832_ (.A1(_01820_),
    .A2(_01947_),
    .B1(_01957_),
    .C1(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__nor4_4 _09833_ (.A(_01959_),
    .B(_01916_),
    .C(_01946_),
    .D(_01909_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor3b_1 _09834_ (.A(_01873_),
    .B(_01885_),
    .C_N(net428),
    .Y(_01961_));
 sky130_fd_sc_hd__o21ai_4 _09835_ (.A1(_01910_),
    .A2(_01912_),
    .B1(_01908_),
    .Y(_01962_));
 sky130_fd_sc_hd__or3_4 _09836_ (.A(_01910_),
    .B(_01912_),
    .C(_01915_),
    .X(_01963_));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(_07672_),
    .X(net414));
 sky130_fd_sc_hd__or2_0 _09838_ (.A(_01940_),
    .B(_01945_),
    .X(_01965_));
 sky130_fd_sc_hd__clkbuf_4 _09839_ (.A(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(net25),
    .B(_01870_),
    .Y(_01967_));
 sky130_fd_sc_hd__xor2_1 _09841_ (.A(_01956_),
    .B(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__a41oi_4 _09842_ (.A1(_01818_),
    .A2(_01962_),
    .A3(_01963_),
    .A4(_01966_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__a211oi_2 _09843_ (.A1(_01820_),
    .A2(_01947_),
    .B1(_01957_),
    .C1(_01958_),
    .Y(_01970_));
 sky130_fd_sc_hd__and4_2 _09844_ (.A(_01869_),
    .B(_01872_),
    .C(_01884_),
    .D(_01970_),
    .X(_01971_));
 sky130_fd_sc_hd__nand4_4 _09845_ (.A(_01962_),
    .B(_01963_),
    .C(_01966_),
    .D(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__o31ai_4 _09846_ (.A1(_01873_),
    .A2(net428),
    .A3(_01969_),
    .B1(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor3_1 _09847_ (.A(_01873_),
    .B(_01881_),
    .C(_01883_),
    .Y(_01974_));
 sky130_fd_sc_hd__and3_1 _09848_ (.A(net25),
    .B(_01840_),
    .C(_01843_),
    .X(_01975_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_01839_),
    .B(_01857_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21oi_1 _09850_ (.A1(_01975_),
    .A2(_01976_),
    .B1(_01875_),
    .Y(_01977_));
 sky130_fd_sc_hd__a21o_1 _09851_ (.A1(net428),
    .A2(_01974_),
    .B1(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__nand2b_1 _09852_ (.A_N(_01975_),
    .B(_01874_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand3_1 _09853_ (.A(_01973_),
    .B(_01978_),
    .C(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__o211ai_1 _09854_ (.A1(_01940_),
    .A2(_01945_),
    .B1(_01869_),
    .C1(_01872_),
    .Y(_01981_));
 sky130_fd_sc_hd__a31oi_1 _09855_ (.A1(_01869_),
    .A2(_01872_),
    .A3(_01884_),
    .B1(_01959_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor4b_2 _09856_ (.A(_01909_),
    .B(_01981_),
    .C(_01916_),
    .D_N(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_1 _09857_ (.A(_01679_),
    .B(_01876_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand3_1 _09858_ (.A(_01829_),
    .B(_01867_),
    .C(_01858_),
    .Y(_01985_));
 sky130_fd_sc_hd__xnor2_2 _09859_ (.A(_01984_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__xnor2_2 _09860_ (.A(_01983_),
    .B(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2b_1 _09861_ (.A(_01882_),
    .B_N(_01840_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand3_1 _09862_ (.A(_01841_),
    .B(_01825_),
    .C(_01829_),
    .Y(_01989_));
 sky130_fd_sc_hd__a311oi_2 _09863_ (.A1(_01839_),
    .A2(_01988_),
    .A3(_01857_),
    .B1(_01989_),
    .C1(_01886_),
    .Y(_01990_));
 sky130_fd_sc_hd__xnor2_1 _09864_ (.A(_01883_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__inv_1 _09865_ (.A(_01881_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand4_1 _09866_ (.A(_01869_),
    .B(_01872_),
    .C(_01992_),
    .D(_01970_),
    .Y(_01993_));
 sky130_fd_sc_hd__o32ai_1 _09867_ (.A1(_01874_),
    .A2(_01875_),
    .A3(_01883_),
    .B1(_01940_),
    .B2(_01945_),
    .Y(_01994_));
 sky130_fd_sc_hd__nor4_1 _09868_ (.A(_01909_),
    .B(_01916_),
    .C(_01993_),
    .D(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__xnor2_2 _09869_ (.A(_01991_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__or3b_1 _09870_ (.A(_01987_),
    .B(_01996_),
    .C_N(_01865_),
    .X(_01997_));
 sky130_fd_sc_hd__nor2_2 _09871_ (.A(_01980_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__o21ai_0 _09872_ (.A1(_01948_),
    .A2(_01953_),
    .B1(_01951_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _09873_ (.A(_01806_),
    .B(_01938_),
    .Y(_02000_));
 sky130_fd_sc_hd__a31oi_4 _09874_ (.A1(_01818_),
    .A2(_01845_),
    .A3(_01857_),
    .B1(_01948_),
    .Y(_02001_));
 sky130_fd_sc_hd__o211a_1 _09875_ (.A1(_01774_),
    .A2(_01801_),
    .B1(_01938_),
    .C1(_01806_),
    .X(_02002_));
 sky130_fd_sc_hd__nor4_1 _09876_ (.A(_01816_),
    .B(_02000_),
    .C(_02001_),
    .D(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__and2_0 _09877_ (.A(_01925_),
    .B(_01937_),
    .X(_02004_));
 sky130_fd_sc_hd__o211ai_4 _09878_ (.A1(_01945_),
    .A2(_02004_),
    .B1(_01929_),
    .C1(_01932_),
    .Y(_02005_));
 sky130_fd_sc_hd__a2111oi_4 _09879_ (.A1(_01966_),
    .A2(_01971_),
    .B1(_02005_),
    .C1(_01916_),
    .D1(_01909_),
    .Y(_02006_));
 sky130_fd_sc_hd__a22oi_2 _09880_ (.A1(_01967_),
    .A2(_01999_),
    .B1(_02003_),
    .B2(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(_01962_),
    .B(_01963_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor3_1 _09882_ (.A(_02008_),
    .B(_01946_),
    .C(_01971_),
    .Y(_02009_));
 sky130_fd_sc_hd__xor2_4 _09883_ (.A(_01953_),
    .B(_02001_),
    .X(_02010_));
 sky130_fd_sc_hd__or3_1 _09884_ (.A(_02000_),
    .B(_02001_),
    .C(_02002_),
    .X(_02011_));
 sky130_fd_sc_hd__o31ai_2 _09885_ (.A1(_01909_),
    .A2(_01916_),
    .A3(_02005_),
    .B1(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor4b_4 _09886_ (.A(_02007_),
    .B(_02009_),
    .C(_02010_),
    .D_N(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_8 _09887_ (.A(_01845_),
    .B(_01820_),
    .Y(_02014_));
 sky130_fd_sc_hd__inv_1 _09888_ (.A(_01937_),
    .Y(_02015_));
 sky130_fd_sc_hd__inv_1 _09889_ (.A(_01932_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand4_4 _09890_ (.A(_01869_),
    .B(_01872_),
    .C(_01884_),
    .D(_01970_),
    .Y(_02017_));
 sky130_fd_sc_hd__o211ai_1 _09891_ (.A1(_01946_),
    .A2(_02017_),
    .B1(_01962_),
    .C1(_01963_),
    .Y(_02018_));
 sky130_fd_sc_hd__or3_2 _09892_ (.A(_01930_),
    .B(_02016_),
    .C(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__nor3_1 _09893_ (.A(_07450_),
    .B(_07432_),
    .C(_01710_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _09894_ (.A(_01711_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor3_1 _09895_ (.A(_07430_),
    .B(_07412_),
    .C(_01570_),
    .Y(_02022_));
 sky130_fd_sc_hd__or2_0 _09896_ (.A(_01571_),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__nor3_1 _09897_ (.A(_07410_),
    .B(_07392_),
    .C(_01476_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor3_1 _09898_ (.A(_07390_),
    .B(_07372_),
    .C(_07371_),
    .Y(_02025_));
 sky130_fd_sc_hd__nor2_4 _09899_ (.A(_07370_),
    .B(_01492_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(_01745_),
    .B(_07388_),
    .Y(_02026_));
 sky130_fd_sc_hd__o31ai_2 _09901_ (.A1(_01344_),
    .A2(_01745_),
    .A3(_02025_),
    .B1(_02026_),
    .Y(_07408_));
 sky130_fd_sc_hd__nand2_1 _09902_ (.A(_01633_),
    .B(_07408_),
    .Y(_02027_));
 sky130_fd_sc_hd__o31ai_2 _09903_ (.A1(_01477_),
    .A2(_01633_),
    .A3(_02024_),
    .B1(_02027_),
    .Y(_07428_));
 sky130_fd_sc_hd__nor2_1 _09904_ (.A(_01733_),
    .B(_07428_),
    .Y(_02028_));
 sky130_fd_sc_hd__a21oi_1 _09905_ (.A1(net33),
    .A2(_02023_),
    .B1(_02028_),
    .Y(_07448_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(_02021_),
    .A1(_07448_),
    .S(_01878_),
    .X(_07468_));
 sky130_fd_sc_hd__nand3_2 _09907_ (.A(_01820_),
    .B(_01845_),
    .C(_07468_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor3_1 _09908_ (.A(_07470_),
    .B(_07452_),
    .C(_01761_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _09909_ (.A(_01762_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__o21ai_2 _09910_ (.A1(_01886_),
    .A2(_01870_),
    .B1(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__a21oi_1 _09911_ (.A1(_02029_),
    .A2(_02032_),
    .B1(_01603_),
    .Y(_02033_));
 sky130_fd_sc_hd__o21a_1 _09912_ (.A1(_07510_),
    .A2(_07509_),
    .B1(_07508_),
    .X(_02034_));
 sky130_fd_sc_hd__o21a_1 _09913_ (.A1(_07507_),
    .A2(_02034_),
    .B1(_07505_),
    .X(_02035_));
 sky130_fd_sc_hd__o21a_1 _09914_ (.A1(_07504_),
    .A2(_02035_),
    .B1(_07502_),
    .X(_02036_));
 sky130_fd_sc_hd__o21a_1 _09915_ (.A1(_02036_),
    .A2(_07501_),
    .B1(_07499_),
    .X(_02037_));
 sky130_fd_sc_hd__o21a_1 _09916_ (.A1(_07498_),
    .A2(_02037_),
    .B1(_07496_),
    .X(_02038_));
 sky130_fd_sc_hd__o21ai_2 _09917_ (.A1(_07495_),
    .A2(_02038_),
    .B1(_07493_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2b_1 _09918_ (.A_N(_07492_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_2 _09919_ (.A(_02040_),
    .B(_01786_),
    .Y(_02041_));
 sky130_fd_sc_hd__a21oi_4 _09920_ (.A1(_02029_),
    .A2(_02032_),
    .B1(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2b_4 _09921_ (.A(_07492_),
    .B_N(_02039_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_2 _09922_ (.A(_02043_),
    .B(_01786_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand3_1 _09923_ (.A(_02044_),
    .B(_02032_),
    .C(_02029_),
    .Y(_02045_));
 sky130_fd_sc_hd__nor3b_4 _09924_ (.A(_02042_),
    .B(_02033_),
    .C_N(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _09925_ (.A(_07472_),
    .B(_01905_),
    .Y(_02047_));
 sky130_fd_sc_hd__xnor2_2 _09926_ (.A(_07490_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__clkbuf_8 _09927_ (.A(_01603_),
    .X(_02049_));
 sky130_fd_sc_hd__nand3_1 _09928_ (.A(_02049_),
    .B(_02041_),
    .C(_02048_),
    .Y(_02050_));
 sky130_fd_sc_hd__o21ai_2 _09929_ (.A1(_02044_),
    .A2(_02048_),
    .B1(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__mux2i_4 _09930_ (.A0(_02046_),
    .A1(_02051_),
    .S(_01972_),
    .Y(_02052_));
 sky130_fd_sc_hd__a311oi_4 _09931_ (.A1(_02014_),
    .A2(_02015_),
    .A3(_02019_),
    .B1(_02006_),
    .C1(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__buf_6 _09932_ (.A(_01878_),
    .X(_02054_));
 sky130_fd_sc_hd__nor3_1 _09933_ (.A(net28),
    .B(_01800_),
    .C(_01917_),
    .Y(_02055_));
 sky130_fd_sc_hd__a21oi_1 _09934_ (.A1(net28),
    .A2(_01933_),
    .B1(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__xor2_1 _09935_ (.A(_01932_),
    .B(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__o211ai_2 _09936_ (.A1(_02008_),
    .A2(_01930_),
    .B1(_02057_),
    .C1(_02014_),
    .Y(_02058_));
 sky130_fd_sc_hd__mux2i_4 _09937_ (.A0(_01798_),
    .A1(_07442_),
    .S(net29),
    .Y(_02059_));
 sky130_fd_sc_hd__o21ai_1 _09938_ (.A1(_01886_),
    .A2(_01870_),
    .B1(_01922_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_2 _09939_ (.A(_02059_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__o2111ai_1 _09940_ (.A1(_01946_),
    .A2(_02017_),
    .B1(_02061_),
    .C1(_01963_),
    .D1(_01962_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_8 _09941_ (.A(_01870_),
    .B(_01886_),
    .Y(_02063_));
 sky130_fd_sc_hd__o21ai_1 _09942_ (.A1(net410),
    .A2(_02056_),
    .B1(_01929_),
    .Y(_02064_));
 sky130_fd_sc_hd__xor2_1 _09943_ (.A(_02062_),
    .B(_02064_),
    .X(_02065_));
 sky130_fd_sc_hd__and2_0 _09944_ (.A(_02058_),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__buf_2 _09945_ (.A(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__a2111oi_2 _09946_ (.A1(net25),
    .A2(_01845_),
    .B1(_01918_),
    .C1(_02059_),
    .D1(_00746_),
    .Y(_02068_));
 sky130_fd_sc_hd__a311o_1 _09947_ (.A1(_01603_),
    .A2(_01918_),
    .A3(_02059_),
    .B1(_01786_),
    .C1(_01913_),
    .X(_02069_));
 sky130_fd_sc_hd__a311oi_4 _09948_ (.A1(_02049_),
    .A2(net410),
    .A3(_02059_),
    .B1(_02068_),
    .C1(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_4 _09949_ (.A(_01910_),
    .B(_01912_),
    .Y(_02071_));
 sky130_fd_sc_hd__o211ai_2 _09950_ (.A1(_02049_),
    .A2(_02061_),
    .B1(_02070_),
    .C1(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__or3_1 _09951_ (.A(_01755_),
    .B(_01913_),
    .C(_07445_),
    .X(_02073_));
 sky130_fd_sc_hd__nand3_1 _09952_ (.A(_01755_),
    .B(_01913_),
    .C(_07445_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor3_1 _09953_ (.A(_01797_),
    .B(_01913_),
    .C(_01888_),
    .Y(_02075_));
 sky130_fd_sc_hd__a311oi_1 _09954_ (.A1(_01797_),
    .A2(_01913_),
    .A3(_01888_),
    .B1(_02075_),
    .C1(net28),
    .Y(_02076_));
 sky130_fd_sc_hd__a31oi_1 _09955_ (.A1(net28),
    .A2(_02073_),
    .A3(_02074_),
    .B1(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _09956_ (.A(_01907_),
    .B(_01899_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_01913_),
    .B(_01911_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _09958_ (.A(_01918_),
    .B(_02059_),
    .Y(_02080_));
 sky130_fd_sc_hd__mux2i_1 _09959_ (.A0(_02078_),
    .A1(_02079_),
    .S(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__mux2i_1 _09960_ (.A0(_02077_),
    .A1(_02081_),
    .S(_02014_),
    .Y(_02082_));
 sky130_fd_sc_hd__a2bb2oi_1 _09961_ (.A1_N(_07207_),
    .A2_N(_02082_),
    .B1(_01909_),
    .B2(_02061_),
    .Y(_02083_));
 sky130_fd_sc_hd__a2111oi_4 _09962_ (.A1(_01786_),
    .A2(_01913_),
    .B1(_01910_),
    .C1(_01912_),
    .D1(_02070_),
    .Y(_02084_));
 sky130_fd_sc_hd__a31oi_4 _09963_ (.A1(_01972_),
    .A2(_02072_),
    .A3(_02083_),
    .B1(_02084_),
    .Y(_02085_));
 sky130_fd_sc_hd__and2_0 _09964_ (.A(_01973_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__nand4_2 _09965_ (.A(_02013_),
    .B(_02053_),
    .C(_02067_),
    .D(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_2 _09966_ (.A(_01998_),
    .B(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__o21ai_2 _09967_ (.A1(_01961_),
    .A2(_02088_),
    .B1(_01986_),
    .Y(_02089_));
 sky130_fd_sc_hd__xnor2_4 _09968_ (.A(_01865_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__and3_2 _09969_ (.A(_02013_),
    .B(_02053_),
    .C(_02067_),
    .X(_02091_));
 sky130_fd_sc_hd__and3_1 _09970_ (.A(_01973_),
    .B(_01978_),
    .C(_01979_),
    .X(_02092_));
 sky130_fd_sc_hd__nor3b_2 _09971_ (.A(_01987_),
    .B(_01996_),
    .C_N(_01865_),
    .Y(_02093_));
 sky130_fd_sc_hd__and3_2 _09972_ (.A(_02092_),
    .B(_02093_),
    .C(_02085_),
    .X(_02094_));
 sky130_fd_sc_hd__nand2_2 _09973_ (.A(_02091_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor3_1 _09974_ (.A(_07453_),
    .B(_07455_),
    .C(_01760_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_4 _09975_ (.A(_07372_),
    .B(_01745_),
    .Y(_07391_));
 sky130_fd_sc_hd__nor3_1 _09976_ (.A(_07393_),
    .B(_07395_),
    .C(_07394_),
    .Y(_02097_));
 sky130_fd_sc_hd__o21ai_2 _09977_ (.A1(_01476_),
    .A2(_02097_),
    .B1(_01619_),
    .Y(_02098_));
 sky130_fd_sc_hd__o21a_1 _09978_ (.A1(_07391_),
    .A2(_01619_),
    .B1(_02098_),
    .X(_07411_));
 sky130_fd_sc_hd__nor3_1 _09979_ (.A(_07413_),
    .B(_07415_),
    .C(_01569_),
    .Y(_02099_));
 sky130_fd_sc_hd__o21ai_0 _09980_ (.A1(_01570_),
    .A2(_02099_),
    .B1(_01733_),
    .Y(_02100_));
 sky130_fd_sc_hd__o21a_1 _09981_ (.A1(_01733_),
    .A2(_07411_),
    .B1(_02100_),
    .X(_07431_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(net28),
    .B(_07431_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor3_1 _09983_ (.A(_07433_),
    .B(_07435_),
    .C(_01709_),
    .Y(_02102_));
 sky130_fd_sc_hd__or3_1 _09984_ (.A(_01710_),
    .B(_02054_),
    .C(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__nand2_1 _09985_ (.A(_02101_),
    .B(_02103_),
    .Y(_07451_));
 sky130_fd_sc_hd__nand2_1 _09986_ (.A(net410),
    .B(_07451_),
    .Y(_02104_));
 sky130_fd_sc_hd__o31ai_2 _09987_ (.A1(_01761_),
    .A2(net410),
    .A3(_02096_),
    .B1(_02104_),
    .Y(_07471_));
 sky130_fd_sc_hd__nor3_1 _09988_ (.A(_07473_),
    .B(_07475_),
    .C(_01904_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _09989_ (.A(_01905_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__mux2i_4 _09990_ (.A0(_07471_),
    .A1(_02106_),
    .S(_01972_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand4_1 _09991_ (.A(_07530_),
    .B(_07522_),
    .C(_07525_),
    .D(_07528_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand3_1 _09992_ (.A(_07513_),
    .B(_07516_),
    .C(_07519_),
    .Y(_02109_));
 sky130_fd_sc_hd__nor3_2 _09993_ (.A(_01114_),
    .B(_02108_),
    .C(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__nand3_1 _09994_ (.A(_07207_),
    .B(_02107_),
    .C(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _09995_ (.A(_01873_),
    .B(_01881_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_02112_),
    .B(net428),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _09997_ (.A(_01840_),
    .B(_01991_),
    .Y(_02114_));
 sky130_fd_sc_hd__o31a_1 _09998_ (.A1(_01885_),
    .A2(_02113_),
    .A3(_02114_),
    .B1(_01978_),
    .X(_02115_));
 sky130_fd_sc_hd__nand3_4 _09999_ (.A(_02013_),
    .B(_02067_),
    .C(_02053_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand2_1 _10000_ (.A(_02093_),
    .B(_02086_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor3_1 _10001_ (.A(_01885_),
    .B(_02113_),
    .C(_02114_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _10002_ (.A(_01979_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__o21ai_0 _10003_ (.A1(_02116_),
    .A2(_02117_),
    .B1(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__o211ai_1 _10004_ (.A1(_02095_),
    .A2(_02111_),
    .B1(_02115_),
    .C1(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__a21oi_1 _10005_ (.A1(_01818_),
    .A2(_02009_),
    .B1(_02007_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand4_2 _10006_ (.A(_01962_),
    .B(_01963_),
    .C(_01966_),
    .D(_02017_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_4 _10007_ (.A(_02123_),
    .B(_02012_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _10008_ (.A(_02010_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__and4_1 _10009_ (.A(_02125_),
    .B(_02053_),
    .C(_02067_),
    .D(_02085_),
    .X(_02126_));
 sky130_fd_sc_hd__o21ai_1 _10010_ (.A1(_01980_),
    .A2(_01997_),
    .B1(_02013_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand3_4 _10011_ (.A(_02053_),
    .B(_02067_),
    .C(_02085_),
    .Y(_02128_));
 sky130_fd_sc_hd__o22a_4 _10012_ (.A1(_02122_),
    .A2(_02126_),
    .B1(_02127_),
    .B2(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2b_1 _10013_ (.A_N(_01996_),
    .B(_02092_),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_1 _10014_ (.A(_01996_),
    .B(_02087_),
    .Y(_02131_));
 sky130_fd_sc_hd__nor2b_1 _10015_ (.A(_01987_),
    .B_N(_01865_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_2 _10016_ (.A(_01973_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__a21oi_1 _10017_ (.A1(_02130_),
    .A2(_02131_),
    .B1(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__nand3_2 _10018_ (.A(_02092_),
    .B(_02093_),
    .C(_02085_),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_8 _10019_ (.A(_02135_),
    .B(_02116_),
    .Y(_02136_));
 sky130_fd_sc_hd__buf_4 _10020_ (.A(_01786_),
    .X(_02137_));
 sky130_fd_sc_hd__nor2_1 _10021_ (.A(_07495_),
    .B(_02038_),
    .Y(_02138_));
 sky130_fd_sc_hd__xnor2_4 _10022_ (.A(_07493_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__xnor2_1 _10023_ (.A(_02137_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__o211ai_2 _10024_ (.A1(_07207_),
    .A2(_02107_),
    .B1(_02094_),
    .C1(_02091_),
    .Y(_02141_));
 sky130_fd_sc_hd__o211ai_4 _10025_ (.A1(_02136_),
    .A2(_02140_),
    .B1(_02141_),
    .C1(_02110_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand4b_2 _10026_ (.A_N(_02121_),
    .B(_02129_),
    .C(_02134_),
    .D(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__buf_4 _10027_ (.A(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__buf_6 _10028_ (.A(_01972_),
    .X(_02145_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_02072_),
    .B(_02083_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor3b_1 _10030_ (.A(net11),
    .B(_02084_),
    .C_N(_02046_),
    .Y(_02147_));
 sky130_fd_sc_hd__a31o_1 _10031_ (.A1(net11),
    .A2(_02051_),
    .A3(_02146_),
    .B1(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__xnor2_1 _10032_ (.A(_02065_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__o21ai_0 _10033_ (.A1(_02116_),
    .A2(_02135_),
    .B1(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__and2_1 _10034_ (.A(_02058_),
    .B(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__xnor2_2 _10035_ (.A(_01786_),
    .B(_01907_),
    .Y(_02152_));
 sky130_fd_sc_hd__a41oi_4 _10036_ (.A1(_01962_),
    .A2(_01963_),
    .A3(_01966_),
    .A4(_01971_),
    .B1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__xor2_4 _10037_ (.A(_02071_),
    .B(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__or3_1 _10038_ (.A(_02052_),
    .B(_02085_),
    .C(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__inv_1 _10039_ (.A(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__xnor2_1 _10040_ (.A(_02018_),
    .B(_02061_),
    .Y(_02157_));
 sky130_fd_sc_hd__o21ai_0 _10041_ (.A1(_02052_),
    .A2(_02154_),
    .B1(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__inv_1 _10042_ (.A(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _10043_ (.A(_02029_),
    .B(_02032_),
    .Y(_07488_));
 sky130_fd_sc_hd__nor2_1 _10044_ (.A(_02071_),
    .B(_07488_),
    .Y(_02160_));
 sky130_fd_sc_hd__xnor2_1 _10045_ (.A(_07207_),
    .B(_01907_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand3_1 _10046_ (.A(_01897_),
    .B(_01900_),
    .C(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__o21ai_0 _10047_ (.A1(_01910_),
    .A2(_01912_),
    .B1(_02152_),
    .Y(_02163_));
 sky130_fd_sc_hd__a21oi_1 _10048_ (.A1(_02162_),
    .A2(_02163_),
    .B1(_02048_),
    .Y(_02164_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(_02160_),
    .A1(_02164_),
    .S(_01972_),
    .X(_02165_));
 sky130_fd_sc_hd__nand4_1 _10050_ (.A(_02092_),
    .B(_02093_),
    .C(_02085_),
    .D(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__xnor2_1 _10051_ (.A(_02049_),
    .B(_02071_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _10052_ (.A(_02153_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__mux2i_4 _10053_ (.A0(_07488_),
    .A1(_02048_),
    .S(net11),
    .Y(_02169_));
 sky130_fd_sc_hd__nand3_1 _10054_ (.A(_02049_),
    .B(_02071_),
    .C(_02161_),
    .Y(_02170_));
 sky130_fd_sc_hd__or3_1 _10055_ (.A(_02049_),
    .B(_02071_),
    .C(_02152_),
    .X(_02171_));
 sky130_fd_sc_hd__a22oi_1 _10056_ (.A1(_01885_),
    .A2(_01960_),
    .B1(_02170_),
    .B2(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor4_1 _10057_ (.A(_02040_),
    .B(_02168_),
    .C(_02169_),
    .D(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__a21o_1 _10058_ (.A1(_02040_),
    .A2(_02165_),
    .B1(_02137_),
    .X(_02174_));
 sky130_fd_sc_hd__a211o_1 _10059_ (.A1(_02154_),
    .A2(_02169_),
    .B1(_07207_),
    .C1(_02040_),
    .X(_02175_));
 sky130_fd_sc_hd__o21bai_1 _10060_ (.A1(_02154_),
    .A2(_02169_),
    .B1_N(_02041_),
    .Y(_02176_));
 sky130_fd_sc_hd__o211ai_1 _10061_ (.A1(_02173_),
    .A2(_02174_),
    .B1(_02175_),
    .C1(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__o21ai_1 _10062_ (.A1(_02116_),
    .A2(_02166_),
    .B1(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__o31a_2 _10063_ (.A1(_02136_),
    .A2(_02156_),
    .A3(_02159_),
    .B1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__a31oi_2 _10064_ (.A1(_02014_),
    .A2(_02015_),
    .A3(_02019_),
    .B1(_02006_),
    .Y(_02180_));
 sky130_fd_sc_hd__a21oi_2 _10065_ (.A1(_02067_),
    .A2(_02148_),
    .B1(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__a21oi_1 _10066_ (.A1(_02122_),
    .A2(_01998_),
    .B1(_02128_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor4_2 _10067_ (.A(_02010_),
    .B(_02124_),
    .C(_02181_),
    .D(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__and3_2 _10068_ (.A(_02151_),
    .B(_02179_),
    .C(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__xnor2_2 _10069_ (.A(_01987_),
    .B(_02088_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand3_1 _10070_ (.A(_02091_),
    .B(_02094_),
    .C(_02107_),
    .Y(_02186_));
 sky130_fd_sc_hd__o211a_2 _10071_ (.A1(_02136_),
    .A2(_02139_),
    .B1(_02186_),
    .C1(_00746_),
    .X(_02187_));
 sky130_fd_sc_hd__o21a_4 _10072_ (.A1(_07530_),
    .A2(_07529_),
    .B1(_07528_),
    .X(_02188_));
 sky130_fd_sc_hd__o21a_1 _10073_ (.A1(_02188_),
    .A2(_07527_),
    .B1(_07525_),
    .X(_02189_));
 sky130_fd_sc_hd__o21a_1 _10074_ (.A1(_07524_),
    .A2(_02189_),
    .B1(_07522_),
    .X(_02190_));
 sky130_fd_sc_hd__o21a_1 _10075_ (.A1(_07521_),
    .A2(_02190_),
    .B1(_07519_),
    .X(_02191_));
 sky130_fd_sc_hd__o21a_2 _10076_ (.A1(_07518_),
    .A2(_02191_),
    .B1(_07516_),
    .X(_02192_));
 sky130_fd_sc_hd__nor2_4 _10077_ (.A(_07515_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__inv_2 _10078_ (.A(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__a21oi_4 _10079_ (.A1(_02194_),
    .A2(_07513_),
    .B1(_07512_),
    .Y(_02195_));
 sky130_fd_sc_hd__nor2_1 _10080_ (.A(_02137_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__or3_4 _10081_ (.A(_02137_),
    .B(_02195_),
    .C(_02139_),
    .X(_02197_));
 sky130_fd_sc_hd__nand3b_4 _10082_ (.A_N(_02195_),
    .B(_02139_),
    .C(_02137_),
    .Y(_02198_));
 sky130_fd_sc_hd__a22oi_4 _10083_ (.A1(_02091_),
    .A2(_02094_),
    .B1(_02198_),
    .B2(_02197_),
    .Y(_02199_));
 sky130_fd_sc_hd__or3_4 _10084_ (.A(_07207_),
    .B(_02195_),
    .C(_02107_),
    .X(_02200_));
 sky130_fd_sc_hd__nor3_4 _10085_ (.A(_02200_),
    .B(_02135_),
    .C(_02116_),
    .Y(_02201_));
 sky130_fd_sc_hd__a311o_4 _10086_ (.A1(_02136_),
    .A2(_02107_),
    .A3(_02196_),
    .B1(_02199_),
    .C1(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__nand2_1 _10087_ (.A(_01973_),
    .B(_02129_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor3_2 _10088_ (.A(_02187_),
    .B(_02202_),
    .C(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__nand4_4 _10089_ (.A(_02144_),
    .B(_02184_),
    .C(_02185_),
    .D(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__xor2_4 _10090_ (.A(_02090_),
    .B(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__nor2_8 _10091_ (.A(_02187_),
    .B(_02202_),
    .Y(_02207_));
 sky130_fd_sc_hd__and2_2 _10092_ (.A(_02151_),
    .B(_02179_),
    .X(_02208_));
 sky130_fd_sc_hd__a21o_1 _10093_ (.A1(_02067_),
    .A2(_02148_),
    .B1(_02180_),
    .X(_02209_));
 sky130_fd_sc_hd__o211ai_4 _10094_ (.A1(_01998_),
    .A2(_02128_),
    .B1(_02209_),
    .C1(_02013_),
    .Y(_02210_));
 sky130_fd_sc_hd__a211oi_4 _10095_ (.A1(_02130_),
    .A2(_02131_),
    .B1(_02210_),
    .C1(_02133_),
    .Y(_02211_));
 sky130_fd_sc_hd__inv_1 _10096_ (.A(_02115_),
    .Y(_02212_));
 sky130_fd_sc_hd__o21ai_0 _10097_ (.A1(_02116_),
    .A2(_02117_),
    .B1(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__a31oi_2 _10098_ (.A1(_02207_),
    .A2(_02208_),
    .A3(_02211_),
    .B1(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__o211ai_2 _10099_ (.A1(_02136_),
    .A2(_02139_),
    .B1(_02186_),
    .C1(_00746_),
    .Y(_02215_));
 sky130_fd_sc_hd__a311oi_4 _10100_ (.A1(_02136_),
    .A2(_02107_),
    .A3(_02196_),
    .B1(_02201_),
    .C1(_02199_),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_4 _10101_ (.A(_02216_),
    .B(_02215_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _10102_ (.A(_02151_),
    .B(_02179_),
    .Y(_02218_));
 sky130_fd_sc_hd__buf_6 _10103_ (.A(_02136_),
    .X(_02219_));
 sky130_fd_sc_hd__o211a_1 _10104_ (.A1(net16),
    .A2(_02140_),
    .B1(_02141_),
    .C1(_02110_),
    .X(_02220_));
 sky130_fd_sc_hd__o21ai_1 _10105_ (.A1(_02220_),
    .A2(_02121_),
    .B1(_02211_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor4_1 _10106_ (.A(_02217_),
    .B(_02212_),
    .C(_02218_),
    .D(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__inv_1 _10107_ (.A(_02132_),
    .Y(_02223_));
 sky130_fd_sc_hd__o21ai_1 _10108_ (.A1(_02223_),
    .A2(_02087_),
    .B1(_01996_),
    .Y(_02224_));
 sky130_fd_sc_hd__or3_1 _10109_ (.A(_02116_),
    .B(_02092_),
    .C(_02117_),
    .X(_02225_));
 sky130_fd_sc_hd__nand2_1 _10110_ (.A(_02119_),
    .B(_02212_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand3_1 _10111_ (.A(_02224_),
    .B(_02225_),
    .C(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__a31o_1 _10112_ (.A1(_02207_),
    .A2(_02208_),
    .A3(_02211_),
    .B1(_02120_),
    .X(_02228_));
 sky130_fd_sc_hd__or4b_4 _10113_ (.A(_02214_),
    .B(_02222_),
    .C(_02227_),
    .D_N(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__nand3_1 _10114_ (.A(_02095_),
    .B(_02155_),
    .C(_02158_),
    .Y(_02230_));
 sky130_fd_sc_hd__and3_1 _10115_ (.A(_02215_),
    .B(_02216_),
    .C(_02178_),
    .X(_02231_));
 sky130_fd_sc_hd__nand3_4 _10116_ (.A(_02151_),
    .B(_02179_),
    .C(_02183_),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_1 _10117_ (.A(_07207_),
    .B(_02043_),
    .Y(_02233_));
 sky130_fd_sc_hd__o21ai_1 _10118_ (.A1(_02116_),
    .A2(_02135_),
    .B1(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__xnor2_2 _10119_ (.A(_02169_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__o21ai_1 _10120_ (.A1(_02187_),
    .A2(_02202_),
    .B1(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__or3_1 _10121_ (.A(_02187_),
    .B(_02202_),
    .C(_02235_),
    .X(_02237_));
 sky130_fd_sc_hd__o211ai_4 _10122_ (.A1(_02144_),
    .A2(_02232_),
    .B1(_02236_),
    .C1(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__o211ai_4 _10123_ (.A1(_02144_),
    .A2(_02232_),
    .B1(_02207_),
    .C1(_02179_),
    .Y(_02239_));
 sky130_fd_sc_hd__and2_2 _10124_ (.A(_02095_),
    .B(_02149_),
    .X(_02240_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(_02052_),
    .B(net16),
    .Y(_02241_));
 sky130_fd_sc_hd__xor2_4 _10126_ (.A(_02154_),
    .B(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__nor2_1 _10127_ (.A(_02240_),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__o2111a_2 _10128_ (.A1(_02230_),
    .A2(_02231_),
    .B1(_02238_),
    .C1(_02239_),
    .D1(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__nand3b_4 _10129_ (.A_N(_02121_),
    .B(_02211_),
    .C(_02142_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand4_1 _10130_ (.A(_02215_),
    .B(_02216_),
    .C(_02150_),
    .D(_02179_),
    .Y(_02246_));
 sky130_fd_sc_hd__and3_1 _10131_ (.A(_02065_),
    .B(_02095_),
    .C(_02148_),
    .X(_02247_));
 sky130_fd_sc_hd__nand2_1 _10132_ (.A(_02019_),
    .B(_02058_),
    .Y(_02248_));
 sky130_fd_sc_hd__xor2_2 _10133_ (.A(_02247_),
    .B(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__a32oi_4 _10134_ (.A1(_02207_),
    .A2(_02208_),
    .A3(_02245_),
    .B1(_02246_),
    .B2(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_2 _10135_ (.A1(_02013_),
    .A2(_01998_),
    .B1(_02128_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor3_1 _10136_ (.A(_02124_),
    .B(_02181_),
    .C(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__and2_1 _10137_ (.A(_02250_),
    .B(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__o21ai_2 _10138_ (.A1(net16),
    .A2(_02139_),
    .B1(_02186_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor3_4 _10139_ (.A(_02143_),
    .B(_02217_),
    .C(_02232_),
    .Y(_02255_));
 sky130_fd_sc_hd__o21a_1 _10140_ (.A1(_07537_),
    .A2(_00584_),
    .B1(_07535_),
    .X(_02256_));
 sky130_fd_sc_hd__nor2_4 _10141_ (.A(_02256_),
    .B(_07534_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_07207_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor3_1 _10143_ (.A(_07476_),
    .B(_07478_),
    .C(_01903_),
    .Y(_02259_));
 sky130_fd_sc_hd__or2_0 _10144_ (.A(_01904_),
    .B(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__nor3_1 _10145_ (.A(_07456_),
    .B(_07458_),
    .C(_01759_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_4 _10146_ (.A(_01633_),
    .B(_07395_),
    .Y(_07414_));
 sky130_fd_sc_hd__nor3_1 _10147_ (.A(_07418_),
    .B(_07416_),
    .C(_07417_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _10148_ (.A(_01569_),
    .B(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__mux2_4 _10149_ (.A0(_07414_),
    .A1(_02263_),
    .S(_01733_),
    .X(_07434_));
 sky130_fd_sc_hd__nor3_1 _10150_ (.A(_07436_),
    .B(_07438_),
    .C(_01708_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor3_1 _10151_ (.A(_01709_),
    .B(_02054_),
    .C(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__a21o_1 _10152_ (.A1(_02054_),
    .A2(_07434_),
    .B1(_02265_),
    .X(_07454_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(_02063_),
    .B(_07454_),
    .Y(_02266_));
 sky130_fd_sc_hd__o31ai_1 _10154_ (.A1(_01760_),
    .A2(_02063_),
    .A3(_02261_),
    .B1(_02266_),
    .Y(_07474_));
 sky130_fd_sc_hd__nor2_1 _10155_ (.A(net11),
    .B(_07474_),
    .Y(_02267_));
 sky130_fd_sc_hd__a21oi_1 _10156_ (.A1(net11),
    .A2(_02260_),
    .B1(_02267_),
    .Y(_07494_));
 sky130_fd_sc_hd__nor3_1 _10157_ (.A(_07496_),
    .B(_07498_),
    .C(_02037_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _10158_ (.A(_02038_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__mux2_2 _10159_ (.A0(_07494_),
    .A1(_02269_),
    .S(_02095_),
    .X(_07511_));
 sky130_fd_sc_hd__o21ai_0 _10160_ (.A1(_00746_),
    .A2(_02258_),
    .B1(_07511_),
    .Y(_02270_));
 sky130_fd_sc_hd__or3_1 _10161_ (.A(_02137_),
    .B(_07511_),
    .C(_02257_),
    .X(_02271_));
 sky130_fd_sc_hd__and2_0 _10162_ (.A(_02270_),
    .B(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__xnor2_1 _10163_ (.A(_02137_),
    .B(_02195_),
    .Y(_02273_));
 sky130_fd_sc_hd__xor2_2 _10164_ (.A(_07513_),
    .B(_02193_),
    .X(_02274_));
 sky130_fd_sc_hd__xnor2_1 _10165_ (.A(_02137_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__o22a_1 _10166_ (.A1(_02049_),
    .A2(_02274_),
    .B1(_02275_),
    .B2(_02257_),
    .X(_02276_));
 sky130_fd_sc_hd__nor3b_2 _10167_ (.A(_02254_),
    .B(_02273_),
    .C_N(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__and3_1 _10168_ (.A(_02254_),
    .B(_02273_),
    .C(_02276_),
    .X(_02278_));
 sky130_fd_sc_hd__o32a_1 _10169_ (.A1(_02217_),
    .A2(_02144_),
    .A3(_02232_),
    .B1(_02277_),
    .B2(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__a31o_4 _10170_ (.A1(_02254_),
    .A2(_02255_),
    .A3(_02272_),
    .B1(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__and3_4 _10171_ (.A(_02244_),
    .B(_02280_),
    .C(_02253_),
    .X(_02281_));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(_02784_),
    .X(net407));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_02003_),
    .B(_02006_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(_02125_),
    .B(_02182_),
    .Y(_02284_));
 sky130_fd_sc_hd__o211ai_2 _10175_ (.A1(_02124_),
    .A2(_02128_),
    .B1(_02123_),
    .C1(_02010_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand3_4 _10176_ (.A(_02283_),
    .B(_02284_),
    .C(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__a21oi_4 _10177_ (.A1(_02017_),
    .A2(net428),
    .B1(_01969_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_2 _10178_ (.A(_02128_),
    .B(_02127_),
    .Y(_02288_));
 sky130_fd_sc_hd__xnor2_4 _10179_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__xor2_1 _10180_ (.A(_02210_),
    .B(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__and2_0 _10181_ (.A(_02286_),
    .B(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__nor2_1 _10182_ (.A(_02286_),
    .B(_02289_),
    .Y(_02292_));
 sky130_fd_sc_hd__nand4_4 _10183_ (.A(_02207_),
    .B(_02208_),
    .C(_02245_),
    .D(_02252_),
    .Y(_02293_));
 sky130_fd_sc_hd__mux2i_4 _10184_ (.A0(_02291_),
    .A1(_02292_),
    .S(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__a21oi_1 _10185_ (.A1(_01869_),
    .A2(_01872_),
    .B1(net428),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _10186_ (.A(_02295_),
    .B(_01961_),
    .Y(_02296_));
 sky130_fd_sc_hd__a21oi_1 _10187_ (.A1(_02287_),
    .A2(_02288_),
    .B1(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _10188_ (.A(_02088_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__clkinv_2 _10189_ (.A(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__nand3_2 _10190_ (.A(_02207_),
    .B(_02144_),
    .C(_02184_),
    .Y(_02300_));
 sky130_fd_sc_hd__xor2_4 _10191_ (.A(_02129_),
    .B(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__nand3_1 _10192_ (.A(_02144_),
    .B(_02184_),
    .C(_02204_),
    .Y(_02302_));
 sky130_fd_sc_hd__xor2_2 _10193_ (.A(_02185_),
    .B(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__nor4_4 _10194_ (.A(_02294_),
    .B(_02299_),
    .C(_02301_),
    .D(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__buf_4 _10195_ (.A(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__nand2_8 _10196_ (.A(_02305_),
    .B(_02281_),
    .Y(_02306_));
 sky130_fd_sc_hd__nor3_4 _10197_ (.A(_02206_),
    .B(_02306_),
    .C(_02229_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor3_1 _10198_ (.A(_07538_),
    .B(_07540_),
    .C(_00583_),
    .Y(_02308_));
 sky130_fd_sc_hd__buf_6 _10199_ (.A(_02255_),
    .X(_02309_));
 sky130_fd_sc_hd__nor3_1 _10200_ (.A(_07519_),
    .B(_07521_),
    .C(_02190_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor3_1 _10201_ (.A(_07502_),
    .B(_07504_),
    .C(_02035_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_2 _10202_ (.A(_07441_),
    .B(_02054_),
    .Y(_07460_));
 sky130_fd_sc_hd__nor3_1 _10203_ (.A(_07464_),
    .B(_07462_),
    .C(_07463_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _10204_ (.A(_01758_),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__mux2_4 _10205_ (.A0(_07460_),
    .A1(_02313_),
    .S(_02014_),
    .X(_07480_));
 sky130_fd_sc_hd__nor3_1 _10206_ (.A(_07482_),
    .B(_07484_),
    .C(_01901_),
    .Y(_02314_));
 sky130_fd_sc_hd__o21ai_0 _10207_ (.A1(_01902_),
    .A2(_02314_),
    .B1(_02145_),
    .Y(_02315_));
 sky130_fd_sc_hd__o21a_1 _10208_ (.A1(_07480_),
    .A2(_02145_),
    .B1(_02315_),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_1 _10209_ (.A(_07500_),
    .B(_02219_),
    .Y(_02316_));
 sky130_fd_sc_hd__o31ai_1 _10210_ (.A1(_02036_),
    .A2(_02219_),
    .A3(_02311_),
    .B1(_02316_),
    .Y(_07517_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(_07517_),
    .B(net8),
    .Y(_02317_));
 sky130_fd_sc_hd__o31ai_2 _10212_ (.A1(_02191_),
    .A2(net8),
    .A3(_02310_),
    .B1(_02317_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(_07536_),
    .B(net2),
    .Y(_02318_));
 sky130_fd_sc_hd__o31ai_2 _10214_ (.A1(_00584_),
    .A2(net2),
    .A3(_02308_),
    .B1(_02318_),
    .Y(_07559_));
 sky130_fd_sc_hd__o21a_1 _10215_ (.A1(_07555_),
    .A2(_07554_),
    .B1(_07553_),
    .X(_02319_));
 sky130_fd_sc_hd__o21a_1 _10216_ (.A1(_07552_),
    .A2(_02319_),
    .B1(_07573_),
    .X(_02320_));
 sky130_fd_sc_hd__o21a_1 _10217_ (.A1(_07572_),
    .A2(_02320_),
    .B1(_07570_),
    .X(_02321_));
 sky130_fd_sc_hd__o21a_1 _10218_ (.A1(_07569_),
    .A2(_02321_),
    .B1(_07567_),
    .X(_02322_));
 sky130_fd_sc_hd__o21a_1 _10219_ (.A1(_07566_),
    .A2(_02322_),
    .B1(_07564_),
    .X(_02323_));
 sky130_fd_sc_hd__o21a_1 _10220_ (.A1(_07563_),
    .A2(_02323_),
    .B1(_07561_),
    .X(_02324_));
 sky130_fd_sc_hd__nor3_1 _10221_ (.A(_07561_),
    .B(_07563_),
    .C(_02323_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _10222_ (.A(_02324_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_2 _10223_ (.A(_02228_),
    .B(_02226_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_2 _10224_ (.A(_02224_),
    .B(_02225_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _10225_ (.A(_02206_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__o31ai_1 _10226_ (.A1(_02217_),
    .A2(_02218_),
    .A3(_02221_),
    .B1(_02225_),
    .Y(_02330_));
 sky130_fd_sc_hd__a21oi_2 _10227_ (.A1(_02115_),
    .A2(_02330_),
    .B1(_02214_),
    .Y(_02331_));
 sky130_fd_sc_hd__a31oi_4 _10228_ (.A1(_02329_),
    .A2(_02281_),
    .A3(_02305_),
    .B1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__or2_2 _10229_ (.A(_02327_),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nor2_4 _10230_ (.A(_02206_),
    .B(_02229_),
    .Y(_02334_));
 sky130_fd_sc_hd__clkbuf_8 _10231_ (.A(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__nand3_4 _10232_ (.A(_02244_),
    .B(_02253_),
    .C(_02280_),
    .Y(_02336_));
 sky130_fd_sc_hd__o41ai_4 _10233_ (.A1(_02336_),
    .A2(_02294_),
    .A3(_02299_),
    .A4(_02301_),
    .B1(_02303_),
    .Y(_02337_));
 sky130_fd_sc_hd__xnor2_4 _10234_ (.A(_02090_),
    .B(_02205_),
    .Y(_02338_));
 sky130_fd_sc_hd__nand4_4 _10235_ (.A(_02207_),
    .B(_02129_),
    .C(_02144_),
    .D(_02184_),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_1 _10236_ (.A(_02133_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__xnor2_1 _10237_ (.A(_02328_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__xnor2_4 _10238_ (.A(_02289_),
    .B(_02339_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _10239_ (.A(_02299_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__and3_1 _10240_ (.A(_02338_),
    .B(_02341_),
    .C(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__o211ai_4 _10241_ (.A1(_02335_),
    .A2(_02306_),
    .B1(_02337_),
    .C1(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__nor2_4 _10242_ (.A(_02333_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__o31ai_1 _10243_ (.A1(_02217_),
    .A2(_02144_),
    .A3(_02232_),
    .B1(_02274_),
    .Y(_02347_));
 sky130_fd_sc_hd__o41a_2 _10244_ (.A1(_02217_),
    .A2(_02144_),
    .A3(_02232_),
    .A4(_07511_),
    .B1(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__xnor2_2 _10245_ (.A(_02137_),
    .B(_02257_),
    .Y(_02349_));
 sky130_fd_sc_hd__xnor2_2 _10246_ (.A(_02348_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__o211ai_4 _10247_ (.A1(_02144_),
    .A2(_02232_),
    .B1(_02235_),
    .C1(_02207_),
    .Y(_02351_));
 sky130_fd_sc_hd__xor2_1 _10248_ (.A(_02351_),
    .B(_02242_),
    .X(_02352_));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_02238_),
    .B(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_2 _10250_ (.A(_02181_),
    .B(_02251_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(_02250_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__or4_2 _10252_ (.A(_02280_),
    .B(_02350_),
    .C(_02353_),
    .D(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__nor2_1 _10253_ (.A(_02255_),
    .B(_02274_),
    .Y(_02357_));
 sky130_fd_sc_hd__a21oi_2 _10254_ (.A1(_02255_),
    .A2(_07511_),
    .B1(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand4_4 _10255_ (.A(_02334_),
    .B(_02281_),
    .C(_02304_),
    .D(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__xnor2_4 _10256_ (.A(_02240_),
    .B(_02239_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_2 _10257_ (.A(_02324_),
    .B(_07560_),
    .Y(_02361_));
 sky130_fd_sc_hd__inv_2 _10258_ (.A(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__a21oi_4 _10259_ (.A1(_02362_),
    .A2(_07558_),
    .B1(_07557_),
    .Y(_02363_));
 sky130_fd_sc_hd__inv_2 _10260_ (.A(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__xnor2_1 _10261_ (.A(_02254_),
    .B(_02273_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21oi_1 _10262_ (.A1(_02270_),
    .A2(_02271_),
    .B1(_02254_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _10263_ (.A(_02255_),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__o31ai_4 _10264_ (.A1(_02255_),
    .A2(_02276_),
    .A3(_02365_),
    .B1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__o21a_1 _10265_ (.A1(_02230_),
    .A2(_02231_),
    .B1(_02239_),
    .X(_02369_));
 sky130_fd_sc_hd__a31oi_2 _10266_ (.A1(_02238_),
    .A2(_02280_),
    .A3(_02352_),
    .B1(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__or4_4 _10267_ (.A(_02360_),
    .B(_02370_),
    .C(_02368_),
    .D(_02364_),
    .X(_02371_));
 sky130_fd_sc_hd__and2_1 _10268_ (.A(_02244_),
    .B(_02253_),
    .X(_02372_));
 sky130_fd_sc_hd__nand4b_2 _10269_ (.A_N(_02242_),
    .B(_02369_),
    .C(_02280_),
    .D(_02238_),
    .Y(_02373_));
 sky130_fd_sc_hd__a31oi_4 _10270_ (.A1(_02334_),
    .A2(_02372_),
    .A3(_02304_),
    .B1(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a211oi_4 _10271_ (.A1(_02356_),
    .A2(_02359_),
    .B1(_02374_),
    .C1(_02371_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _10272_ (.A(_02217_),
    .B(_02218_),
    .Y(_02376_));
 sky130_fd_sc_hd__a31oi_4 _10273_ (.A1(_02376_),
    .A2(_02245_),
    .A3(_02354_),
    .B1(_02251_),
    .Y(_02377_));
 sky130_fd_sc_hd__xor2_4 _10274_ (.A(_02124_),
    .B(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__a31oi_4 _10275_ (.A1(_02335_),
    .A2(_02305_),
    .A3(_02378_),
    .B1(_02336_),
    .Y(_02379_));
 sky130_fd_sc_hd__xnor2_4 _10276_ (.A(_02286_),
    .B(_02293_),
    .Y(_02380_));
 sky130_fd_sc_hd__clkbuf_4 _10277_ (.A(_02280_),
    .X(_02381_));
 sky130_fd_sc_hd__a41oi_4 _10278_ (.A1(_02244_),
    .A2(_02250_),
    .A3(_02354_),
    .A4(_02381_),
    .B1(_02378_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor3_4 _10279_ (.A(_02379_),
    .B(_02380_),
    .C(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__a211oi_4 _10280_ (.A1(_02334_),
    .A2(_02304_),
    .B1(_02380_),
    .C1(_02336_),
    .Y(_02384_));
 sky130_fd_sc_hd__xnor2_4 _10281_ (.A(_02301_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__and3_4 _10282_ (.A(_02383_),
    .B(_02385_),
    .C(_02375_),
    .X(_02386_));
 sky130_fd_sc_hd__nand2_2 _10283_ (.A(_02346_),
    .B(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(_07559_),
    .A1(_02326_),
    .S(_02387_),
    .X(_07582_));
 sky130_fd_sc_hd__or2_4 _10285_ (.A(_02333_),
    .B(_02345_),
    .X(_02388_));
 sky130_fd_sc_hd__nand3_4 _10286_ (.A(_02383_),
    .B(_02375_),
    .C(_02385_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_8 _10287_ (.A(_02389_),
    .B(_02388_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_2 _10288_ (.A(_02364_),
    .B(_02368_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_2 _10289_ (.A(_02238_),
    .B(_02381_),
    .Y(_02392_));
 sky130_fd_sc_hd__o31ai_2 _10290_ (.A1(_02381_),
    .A2(_02350_),
    .A3(_02392_),
    .B1(_02359_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand3_1 _10291_ (.A(_02376_),
    .B(_02245_),
    .C(_02354_),
    .Y(_02394_));
 sky130_fd_sc_hd__o21ai_1 _10292_ (.A1(_02376_),
    .A2(_02354_),
    .B1(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_02244_),
    .B(_02381_),
    .Y(_02396_));
 sky130_fd_sc_hd__xor2_1 _10294_ (.A(_02250_),
    .B(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__xnor2_2 _10295_ (.A(_02351_),
    .B(_02242_),
    .Y(_02398_));
 sky130_fd_sc_hd__a21oi_1 _10296_ (.A1(_02238_),
    .A2(_02381_),
    .B1(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__and3_1 _10297_ (.A(_02238_),
    .B(_02280_),
    .C(_02398_),
    .X(_02400_));
 sky130_fd_sc_hd__o21ai_1 _10298_ (.A1(_02399_),
    .A2(_02400_),
    .B1(_02369_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand3_4 _10299_ (.A(_02335_),
    .B(_02281_),
    .C(_02305_),
    .Y(_02402_));
 sky130_fd_sc_hd__o31ai_1 _10300_ (.A1(_02395_),
    .A2(_02397_),
    .A3(_02401_),
    .B1(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__and4b_1 _10301_ (.A_N(_02360_),
    .B(_02393_),
    .C(_02383_),
    .D(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__nand4_4 _10302_ (.A(_02391_),
    .B(_02343_),
    .C(_02385_),
    .D(_02404_),
    .Y(_02405_));
 sky130_fd_sc_hd__nor2b_2 _10303_ (.A(_02301_),
    .B_N(_02384_),
    .Y(_02406_));
 sky130_fd_sc_hd__xor2_2 _10304_ (.A(_02342_),
    .B(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__a21oi_4 _10305_ (.A1(_02375_),
    .A2(_02383_),
    .B1(_02385_),
    .Y(_02408_));
 sky130_fd_sc_hd__a211oi_4 _10306_ (.A1(_02388_),
    .A2(_02386_),
    .B1(_02407_),
    .C1(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__inv_1 _10307_ (.A(_02300_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2b_1 _10308_ (.A(_02289_),
    .B_N(_02129_),
    .Y(_02411_));
 sky130_fd_sc_hd__o21ai_1 _10309_ (.A1(_02410_),
    .A2(_02384_),
    .B1(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__xnor2_2 _10310_ (.A(_02299_),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__o31ai_4 _10311_ (.A1(_02342_),
    .A2(_02346_),
    .A3(_02389_),
    .B1(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__o211ai_4 _10312_ (.A1(_02390_),
    .A2(_02405_),
    .B1(_02409_),
    .C1(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__or3_1 _10313_ (.A(_02379_),
    .B(_02380_),
    .C(_02382_),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_1 _10314_ (.A(_02402_),
    .B(_02397_),
    .Y(_02417_));
 sky130_fd_sc_hd__or3_1 _10315_ (.A(_02381_),
    .B(_02350_),
    .C(_02353_),
    .X(_02418_));
 sky130_fd_sc_hd__a21oi_2 _10316_ (.A1(_02418_),
    .A2(_02359_),
    .B1(_02371_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand3_1 _10317_ (.A(_02244_),
    .B(_02250_),
    .C(_02381_),
    .Y(_02420_));
 sky130_fd_sc_hd__a31oi_1 _10318_ (.A1(_02335_),
    .A2(_02281_),
    .A3(_02305_),
    .B1(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__xnor2_1 _10319_ (.A(_02395_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21oi_2 _10320_ (.A1(_02417_),
    .A2(_02419_),
    .B1(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__o32ai_4 _10321_ (.A1(_02375_),
    .A2(_02416_),
    .A3(_02423_),
    .B1(_02389_),
    .B2(_02388_),
    .Y(_02424_));
 sky130_fd_sc_hd__clkinvlp_4 _10322_ (.A(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__o21ai_4 _10323_ (.A1(_02335_),
    .A2(_02306_),
    .B1(_02337_),
    .Y(_02426_));
 sky130_fd_sc_hd__or3_2 _10324_ (.A(_02206_),
    .B(_02426_),
    .C(_02333_),
    .X(_02427_));
 sky130_fd_sc_hd__o32ai_4 _10325_ (.A1(_02206_),
    .A2(_02335_),
    .A3(_02306_),
    .B1(_02339_),
    .B2(_02133_),
    .Y(_02428_));
 sky130_fd_sc_hd__xor2_4 _10326_ (.A(_02328_),
    .B(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__o21a_1 _10327_ (.A1(net13),
    .A2(_02405_),
    .B1(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__nor4_4 _10328_ (.A(_02415_),
    .B(_02425_),
    .C(_02427_),
    .D(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__and2_1 _10329_ (.A(_02402_),
    .B(_02401_),
    .X(_02432_));
 sky130_fd_sc_hd__and2_0 _10330_ (.A(_02402_),
    .B(_02397_),
    .X(_02433_));
 sky130_fd_sc_hd__a31o_1 _10331_ (.A1(_02335_),
    .A2(_02372_),
    .A3(_02305_),
    .B1(_02373_),
    .X(_02434_));
 sky130_fd_sc_hd__nand3_1 _10332_ (.A(_02402_),
    .B(_02397_),
    .C(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__mux2i_2 _10333_ (.A0(_02433_),
    .A1(_02435_),
    .S(_02419_),
    .Y(_02436_));
 sky130_fd_sc_hd__a21oi_4 _10334_ (.A1(_02346_),
    .A2(_02386_),
    .B1(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor3_4 _10335_ (.A(_02360_),
    .B(_02432_),
    .C(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__o21ai_2 _10336_ (.A1(_02381_),
    .A2(_02350_),
    .B1(_02359_),
    .Y(_02439_));
 sky130_fd_sc_hd__and3_2 _10337_ (.A(_02392_),
    .B(_02391_),
    .C(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__nand3_1 _10338_ (.A(_02335_),
    .B(_02372_),
    .C(_02305_),
    .Y(_02441_));
 sky130_fd_sc_hd__and3_2 _10339_ (.A(_02238_),
    .B(_02381_),
    .C(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__a211oi_4 _10340_ (.A1(_02391_),
    .A2(_02439_),
    .B1(_02442_),
    .C1(_02392_),
    .Y(_02443_));
 sky130_fd_sc_hd__o21a_1 _10341_ (.A1(_07575_),
    .A2(_07574_),
    .B1(_07581_),
    .X(_02444_));
 sky130_fd_sc_hd__o21a_1 _10342_ (.A1(_07580_),
    .A2(_02444_),
    .B1(_07578_),
    .X(_02445_));
 sky130_fd_sc_hd__o21a_1 _10343_ (.A1(_07577_),
    .A2(_02445_),
    .B1(_07596_),
    .X(_02446_));
 sky130_fd_sc_hd__o21a_1 _10344_ (.A1(_07595_),
    .A2(_02446_),
    .B1(_07593_),
    .X(_02447_));
 sky130_fd_sc_hd__o21a_1 _10345_ (.A1(_07592_),
    .A2(_02447_),
    .B1(_07590_),
    .X(_02448_));
 sky130_fd_sc_hd__o21a_1 _10346_ (.A1(_07589_),
    .A2(_02448_),
    .B1(_07587_),
    .X(_02449_));
 sky130_fd_sc_hd__or2_4 _10347_ (.A(_07586_),
    .B(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__a21oi_4 _10348_ (.A1(_02450_),
    .A2(_07584_),
    .B1(_07583_),
    .Y(_02451_));
 sky130_fd_sc_hd__nor3_1 _10349_ (.A(_07516_),
    .B(_07518_),
    .C(_02191_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor3_1 _10350_ (.A(_07499_),
    .B(_07501_),
    .C(_02036_),
    .Y(_02453_));
 sky130_fd_sc_hd__nor3_1 _10351_ (.A(_07479_),
    .B(_07481_),
    .C(_01902_),
    .Y(_02454_));
 sky130_fd_sc_hd__or2_0 _10352_ (.A(_01903_),
    .B(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__nor3_1 _10353_ (.A(_07459_),
    .B(_07461_),
    .C(_01758_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor3_1 _10354_ (.A(_07441_),
    .B(_07439_),
    .C(_07440_),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _10355_ (.A(_01708_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__a21oi_4 _10356_ (.A1(_01730_),
    .A2(_01658_),
    .B1(_07418_),
    .Y(_07437_));
 sky130_fd_sc_hd__mux2_4 _10357_ (.A0(_02458_),
    .A1(_07437_),
    .S(_02054_),
    .X(_07457_));
 sky130_fd_sc_hd__nand2_1 _10358_ (.A(_02063_),
    .B(_07457_),
    .Y(_02459_));
 sky130_fd_sc_hd__o31ai_1 _10359_ (.A1(_01759_),
    .A2(_02063_),
    .A3(_02456_),
    .B1(_02459_),
    .Y(_07477_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_02145_),
    .B(_07477_),
    .Y(_02460_));
 sky130_fd_sc_hd__a21oi_1 _10361_ (.A1(_02145_),
    .A2(_02455_),
    .B1(_02460_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(net16),
    .B(_07497_),
    .Y(_02461_));
 sky130_fd_sc_hd__o31ai_2 _10363_ (.A1(_02037_),
    .A2(net16),
    .A3(_02453_),
    .B1(_02461_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand2_1 _10364_ (.A(net8),
    .B(_07514_),
    .Y(_02462_));
 sky130_fd_sc_hd__o31ai_4 _10365_ (.A1(_02192_),
    .A2(_02255_),
    .A3(_02452_),
    .B1(_02462_),
    .Y(_07533_));
 sky130_fd_sc_hd__nor2_1 _10366_ (.A(_02348_),
    .B(_07533_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor3_1 _10367_ (.A(_07535_),
    .B(_07537_),
    .C(_00584_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _10368_ (.A(_02256_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__nor2_1 _10369_ (.A(_02350_),
    .B(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__mux2_1 _10370_ (.A0(_02463_),
    .A1(_02466_),
    .S(_02402_),
    .X(_02467_));
 sky130_fd_sc_hd__nand2_2 _10371_ (.A(_02467_),
    .B(_02451_),
    .Y(_02468_));
 sky130_fd_sc_hd__a21oi_1 _10372_ (.A1(_02381_),
    .A2(_02441_),
    .B1(_02368_),
    .Y(_02469_));
 sky130_fd_sc_hd__xor2_1 _10373_ (.A(_07558_),
    .B(_02361_),
    .X(_02470_));
 sky130_fd_sc_hd__nand2_1 _10374_ (.A(_02451_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__inv_1 _10375_ (.A(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__a31oi_4 _10376_ (.A1(_02335_),
    .A2(_02281_),
    .A3(_02305_),
    .B1(_02349_),
    .Y(_02473_));
 sky130_fd_sc_hd__xnor3_1 _10377_ (.A(_02348_),
    .B(_02363_),
    .C(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__nand3_1 _10378_ (.A(_02469_),
    .B(_02472_),
    .C(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__o31ai_4 _10379_ (.A1(_02468_),
    .A2(_02389_),
    .A3(_02388_),
    .B1(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__o31a_4 _10380_ (.A1(_02390_),
    .A2(_02440_),
    .A3(_02443_),
    .B1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__a21boi_4 _10381_ (.A1(_02431_),
    .A2(_02438_),
    .B1_N(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_2 _10382_ (.A(_02370_),
    .B(_02374_),
    .Y(_02479_));
 sky130_fd_sc_hd__or3_2 _10383_ (.A(net13),
    .B(_02440_),
    .C(_02443_),
    .X(_02480_));
 sky130_fd_sc_hd__or2_0 _10384_ (.A(_02480_),
    .B(_02476_),
    .X(_02481_));
 sky130_fd_sc_hd__o21bai_4 _10385_ (.A1(_02398_),
    .A2(_02442_),
    .B1_N(_02400_),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _10386_ (.A(_02391_),
    .B(_02439_),
    .Y(_02483_));
 sky130_fd_sc_hd__nor3_4 _10387_ (.A(_02392_),
    .B(_02390_),
    .C(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__xor2_4 _10388_ (.A(_02482_),
    .B(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__nand3_2 _10389_ (.A(_02479_),
    .B(_02481_),
    .C(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__o21a_1 _10390_ (.A1(_07607_),
    .A2(_07606_),
    .B1(_07605_),
    .X(_02487_));
 sky130_fd_sc_hd__o21a_1 _10391_ (.A1(_07604_),
    .A2(_02487_),
    .B1(_07602_),
    .X(_02488_));
 sky130_fd_sc_hd__o21a_1 _10392_ (.A1(_07601_),
    .A2(_02488_),
    .B1(_07599_),
    .X(_02489_));
 sky130_fd_sc_hd__o21a_1 _10393_ (.A1(_07598_),
    .A2(_02489_),
    .B1(_07619_),
    .X(_02490_));
 sky130_fd_sc_hd__o21a_1 _10394_ (.A1(_07618_),
    .A2(_02490_),
    .B1(_07616_),
    .X(_02491_));
 sky130_fd_sc_hd__o21ai_2 _10395_ (.A1(_07615_),
    .A2(_02491_),
    .B1(_07613_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand2b_1 _10396_ (.A_N(_07612_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__a21oi_2 _10397_ (.A1(_02493_),
    .A2(_07610_),
    .B1(_07609_),
    .Y(_02494_));
 sky130_fd_sc_hd__and4b_2 _10398_ (.A_N(_07582_),
    .B(_02438_),
    .C(_02494_),
    .D(_02477_),
    .X(_02495_));
 sky130_fd_sc_hd__xnor2_2 _10399_ (.A(_02348_),
    .B(_02473_),
    .Y(_02496_));
 sky130_fd_sc_hd__xnor2_1 _10400_ (.A(_02363_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__nor2_1 _10401_ (.A(_02451_),
    .B(_02470_),
    .Y(_02498_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(_07533_),
    .A1(_02465_),
    .S(_02402_),
    .X(_07556_));
 sky130_fd_sc_hd__xnor2_1 _10403_ (.A(_02451_),
    .B(_07556_),
    .Y(_02499_));
 sky130_fd_sc_hd__nand2_1 _10404_ (.A(_02496_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__o32a_1 _10405_ (.A1(_02472_),
    .A2(_02497_),
    .A3(_02498_),
    .B1(_02500_),
    .B2(_02387_),
    .X(_02501_));
 sky130_fd_sc_hd__xor2_1 _10406_ (.A(_07584_),
    .B(_02450_),
    .X(_02502_));
 sky130_fd_sc_hd__a21o_1 _10407_ (.A1(_07610_),
    .A2(_02493_),
    .B1(_07609_),
    .X(_02503_));
 sky130_fd_sc_hd__nor3_2 _10408_ (.A(_02501_),
    .B(_02502_),
    .C(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__a21oi_4 _10409_ (.A1(_02495_),
    .A2(_02431_),
    .B1(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21oi_1 _10410_ (.A1(_02363_),
    .A2(_02496_),
    .B1(_02469_),
    .Y(_02506_));
 sky130_fd_sc_hd__a21oi_1 _10411_ (.A1(_02346_),
    .A2(_02386_),
    .B1(_02483_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _10412_ (.A(_02472_),
    .B(_02474_),
    .Y(_02508_));
 sky130_fd_sc_hd__o221ai_2 _10413_ (.A1(_02387_),
    .A2(_02468_),
    .B1(_02506_),
    .B2(_02507_),
    .C1(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__and3_1 _10414_ (.A(_02480_),
    .B(_02438_),
    .C(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__and2b_1 _10415_ (.A_N(_02476_),
    .B(_02509_),
    .X(_02511_));
 sky130_fd_sc_hd__a21oi_2 _10416_ (.A1(_02431_),
    .A2(_02510_),
    .B1(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__or4_1 _10417_ (.A(_02478_),
    .B(_02486_),
    .C(_02505_),
    .D(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__buf_6 _10418_ (.A(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__nor2_1 _10419_ (.A(_02379_),
    .B(_02382_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand2_1 _10420_ (.A(_02346_),
    .B(_02385_),
    .Y(_02516_));
 sky130_fd_sc_hd__and2_0 _10421_ (.A(_02375_),
    .B(_02515_),
    .X(_02517_));
 sky130_fd_sc_hd__o21ai_1 _10422_ (.A1(_02380_),
    .A2(_02516_),
    .B1(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__o21a_1 _10423_ (.A1(net3),
    .A2(_02515_),
    .B1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__buf_6 _10424_ (.A(_02390_),
    .X(_02520_));
 sky130_fd_sc_hd__o211a_1 _10425_ (.A1(_02520_),
    .A2(_02405_),
    .B1(_02409_),
    .C1(_02414_),
    .X(_02521_));
 sky130_fd_sc_hd__nand2b_1 _10426_ (.A_N(_02426_),
    .B(_02338_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor2_1 _10427_ (.A(_02333_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__o21ai_4 _10428_ (.A1(_02390_),
    .A2(_02405_),
    .B1(_02429_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand4_4 _10429_ (.A(_02521_),
    .B(_02424_),
    .C(_02523_),
    .D(_02524_),
    .Y(_02525_));
 sky130_fd_sc_hd__nor2_1 _10430_ (.A(_02360_),
    .B(_02432_),
    .Y(_02526_));
 sky130_fd_sc_hd__o311a_1 _10431_ (.A1(_02520_),
    .A2(_02440_),
    .A3(_02443_),
    .B1(_02476_),
    .C1(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__nand2_1 _10432_ (.A(_02525_),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__buf_6 _10433_ (.A(_02387_),
    .X(_02529_));
 sky130_fd_sc_hd__a21o_2 _10434_ (.A1(net3),
    .A2(net12),
    .B1(_02423_),
    .X(_02530_));
 sky130_fd_sc_hd__nand2b_1 _10435_ (.A_N(_02360_),
    .B(_02374_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _10436_ (.A(_02391_),
    .B(_02393_),
    .Y(_02532_));
 sky130_fd_sc_hd__o211ai_2 _10437_ (.A1(_02432_),
    .A2(_02532_),
    .B1(_02360_),
    .C1(_02434_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _10438_ (.A(_02419_),
    .B(_02387_),
    .Y(_02534_));
 sky130_fd_sc_hd__nand2_1 _10439_ (.A(_02402_),
    .B(_02401_),
    .Y(_02535_));
 sky130_fd_sc_hd__a32oi_4 _10440_ (.A1(_02531_),
    .A2(_02533_),
    .A3(_02534_),
    .B1(_02477_),
    .B2(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor3_1 _10441_ (.A(_02437_),
    .B(_02530_),
    .C(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand3_2 _10442_ (.A(_02519_),
    .B(_02528_),
    .C(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_2 _10443_ (.A(_02514_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__clkbuf_4 _10444_ (.A(_02431_),
    .X(_02540_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(net3),
    .B(_02423_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21o_1 _10446_ (.A1(_02515_),
    .A2(_02541_),
    .B1(_02520_),
    .X(_02542_));
 sky130_fd_sc_hd__nand3_1 _10447_ (.A(_02438_),
    .B(_02477_),
    .C(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__a21oi_1 _10448_ (.A1(_02516_),
    .A2(_02517_),
    .B1(_02379_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _10449_ (.A(_02379_),
    .B(_02517_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_02380_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__o21a_1 _10451_ (.A1(_02380_),
    .A2(_02544_),
    .B1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__o21ai_2 _10452_ (.A1(_02540_),
    .A2(_02543_),
    .B1(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_8 _10453_ (.A(_02438_),
    .B(_02477_),
    .Y(_02549_));
 sky130_fd_sc_hd__or4b_2 _10454_ (.A(_02431_),
    .B(_02549_),
    .C(_02547_),
    .D_N(_02542_),
    .X(_02550_));
 sky130_fd_sc_hd__o21ai_4 _10455_ (.A1(net23),
    .A2(_02405_),
    .B1(_02414_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2b_1 _10456_ (.A(_02437_),
    .B_N(_02424_),
    .Y(_02552_));
 sky130_fd_sc_hd__o211ai_2 _10457_ (.A1(_02427_),
    .A2(_02430_),
    .B1(_02527_),
    .C1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _10458_ (.A(net23),
    .B(_02405_),
    .Y(_02554_));
 sky130_fd_sc_hd__xnor2_1 _10459_ (.A(_02426_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__o311ai_4 _10460_ (.A1(net13),
    .A2(_02440_),
    .A3(_02443_),
    .B1(_02476_),
    .C1(_02526_),
    .Y(_02556_));
 sky130_fd_sc_hd__o31ai_2 _10461_ (.A1(_02425_),
    .A2(_02437_),
    .A3(_02556_),
    .B1(_02551_),
    .Y(_02557_));
 sky130_fd_sc_hd__o2111ai_2 _10462_ (.A1(_02551_),
    .A2(_02553_),
    .B1(_02555_),
    .C1(_02409_),
    .D1(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__a21o_2 _10463_ (.A1(_02548_),
    .A2(_02550_),
    .B1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__nor3_1 _10464_ (.A(_02425_),
    .B(_02437_),
    .C(_02556_),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _10465_ (.A(_02335_),
    .B(_02306_),
    .Y(_02561_));
 sky130_fd_sc_hd__a21oi_1 _10466_ (.A1(_02281_),
    .A2(_02305_),
    .B1(_02338_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21oi_2 _10467_ (.A1(_02338_),
    .A2(_02561_),
    .B1(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor3_1 _10468_ (.A(_02426_),
    .B(net13),
    .C(_02405_),
    .Y(_02564_));
 sky130_fd_sc_hd__xnor2_1 _10469_ (.A(_02563_),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_2 _10470_ (.A(_02327_),
    .B(_02332_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor4_1 _10471_ (.A(_02360_),
    .B(_02379_),
    .C(_02380_),
    .D(_02382_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand4_1 _10472_ (.A(_07555_),
    .B(_07558_),
    .C(_07561_),
    .D(_07567_),
    .Y(_02568_));
 sky130_fd_sc_hd__nand4_1 _10473_ (.A(_07553_),
    .B(_07564_),
    .C(_07570_),
    .D(_07573_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor4_1 _10474_ (.A(_01114_),
    .B(_02368_),
    .C(_02568_),
    .D(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand4_2 _10475_ (.A(_02393_),
    .B(_02403_),
    .C(_02567_),
    .D(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__a211oi_4 _10476_ (.A1(_02566_),
    .A2(_02571_),
    .B1(_02389_),
    .C1(_02345_),
    .Y(_02572_));
 sky130_fd_sc_hd__o31a_1 _10477_ (.A1(_02522_),
    .A2(net23),
    .A3(_02405_),
    .B1(_02429_),
    .X(_02573_));
 sky130_fd_sc_hd__nor2_4 _10478_ (.A(_02572_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__a311oi_4 _10479_ (.A1(_02338_),
    .A2(_02566_),
    .A3(_02524_),
    .B1(_02415_),
    .C1(_02426_),
    .Y(_02575_));
 sky130_fd_sc_hd__and3_1 _10480_ (.A(_02565_),
    .B(_02574_),
    .C(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__nor2_1 _10481_ (.A(_02214_),
    .B(_02222_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand4_2 _10482_ (.A(_02577_),
    .B(_02329_),
    .C(_02281_),
    .D(_02305_),
    .Y(_02578_));
 sky130_fd_sc_hd__inv_1 _10483_ (.A(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__a21oi_2 _10484_ (.A1(_02327_),
    .A2(_02579_),
    .B1(_02332_),
    .Y(_02580_));
 sky130_fd_sc_hd__xor2_4 _10485_ (.A(_02572_),
    .B(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__o311ai_4 _10486_ (.A1(_02332_),
    .A2(_02345_),
    .A3(_02389_),
    .B1(_02578_),
    .C1(_02327_),
    .Y(_02582_));
 sky130_fd_sc_hd__and2_0 _10487_ (.A(_02581_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__xor2_1 _10488_ (.A(_02563_),
    .B(_02564_),
    .X(_02584_));
 sky130_fd_sc_hd__and3_1 _10489_ (.A(_02584_),
    .B(_02574_),
    .C(_02583_),
    .X(_02585_));
 sky130_fd_sc_hd__a31oi_2 _10490_ (.A1(_02560_),
    .A2(_02576_),
    .A3(_02583_),
    .B1(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand4_1 _10491_ (.A(_02521_),
    .B(_02523_),
    .C(_02524_),
    .D(_02552_),
    .Y(_02587_));
 sky130_fd_sc_hd__a21o_2 _10492_ (.A1(_02527_),
    .A2(_02587_),
    .B1(_02536_),
    .X(_02588_));
 sky130_fd_sc_hd__o32ai_2 _10493_ (.A1(_07582_),
    .A2(_02525_),
    .A3(_02549_),
    .B1(_02501_),
    .B2(_02502_),
    .Y(_02589_));
 sky130_fd_sc_hd__a21o_1 _10494_ (.A1(_02540_),
    .A2(_02510_),
    .B1(_02511_),
    .X(_02590_));
 sky130_fd_sc_hd__nand4_1 _10495_ (.A(_07599_),
    .B(_07607_),
    .C(_07610_),
    .D(_07602_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand4_1 _10496_ (.A(_07605_),
    .B(_07613_),
    .C(_07616_),
    .D(_07619_),
    .Y(_02592_));
 sky130_fd_sc_hd__nor3_2 _10497_ (.A(_01114_),
    .B(_02591_),
    .C(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__and4b_1 _10498_ (.A_N(_02588_),
    .B(_02589_),
    .C(_02590_),
    .D(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__nor3_2 _10499_ (.A(_02559_),
    .B(_02586_),
    .C(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__clkbuf_4 _10500_ (.A(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_4 _10501_ (.A(_02539_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__or3_1 _10502_ (.A(_07613_),
    .B(_07615_),
    .C(_02491_),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_1 _10503_ (.A(_02492_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__nor2_8 _10504_ (.A(_02549_),
    .B(_02525_),
    .Y(_02600_));
 sky130_fd_sc_hd__nor3_1 _10505_ (.A(_07590_),
    .B(_07592_),
    .C(_02447_),
    .Y(_02601_));
 sky130_fd_sc_hd__nor3_1 _10506_ (.A(_07567_),
    .B(_07569_),
    .C(_02321_),
    .Y(_02602_));
 sky130_fd_sc_hd__or2_0 _10507_ (.A(_02322_),
    .B(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__nor3_1 _10508_ (.A(_07544_),
    .B(_07546_),
    .C(_00581_),
    .Y(_02604_));
 sky130_fd_sc_hd__nor3_1 _10509_ (.A(_07525_),
    .B(_07527_),
    .C(_02188_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor3_1 _10510_ (.A(_07510_),
    .B(_07508_),
    .C(_07509_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21oi_2 _10511_ (.A1(_01885_),
    .A2(_01960_),
    .B1(_07487_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(_02219_),
    .B(_07506_),
    .Y(_02607_));
 sky130_fd_sc_hd__o31ai_4 _10513_ (.A1(_02034_),
    .A2(_02219_),
    .A3(_02606_),
    .B1(_02607_),
    .Y(_07523_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(_02309_),
    .B(_07523_),
    .Y(_02608_));
 sky130_fd_sc_hd__o31ai_2 _10515_ (.A1(_02189_),
    .A2(_02309_),
    .A3(_02605_),
    .B1(_02608_),
    .Y(_07542_));
 sky130_fd_sc_hd__nand2_1 _10516_ (.A(_02307_),
    .B(_07542_),
    .Y(_02609_));
 sky130_fd_sc_hd__o31ai_2 _10517_ (.A1(_00582_),
    .A2(_02307_),
    .A3(_02604_),
    .B1(_02609_),
    .Y(_07565_));
 sky130_fd_sc_hd__nor2_1 _10518_ (.A(net12),
    .B(_07565_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21oi_1 _10519_ (.A1(net12),
    .A2(_02603_),
    .B1(_02610_),
    .Y(_07588_));
 sky130_fd_sc_hd__buf_6 _10520_ (.A(_02600_),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _10521_ (.A(_07588_),
    .B(net19),
    .Y(_02612_));
 sky130_fd_sc_hd__o31ai_1 _10522_ (.A1(_02448_),
    .A2(_02600_),
    .A3(_02601_),
    .B1(_02612_),
    .Y(_07611_));
 sky130_fd_sc_hd__nor2_1 _10523_ (.A(_07611_),
    .B(_02597_),
    .Y(_02613_));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(_02597_),
    .A2(_02599_),
    .B1(_02613_),
    .Y(_07640_));
 sky130_fd_sc_hd__inv_1 _10525_ (.A(\butterfly_count[1] ),
    .Y(_07666_));
 sky130_fd_sc_hd__inv_2 _10526_ (.A(\butterfly_count[0] ),
    .Y(_07716_));
 sky130_fd_sc_hd__o21a_1 _10527_ (.A1(_07621_),
    .A2(_07620_),
    .B1(_07627_),
    .X(_02614_));
 sky130_fd_sc_hd__o21a_1 _10528_ (.A1(_07626_),
    .A2(_02614_),
    .B1(_07624_),
    .X(_02615_));
 sky130_fd_sc_hd__o21a_1 _10529_ (.A1(_07623_),
    .A2(_02615_),
    .B1(_07633_),
    .X(_02616_));
 sky130_fd_sc_hd__o21a_1 _10530_ (.A1(_07632_),
    .A2(_02616_),
    .B1(_07630_),
    .X(_02617_));
 sky130_fd_sc_hd__o21a_1 _10531_ (.A1(_02617_),
    .A2(_07629_),
    .B1(_07639_),
    .X(_02618_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(_07638_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__xnor2_1 _10533_ (.A(_07636_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__or2_4 _10534_ (.A(_02514_),
    .B(_02538_),
    .X(_02621_));
 sky130_fd_sc_hd__nand4b_1 _10535_ (.A_N(_02588_),
    .B(_02589_),
    .C(_02590_),
    .D(_02593_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand2b_2 _10536_ (.A_N(_02586_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__nor3_4 _10537_ (.A(_02623_),
    .B(_02559_),
    .C(_02621_),
    .Y(_02624_));
 sky130_fd_sc_hd__nor3_1 _10538_ (.A(_07616_),
    .B(_07618_),
    .C(_02490_),
    .Y(_02625_));
 sky130_fd_sc_hd__buf_6 _10539_ (.A(_02624_),
    .X(_02626_));
 sky130_fd_sc_hd__nor3_1 _10540_ (.A(_07593_),
    .B(_07595_),
    .C(_02446_),
    .Y(_02627_));
 sky130_fd_sc_hd__nor3_1 _10541_ (.A(_07570_),
    .B(_07572_),
    .C(_02320_),
    .Y(_02628_));
 sky130_fd_sc_hd__or2_0 _10542_ (.A(_02321_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__nor3_1 _10543_ (.A(_07547_),
    .B(_07549_),
    .C(_00580_),
    .Y(_02630_));
 sky130_fd_sc_hd__nor3_1 _10544_ (.A(_07530_),
    .B(_07528_),
    .C(_07529_),
    .Y(_02631_));
 sky130_fd_sc_hd__nor2_4 _10545_ (.A(_07510_),
    .B(_02219_),
    .Y(_07526_));
 sky130_fd_sc_hd__nand2_1 _10546_ (.A(_02309_),
    .B(_07526_),
    .Y(_02632_));
 sky130_fd_sc_hd__o31ai_4 _10547_ (.A1(_02188_),
    .A2(_02309_),
    .A3(_02631_),
    .B1(_02632_),
    .Y(_07545_));
 sky130_fd_sc_hd__nand2_1 _10548_ (.A(_02307_),
    .B(_07545_),
    .Y(_02633_));
 sky130_fd_sc_hd__o31ai_2 _10549_ (.A1(_00581_),
    .A2(_02307_),
    .A3(_02630_),
    .B1(_02633_),
    .Y(_07568_));
 sky130_fd_sc_hd__nor2_1 _10550_ (.A(_02529_),
    .B(_07568_),
    .Y(_02634_));
 sky130_fd_sc_hd__a21oi_1 _10551_ (.A1(_02529_),
    .A2(_02629_),
    .B1(_02634_),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(net19),
    .B(_07591_),
    .Y(_02635_));
 sky130_fd_sc_hd__o31ai_1 _10553_ (.A1(_02447_),
    .A2(net19),
    .A3(_02627_),
    .B1(_02635_),
    .Y(_07614_));
 sky130_fd_sc_hd__nand2_1 _10554_ (.A(net7),
    .B(_07614_),
    .Y(_02636_));
 sky130_fd_sc_hd__o31ai_1 _10555_ (.A1(_02491_),
    .A2(_02624_),
    .A3(_02625_),
    .B1(_02636_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_02437_),
    .B(_02556_),
    .Y(_02637_));
 sky130_fd_sc_hd__o21ai_4 _10557_ (.A1(_02540_),
    .A2(_02549_),
    .B1(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__xnor2_1 _10558_ (.A(_02514_),
    .B(_02588_),
    .Y(_02639_));
 sky130_fd_sc_hd__nor2_1 _10559_ (.A(_02638_),
    .B(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(_02528_),
    .B(_02537_),
    .Y(_02641_));
 sky130_fd_sc_hd__nor3_1 _10561_ (.A(_02540_),
    .B(_02549_),
    .C(_02530_),
    .Y(_02642_));
 sky130_fd_sc_hd__xnor2_1 _10562_ (.A(_02519_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__o21ai_1 _10563_ (.A1(_02514_),
    .A2(_02641_),
    .B1(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__o21a_1 _10564_ (.A1(_02478_),
    .A2(_02484_),
    .B1(_02482_),
    .X(_02645_));
 sky130_fd_sc_hd__o21ai_1 _10565_ (.A1(_02478_),
    .A2(_02484_),
    .B1(_02535_),
    .Y(_02646_));
 sky130_fd_sc_hd__o21ai_4 _10566_ (.A1(_02479_),
    .A2(_02645_),
    .B1(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__nor2_1 _10567_ (.A(_02540_),
    .B(_02549_),
    .Y(_02648_));
 sky130_fd_sc_hd__xor2_1 _10568_ (.A(_02530_),
    .B(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__a211oi_1 _10569_ (.A1(_02548_),
    .A2(_02550_),
    .B1(_02647_),
    .C1(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__o211a_1 _10570_ (.A1(_02624_),
    .A2(_02640_),
    .B1(_02644_),
    .C1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__o21ai_0 _10571_ (.A1(_02505_),
    .A2(_02512_),
    .B1(_02485_),
    .Y(_02652_));
 sky130_fd_sc_hd__nor3_2 _10572_ (.A(net23),
    .B(_02440_),
    .C(_02443_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand2_1 _10573_ (.A(_02653_),
    .B(_02485_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21o_1 _10574_ (.A1(_02540_),
    .A2(_02495_),
    .B1(_02504_),
    .X(_02655_));
 sky130_fd_sc_hd__a21oi_1 _10575_ (.A1(_02655_),
    .A2(_02590_),
    .B1(_02481_),
    .Y(_02656_));
 sky130_fd_sc_hd__a211oi_1 _10576_ (.A1(_02652_),
    .A2(_02654_),
    .B1(_02478_),
    .C1(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__a21oi_1 _10577_ (.A1(_02539_),
    .A2(_02596_),
    .B1(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__a21o_1 _10578_ (.A1(_07584_),
    .A2(_02450_),
    .B1(_07583_),
    .X(_02659_));
 sky130_fd_sc_hd__nand3_1 _10579_ (.A(_02346_),
    .B(_02386_),
    .C(_07556_),
    .Y(_02660_));
 sky130_fd_sc_hd__o21ai_0 _10580_ (.A1(net23),
    .A2(_02470_),
    .B1(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__or2_1 _10581_ (.A(_02659_),
    .B(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_02659_),
    .B(_02661_),
    .Y(_02663_));
 sky130_fd_sc_hd__o21ai_2 _10583_ (.A1(_02600_),
    .A2(_02662_),
    .B1(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__and2_0 _10584_ (.A(_02438_),
    .B(_02477_),
    .X(_02665_));
 sky130_fd_sc_hd__nand3_1 _10585_ (.A(_07582_),
    .B(_02540_),
    .C(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__o21ai_0 _10586_ (.A1(_02525_),
    .A2(_02549_),
    .B1(_02502_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand3_1 _10587_ (.A(_02494_),
    .B(_02666_),
    .C(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__nor3_1 _10588_ (.A(_02655_),
    .B(_02664_),
    .C(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a21oi_1 _10589_ (.A1(_02540_),
    .A2(_02665_),
    .B1(_02662_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand3_1 _10590_ (.A(_02363_),
    .B(net12),
    .C(_02496_),
    .Y(_02671_));
 sky130_fd_sc_hd__o21ai_1 _10591_ (.A1(_02363_),
    .A2(_02496_),
    .B1(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__xnor2_1 _10592_ (.A(_02670_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__and2_0 _10593_ (.A(_02505_),
    .B(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__a211o_2 _10594_ (.A1(_02539_),
    .A2(_02595_),
    .B1(_02669_),
    .C1(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__nor3_1 _10595_ (.A(_07587_),
    .B(_07589_),
    .C(_02448_),
    .Y(_02676_));
 sky130_fd_sc_hd__o21ai_0 _10596_ (.A1(_02449_),
    .A2(_02676_),
    .B1(_02662_),
    .Y(_02677_));
 sky130_fd_sc_hd__nor3_1 _10597_ (.A(_07541_),
    .B(_07543_),
    .C(_00582_),
    .Y(_02678_));
 sky130_fd_sc_hd__nor3_1 _10598_ (.A(_07522_),
    .B(_07524_),
    .C(_02189_),
    .Y(_02679_));
 sky130_fd_sc_hd__nor2_1 _10599_ (.A(_07464_),
    .B(_02063_),
    .Y(_07483_));
 sky130_fd_sc_hd__nor3_1 _10600_ (.A(_07487_),
    .B(_07485_),
    .C(_07486_),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_1 _10601_ (.A(_01901_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__mux2_4 _10602_ (.A0(_07483_),
    .A1(_02681_),
    .S(_02145_),
    .X(_07503_));
 sky130_fd_sc_hd__nor3_1 _10603_ (.A(_07505_),
    .B(_07507_),
    .C(_02034_),
    .Y(_02682_));
 sky130_fd_sc_hd__o21ai_0 _10604_ (.A1(_02035_),
    .A2(_02682_),
    .B1(_02095_),
    .Y(_02683_));
 sky130_fd_sc_hd__o21a_1 _10605_ (.A1(_02095_),
    .A2(_07503_),
    .B1(_02683_),
    .X(_07520_));
 sky130_fd_sc_hd__nand2_1 _10606_ (.A(net8),
    .B(_07520_),
    .Y(_02684_));
 sky130_fd_sc_hd__o31ai_2 _10607_ (.A1(_02190_),
    .A2(net8),
    .A3(_02679_),
    .B1(_02684_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_1 _10608_ (.A(net2),
    .B(_07539_),
    .Y(_02685_));
 sky130_fd_sc_hd__o31ai_2 _10609_ (.A1(_00583_),
    .A2(net2),
    .A3(_02678_),
    .B1(_02685_),
    .Y(_07562_));
 sky130_fd_sc_hd__nor3_1 _10610_ (.A(_07564_),
    .B(_07566_),
    .C(_02322_),
    .Y(_02686_));
 sky130_fd_sc_hd__nor2_1 _10611_ (.A(_02323_),
    .B(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__mux2i_1 _10612_ (.A0(_07562_),
    .A1(_02687_),
    .S(net12),
    .Y(_02688_));
 sky130_fd_sc_hd__nand2_1 _10613_ (.A(_02600_),
    .B(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__o21ai_1 _10614_ (.A1(_02618_),
    .A2(_07638_),
    .B1(_07636_),
    .Y(_02690_));
 sky130_fd_sc_hd__nand2b_1 _10615_ (.A_N(_07635_),
    .B(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21oi_4 _10616_ (.A1(_02691_),
    .A2(_07642_),
    .B1(_07641_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _10617_ (.A(_02692_),
    .B(_02663_),
    .Y(_02693_));
 sky130_fd_sc_hd__a21oi_2 _10618_ (.A1(_02677_),
    .A2(_02689_),
    .B1(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__xor2_1 _10619_ (.A(_07610_),
    .B(_02493_),
    .X(_02695_));
 sky130_fd_sc_hd__nand2b_1 _10620_ (.A_N(_02695_),
    .B(_02692_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2_1 _10621_ (.A(_02664_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__nand2_1 _10622_ (.A(_02666_),
    .B(_02667_),
    .Y(_02698_));
 sky130_fd_sc_hd__xnor2_1 _10623_ (.A(_02494_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__a32o_2 _10624_ (.A1(_02539_),
    .A2(_02694_),
    .A3(_02595_),
    .B1(_02697_),
    .B2(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__and4bb_4 _10625_ (.A_N(_02512_),
    .B_N(_02658_),
    .C(_02700_),
    .D(_02675_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2_8 _10626_ (.A(_02701_),
    .B(_02651_),
    .Y(_02702_));
 sky130_fd_sc_hd__o21ai_2 _10627_ (.A1(net3),
    .A2(_02515_),
    .B1(_02518_),
    .Y(_02703_));
 sky130_fd_sc_hd__nor2_1 _10628_ (.A(_02703_),
    .B(_02584_),
    .Y(_02704_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(_02703_),
    .A1(_02704_),
    .S(_02642_),
    .X(_02705_));
 sky130_fd_sc_hd__nor4_2 _10630_ (.A(_02514_),
    .B(_02641_),
    .C(_02559_),
    .D(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__nor2_1 _10631_ (.A(_02565_),
    .B(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nor4_4 _10632_ (.A(_02478_),
    .B(_02486_),
    .C(_02505_),
    .D(_02512_),
    .Y(_02708_));
 sky130_fd_sc_hd__and4_1 _10633_ (.A(_02519_),
    .B(_02528_),
    .C(_02537_),
    .D(_02547_),
    .X(_02709_));
 sky130_fd_sc_hd__nand3_1 _10634_ (.A(_02521_),
    .B(_02708_),
    .C(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2_1 _10635_ (.A(_02415_),
    .B(_02553_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_1 _10636_ (.A(_02575_),
    .B(_02560_),
    .Y(_02712_));
 sky130_fd_sc_hd__o21ai_2 _10637_ (.A1(_02555_),
    .A2(_02711_),
    .B1(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__nand2_1 _10638_ (.A(_02710_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21ai_2 _10639_ (.A1(_02624_),
    .A2(_02707_),
    .B1(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__inv_1 _10640_ (.A(_02581_),
    .Y(_02716_));
 sky130_fd_sc_hd__nor3_1 _10641_ (.A(_02530_),
    .B(_02588_),
    .C(_02638_),
    .Y(_02717_));
 sky130_fd_sc_hd__a21oi_1 _10642_ (.A1(_02548_),
    .A2(_02550_),
    .B1(_02558_),
    .Y(_02718_));
 sky130_fd_sc_hd__nor2_1 _10643_ (.A(_02703_),
    .B(_02565_),
    .Y(_02719_));
 sky130_fd_sc_hd__and3_1 _10644_ (.A(_02584_),
    .B(_02575_),
    .C(_02560_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_2 _10645_ (.A(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__a41oi_1 _10646_ (.A1(_02708_),
    .A2(_02717_),
    .A3(_02718_),
    .A4(_02719_),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__xor2_1 _10647_ (.A(_02574_),
    .B(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__o21a_1 _10648_ (.A1(_02716_),
    .A2(_02723_),
    .B1(_02597_),
    .X(_02724_));
 sky130_fd_sc_hd__nand2_2 _10649_ (.A(_02708_),
    .B(_02709_),
    .Y(_02725_));
 sky130_fd_sc_hd__nor3_1 _10650_ (.A(_02415_),
    .B(_02596_),
    .C(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand4_2 _10651_ (.A(_02708_),
    .B(_02717_),
    .C(_02718_),
    .D(_02719_),
    .Y(_02727_));
 sky130_fd_sc_hd__nor4_1 _10652_ (.A(_02514_),
    .B(_02538_),
    .C(_02586_),
    .D(_02594_),
    .Y(_02728_));
 sky130_fd_sc_hd__o21ai_1 _10653_ (.A1(_02574_),
    .A2(_02721_),
    .B1(_02581_),
    .Y(_02729_));
 sky130_fd_sc_hd__a31oi_2 _10654_ (.A1(_02574_),
    .A2(_02581_),
    .A3(_02721_),
    .B1(_02582_),
    .Y(_02730_));
 sky130_fd_sc_hd__o31ai_4 _10655_ (.A1(_02727_),
    .A2(_02728_),
    .A3(_02729_),
    .B1(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__nor2_1 _10656_ (.A(_02346_),
    .B(_02389_),
    .Y(_02732_));
 sky130_fd_sc_hd__nor2_1 _10657_ (.A(_02732_),
    .B(_02408_),
    .Y(_02733_));
 sky130_fd_sc_hd__nor3_2 _10658_ (.A(_02425_),
    .B(_02540_),
    .C(_02549_),
    .Y(_02734_));
 sky130_fd_sc_hd__xnor2_2 _10659_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor2_1 _10660_ (.A(_02406_),
    .B(_02732_),
    .Y(_02736_));
 sky130_fd_sc_hd__xnor2_1 _10661_ (.A(_02342_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__a211o_1 _10662_ (.A1(_02708_),
    .A2(_02709_),
    .B1(_02735_),
    .C1(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__xor2_1 _10663_ (.A(_02342_),
    .B(_02736_),
    .X(_02739_));
 sky130_fd_sc_hd__nand4b_2 _10664_ (.A_N(_02733_),
    .B(_02708_),
    .C(_02739_),
    .D(_02709_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand3b_4 _10665_ (.A_N(_02596_),
    .B(_02738_),
    .C(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__or3_1 _10666_ (.A(_02732_),
    .B(_02407_),
    .C(_02408_),
    .X(_02742_));
 sky130_fd_sc_hd__o21ai_0 _10667_ (.A1(_02427_),
    .A2(_02430_),
    .B1(_02552_),
    .Y(_02743_));
 sky130_fd_sc_hd__o31ai_2 _10668_ (.A1(_02415_),
    .A2(_02556_),
    .A3(_02743_),
    .B1(_02557_),
    .Y(_02744_));
 sky130_fd_sc_hd__a22oi_2 _10669_ (.A1(_02551_),
    .A2(_02742_),
    .B1(_02725_),
    .B2(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand4b_1 _10670_ (.A_N(_02726_),
    .B(_02731_),
    .C(_02741_),
    .D(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__or3_1 _10671_ (.A(_02715_),
    .B(_02724_),
    .C(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_4 _10672_ (.A(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__nor2_8 _10673_ (.A(_02748_),
    .B(_02702_),
    .Y(_02749_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(_02620_),
    .A1(_07634_),
    .S(_02749_),
    .X(_07660_));
 sky130_fd_sc_hd__o21ai_2 _10675_ (.A1(_02702_),
    .A2(_02748_),
    .B1(net396),
    .Y(_02750_));
 sky130_fd_sc_hd__maj3_1 _10676_ (.A(_02503_),
    .B(_02698_),
    .C(_02696_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_02664_),
    .B(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__o21ai_1 _10678_ (.A1(_02664_),
    .A2(_02668_),
    .B1(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _10679_ (.A(_02655_),
    .B(_02590_),
    .Y(_02754_));
 sky130_fd_sc_hd__a221o_1 _10680_ (.A1(_02655_),
    .A2(_02597_),
    .B1(_02673_),
    .B2(_02700_),
    .C1(_02590_),
    .X(_02755_));
 sky130_fd_sc_hd__o21ai_2 _10681_ (.A1(_02754_),
    .A2(net1),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21oi_1 _10682_ (.A1(_02597_),
    .A2(_02753_),
    .B1(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand4_1 _10683_ (.A(_02485_),
    .B(_02675_),
    .C(_02750_),
    .D(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand3_1 _10684_ (.A(_02540_),
    .B(_02480_),
    .C(_02438_),
    .Y(_02759_));
 sky130_fd_sc_hd__and2_0 _10685_ (.A(_02590_),
    .B(_02675_),
    .X(_02760_));
 sky130_fd_sc_hd__nor2_1 _10686_ (.A(_02754_),
    .B(net1),
    .Y(_02761_));
 sky130_fd_sc_hd__a221o_1 _10687_ (.A1(_02476_),
    .A2(_02759_),
    .B1(_02700_),
    .B2(_02760_),
    .C1(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__nand2_1 _10688_ (.A(_02759_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__xnor2_1 _10689_ (.A(_02653_),
    .B(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__nor2_1 _10690_ (.A(_02449_),
    .B(_02676_),
    .Y(_02765_));
 sky130_fd_sc_hd__o21a_1 _10691_ (.A1(net19),
    .A2(_02765_),
    .B1(_02689_),
    .X(_07608_));
 sky130_fd_sc_hd__mux2i_4 _10692_ (.A0(_02695_),
    .A1(_07608_),
    .S(_02624_),
    .Y(_02766_));
 sky130_fd_sc_hd__xnor2_1 _10693_ (.A(_02692_),
    .B(_02766_),
    .Y(_02767_));
 sky130_fd_sc_hd__xnor2_1 _10694_ (.A(_07642_),
    .B(_02691_),
    .Y(_02768_));
 sky130_fd_sc_hd__inv_1 _10695_ (.A(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__o32a_1 _10696_ (.A1(_07640_),
    .A2(_02702_),
    .A3(_02748_),
    .B1(_02767_),
    .B2(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__nor2_1 _10697_ (.A(net1),
    .B(_02668_),
    .Y(_02771_));
 sky130_fd_sc_hd__a21oi_2 _10698_ (.A1(_02503_),
    .A2(_02698_),
    .B1(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__o21a_1 _10699_ (.A1(_07647_),
    .A2(_07646_),
    .B1(_07645_),
    .X(_02773_));
 sky130_fd_sc_hd__o21a_1 _10700_ (.A1(_07644_),
    .A2(_02773_),
    .B1(_07659_),
    .X(_02774_));
 sky130_fd_sc_hd__o21a_1 _10701_ (.A1(_07658_),
    .A2(_02774_),
    .B1(_07656_),
    .X(_02775_));
 sky130_fd_sc_hd__o21a_1 _10702_ (.A1(_07655_),
    .A2(_02775_),
    .B1(_07653_),
    .X(_02776_));
 sky130_fd_sc_hd__o21a_1 _10703_ (.A1(_02776_),
    .A2(_07652_),
    .B1(_07650_),
    .X(_02777_));
 sky130_fd_sc_hd__nor2_2 _10704_ (.A(_07649_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nor2b_1 _10705_ (.A(_02778_),
    .B_N(_07665_),
    .Y(_02779_));
 sky130_fd_sc_hd__nor2_2 _10706_ (.A(_02779_),
    .B(_07664_),
    .Y(_02780_));
 sky130_fd_sc_hd__clkinv_2 _10707_ (.A(_02780_),
    .Y(_02781_));
 sky130_fd_sc_hd__a21oi_4 _10708_ (.A1(_02781_),
    .A2(_07662_),
    .B1(_07661_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_2 _10709_ (.A(_02772_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__nor2_4 _10710_ (.A(_02783_),
    .B(_02770_),
    .Y(_02784_));
 sky130_fd_sc_hd__nor3b_4 _10711_ (.A(_02758_),
    .B(_02764_),
    .C_N(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__nor3_1 _10712_ (.A(_02514_),
    .B(_02588_),
    .C(net1),
    .Y(_02786_));
 sky130_fd_sc_hd__a21oi_1 _10713_ (.A1(_02514_),
    .A2(_02588_),
    .B1(_02786_),
    .Y(_02787_));
 sky130_fd_sc_hd__inv_1 _10714_ (.A(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__xnor2_2 _10715_ (.A(_02482_),
    .B(_02484_),
    .Y(_02789_));
 sky130_fd_sc_hd__a2111oi_4 _10716_ (.A1(_02539_),
    .A2(_02596_),
    .B1(_02653_),
    .C1(_02789_),
    .D1(_02754_),
    .Y(_02790_));
 sky130_fd_sc_hd__xnor2_4 _10717_ (.A(_02647_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__o21ai_2 _10718_ (.A1(_02702_),
    .A2(_02748_),
    .B1(net390),
    .Y(_02792_));
 sky130_fd_sc_hd__xor2_4 _10719_ (.A(_02791_),
    .B(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__o21ai_1 _10720_ (.A1(_02621_),
    .A2(_02596_),
    .B1(_02644_),
    .Y(_02794_));
 sky130_fd_sc_hd__and2_0 _10721_ (.A(_02651_),
    .B(_02701_),
    .X(_02795_));
 sky130_fd_sc_hd__clkbuf_4 _10722_ (.A(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__nor3_1 _10723_ (.A(_02715_),
    .B(_02724_),
    .C(_02746_),
    .Y(_02797_));
 sky130_fd_sc_hd__xnor2_2 _10724_ (.A(_02530_),
    .B(_02648_),
    .Y(_02798_));
 sky130_fd_sc_hd__o21ai_1 _10725_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02597_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand4_1 _10726_ (.A(_02798_),
    .B(_02799_),
    .C(_02701_),
    .D(_02791_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21oi_1 _10727_ (.A1(_02796_),
    .A2(_02797_),
    .B1(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__xor2_1 _10728_ (.A(_02794_),
    .B(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__nand2_1 _10729_ (.A(_02708_),
    .B(_02597_),
    .Y(_02803_));
 sky130_fd_sc_hd__nor3_1 _10730_ (.A(_02588_),
    .B(_02638_),
    .C(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__xnor2_1 _10731_ (.A(_02649_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2b_1 _10732_ (.A_N(_02638_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__nor4_1 _10733_ (.A(_02788_),
    .B(_02793_),
    .C(_02802_),
    .D(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__nor2_1 _10734_ (.A(_02596_),
    .B(_02725_),
    .Y(_02808_));
 sky130_fd_sc_hd__xnor2_1 _10735_ (.A(_02735_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__and3_1 _10736_ (.A(_02796_),
    .B(_02809_),
    .C(_02747_),
    .X(_02810_));
 sky130_fd_sc_hd__o21bai_2 _10737_ (.A1(_02796_),
    .A2(_02809_),
    .B1_N(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__and4b_1 _10738_ (.A_N(_02794_),
    .B(_02791_),
    .C(_02798_),
    .D(_02799_),
    .X(_02812_));
 sky130_fd_sc_hd__o211ai_1 _10739_ (.A1(_02702_),
    .A2(_02748_),
    .B1(_02812_),
    .C1(net390),
    .Y(_02813_));
 sky130_fd_sc_hd__a31o_1 _10740_ (.A1(_02621_),
    .A2(_02548_),
    .A3(_02550_),
    .B1(_02808_),
    .X(_02814_));
 sky130_fd_sc_hd__xor2_1 _10741_ (.A(_02813_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__nor2b_1 _10742_ (.A(_02811_),
    .B_N(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__nand2_1 _10743_ (.A(_02733_),
    .B(_02734_),
    .Y(_02817_));
 sky130_fd_sc_hd__xnor2_1 _10744_ (.A(_02739_),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__o31ai_1 _10745_ (.A1(_02742_),
    .A2(net1),
    .A3(_02725_),
    .B1(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__or2_0 _10746_ (.A(_02596_),
    .B(_02725_),
    .X(_02820_));
 sky130_fd_sc_hd__nor3_1 _10747_ (.A(_02409_),
    .B(_02596_),
    .C(_02725_),
    .Y(_02821_));
 sky130_fd_sc_hd__a41oi_1 _10748_ (.A1(_02796_),
    .A2(_02820_),
    .A3(_02748_),
    .A4(_02819_),
    .B1(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__o22a_2 _10749_ (.A1(_02810_),
    .A2(_02819_),
    .B1(_02822_),
    .B2(_02735_),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_1 _10750_ (.A(_02738_),
    .B(_02740_),
    .Y(_02824_));
 sky130_fd_sc_hd__nor2_1 _10751_ (.A(_02596_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__a22o_1 _10752_ (.A1(_02551_),
    .A2(_02742_),
    .B1(_02725_),
    .B2(_02744_),
    .X(_02826_));
 sky130_fd_sc_hd__nor2_1 _10753_ (.A(_02826_),
    .B(_02726_),
    .Y(_02827_));
 sky130_fd_sc_hd__a22oi_4 _10754_ (.A1(_02710_),
    .A2(_02713_),
    .B1(_02706_),
    .B2(_02623_),
    .Y(_02828_));
 sky130_fd_sc_hd__o211ai_1 _10755_ (.A1(_02702_),
    .A2(_02825_),
    .B1(_02827_),
    .C1(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__o21ai_2 _10756_ (.A1(_02415_),
    .A2(_02820_),
    .B1(_02745_),
    .Y(_02830_));
 sky130_fd_sc_hd__inv_1 _10757_ (.A(_02731_),
    .Y(_02831_));
 sky130_fd_sc_hd__o21ai_0 _10758_ (.A1(_02826_),
    .A2(_02726_),
    .B1(_02828_),
    .Y(_02832_));
 sky130_fd_sc_hd__o41ai_1 _10759_ (.A1(_02830_),
    .A2(_02715_),
    .A3(_02724_),
    .A4(_02831_),
    .B1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand3_1 _10760_ (.A(_02796_),
    .B(_02741_),
    .C(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__and3_1 _10761_ (.A(_02708_),
    .B(_02717_),
    .C(_02719_),
    .X(_02835_));
 sky130_fd_sc_hd__a21oi_1 _10762_ (.A1(_02575_),
    .A2(_02560_),
    .B1(_02584_),
    .Y(_02836_));
 sky130_fd_sc_hd__nor2_1 _10763_ (.A(_02836_),
    .B(_02721_),
    .Y(_02837_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(_02706_),
    .B(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__a31oi_2 _10765_ (.A1(_02623_),
    .A2(_02706_),
    .A3(_02835_),
    .B1(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__inv_1 _10766_ (.A(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__nor3_2 _10767_ (.A(_02825_),
    .B(_02830_),
    .C(_02715_),
    .Y(_02841_));
 sky130_fd_sc_hd__nand2_1 _10768_ (.A(_02597_),
    .B(_02723_),
    .Y(_02842_));
 sky130_fd_sc_hd__a31oi_2 _10769_ (.A1(_02796_),
    .A2(_02748_),
    .A3(_02841_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__and4_1 _10770_ (.A(_02796_),
    .B(_02842_),
    .C(_02748_),
    .D(_02841_),
    .X(_02844_));
 sky130_fd_sc_hd__a2111oi_1 _10771_ (.A1(_02829_),
    .A2(_02834_),
    .B1(_02840_),
    .C1(_02843_),
    .D1(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__inv_1 _10772_ (.A(_02724_),
    .Y(_02846_));
 sky130_fd_sc_hd__and3_1 _10773_ (.A(_02795_),
    .B(_02747_),
    .C(_02841_),
    .X(_02847_));
 sky130_fd_sc_hd__inv_1 _10774_ (.A(_02727_),
    .Y(_02848_));
 sky130_fd_sc_hd__nor3_1 _10775_ (.A(_02581_),
    .B(_02721_),
    .C(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__inv_1 _10776_ (.A(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__a31oi_2 _10777_ (.A1(_02795_),
    .A2(_02747_),
    .A3(_02841_),
    .B1(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__o31ai_1 _10778_ (.A1(_02478_),
    .A2(_02486_),
    .A3(_02622_),
    .B1(_02582_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_1 _10779_ (.A1(_02848_),
    .A2(_02852_),
    .B1(_02721_),
    .X(_02853_));
 sky130_fd_sc_hd__nand3_1 _10780_ (.A(_02574_),
    .B(_02581_),
    .C(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__o21ai_2 _10781_ (.A1(_02574_),
    .A2(_02581_),
    .B1(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__nor2_1 _10782_ (.A(_02715_),
    .B(_02724_),
    .Y(_02856_));
 sky130_fd_sc_hd__a41oi_4 _10783_ (.A1(_02796_),
    .A2(_02741_),
    .A3(_02827_),
    .A4(_02856_),
    .B1(_02731_),
    .Y(_02857_));
 sky130_fd_sc_hd__a2111oi_4 _10784_ (.A1(_02846_),
    .A2(_02847_),
    .B1(_02851_),
    .C1(_02855_),
    .D1(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__and3b_1 _10785_ (.A_N(_02823_),
    .B(_02845_),
    .C(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__and4_1 _10786_ (.A(_02785_),
    .B(_02807_),
    .C(_02816_),
    .D(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__buf_6 _10787_ (.A(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__inv_8 _10788_ (.A(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__buf_8 _10789_ (.A(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__buf_8 _10790_ (.A(_02863_),
    .X(_00553_));
 sky130_fd_sc_hd__nor3_1 _10791_ (.A(_07650_),
    .B(_07652_),
    .C(_02776_),
    .Y(_02864_));
 sky130_fd_sc_hd__or2_0 _10792_ (.A(_02777_),
    .B(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__buf_6 _10793_ (.A(_02749_),
    .X(_02866_));
 sky130_fd_sc_hd__nor3_1 _10794_ (.A(_07630_),
    .B(_07632_),
    .C(_02616_),
    .Y(_02867_));
 sky130_fd_sc_hd__nor3_1 _10795_ (.A(_07599_),
    .B(_07601_),
    .C(_02488_),
    .Y(_02868_));
 sky130_fd_sc_hd__nor3_1 _10796_ (.A(_07578_),
    .B(_07580_),
    .C(_02444_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor3_1 _10797_ (.A(_07553_),
    .B(_07555_),
    .C(_07554_),
    .Y(_02870_));
 sky130_fd_sc_hd__or3_4 _10798_ (.A(_02520_),
    .B(_02319_),
    .C(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__o31ai_4 _10799_ (.A1(_07532_),
    .A2(net2),
    .A3(_02529_),
    .B1(_02871_),
    .Y(_07576_));
 sky130_fd_sc_hd__nand2_1 _10800_ (.A(_02611_),
    .B(_07576_),
    .Y(_02872_));
 sky130_fd_sc_hd__o31ai_1 _10801_ (.A1(_02445_),
    .A2(_02611_),
    .A3(_02869_),
    .B1(_02872_),
    .Y(_07597_));
 sky130_fd_sc_hd__nand2_1 _10802_ (.A(net7),
    .B(_07597_),
    .Y(_02873_));
 sky130_fd_sc_hd__o31ai_1 _10803_ (.A1(_02489_),
    .A2(net7),
    .A3(_02868_),
    .B1(_02873_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_1 _10804_ (.A(net18),
    .B(_07628_),
    .Y(_02874_));
 sky130_fd_sc_hd__o31ai_1 _10805_ (.A1(_02617_),
    .A2(net18),
    .A3(_02867_),
    .B1(_02874_),
    .Y(_07648_));
 sky130_fd_sc_hd__nor2_1 _10806_ (.A(_07648_),
    .B(net434),
    .Y(_02875_));
 sky130_fd_sc_hd__a21oi_1 _10807_ (.A1(net434),
    .A2(_02865_),
    .B1(_02875_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(_02597_),
    .B(_02753_),
    .Y(_02876_));
 sky130_fd_sc_hd__inv_1 _10809_ (.A(_02750_),
    .Y(_02877_));
 sky130_fd_sc_hd__a31oi_2 _10810_ (.A1(net393),
    .A2(_02876_),
    .A3(net38),
    .B1(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__xnor2_2 _10811_ (.A(_02675_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__or3b_1 _10812_ (.A(_02758_),
    .B(_02764_),
    .C_N(net407),
    .X(_02880_));
 sky130_fd_sc_hd__buf_4 _10813_ (.A(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__or2_0 _10814_ (.A(_02788_),
    .B(_02793_),
    .X(_02882_));
 sky130_fd_sc_hd__nor2_1 _10815_ (.A(_02881_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2b_1 _10816_ (.A_N(_02792_),
    .B(_02791_),
    .Y(_02884_));
 sky130_fd_sc_hd__a21oi_1 _10817_ (.A1(_02884_),
    .A2(_02803_),
    .B1(_02588_),
    .Y(_02885_));
 sky130_fd_sc_hd__xor2_1 _10818_ (.A(_02638_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__a21o_1 _10819_ (.A1(net425),
    .A2(_02883_),
    .B1(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__nand3_1 _10820_ (.A(_02863_),
    .B(_02886_),
    .C(_02883_),
    .Y(_02888_));
 sky130_fd_sc_hd__nand3_1 _10821_ (.A(_02480_),
    .B(_02485_),
    .C(_02763_),
    .Y(_02889_));
 sky130_fd_sc_hd__nor2_1 _10822_ (.A(_02480_),
    .B(_02789_),
    .Y(_02890_));
 sky130_fd_sc_hd__and2_0 _10823_ (.A(_02675_),
    .B(_02750_),
    .X(_02891_));
 sky130_fd_sc_hd__and3_1 _10824_ (.A(net392),
    .B(_02757_),
    .C(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__nand3_1 _10825_ (.A(_02890_),
    .B(_02763_),
    .C(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__or2_0 _10826_ (.A(_02892_),
    .B(_02889_),
    .X(_02894_));
 sky130_fd_sc_hd__nand3_1 _10827_ (.A(_02759_),
    .B(_02890_),
    .C(_02762_),
    .Y(_02895_));
 sky130_fd_sc_hd__o2111a_1 _10828_ (.A1(_02889_),
    .A2(net424),
    .B1(_02893_),
    .C1(_02894_),
    .D1(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__xnor2_1 _10829_ (.A(_02788_),
    .B(_02884_),
    .Y(_02897_));
 sky130_fd_sc_hd__a211oi_2 _10830_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02896_),
    .C1(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _10831_ (.A(_02879_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__clkbuf_4 _10832_ (.A(_02137_),
    .X(_02900_));
 sky130_fd_sc_hd__and2_0 _10833_ (.A(_02816_),
    .B(_02859_),
    .X(_02901_));
 sky130_fd_sc_hd__clkbuf_4 _10834_ (.A(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__or4_4 _10835_ (.A(_02788_),
    .B(_02793_),
    .C(_02802_),
    .D(_02806_),
    .X(_02903_));
 sky130_fd_sc_hd__nor3_1 _10836_ (.A(_07639_),
    .B(_07629_),
    .C(_02617_),
    .Y(_02904_));
 sky130_fd_sc_hd__nor3_1 _10837_ (.A(_07619_),
    .B(_07598_),
    .C(_02489_),
    .Y(_02905_));
 sky130_fd_sc_hd__nor3_1 _10838_ (.A(_07596_),
    .B(_07577_),
    .C(_02445_),
    .Y(_02906_));
 sky130_fd_sc_hd__nor2_8 _10839_ (.A(_07530_),
    .B(_02309_),
    .Y(_07548_));
 sky130_fd_sc_hd__nor3_1 _10840_ (.A(_07532_),
    .B(_07550_),
    .C(_07531_),
    .Y(_02907_));
 sky130_fd_sc_hd__nor2_1 _10841_ (.A(_00580_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(_07548_),
    .A1(_02908_),
    .S(_02402_),
    .X(_07571_));
 sky130_fd_sc_hd__nor3_1 _10843_ (.A(_07573_),
    .B(_07552_),
    .C(_02319_),
    .Y(_02909_));
 sky130_fd_sc_hd__o21ai_0 _10844_ (.A1(_02320_),
    .A2(_02909_),
    .B1(_02529_),
    .Y(_02910_));
 sky130_fd_sc_hd__o21a_1 _10845_ (.A1(_02529_),
    .A2(_07571_),
    .B1(_02910_),
    .X(_07594_));
 sky130_fd_sc_hd__nand2_1 _10846_ (.A(_02611_),
    .B(_07594_),
    .Y(_02911_));
 sky130_fd_sc_hd__o31ai_1 _10847_ (.A1(_02446_),
    .A2(net19),
    .A3(_02906_),
    .B1(_02911_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand2_1 _10848_ (.A(net7),
    .B(_07617_),
    .Y(_02912_));
 sky130_fd_sc_hd__o31ai_1 _10849_ (.A1(_02490_),
    .A2(net7),
    .A3(_02905_),
    .B1(_02912_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_1 _10850_ (.A(_02749_),
    .B(_07637_),
    .Y(_02913_));
 sky130_fd_sc_hd__o31ai_2 _10851_ (.A1(_02618_),
    .A2(_02749_),
    .A3(_02904_),
    .B1(_02913_),
    .Y(_07663_));
 sky130_fd_sc_hd__nor3_2 _10852_ (.A(_02880_),
    .B(_02903_),
    .C(_07663_),
    .Y(_02914_));
 sky130_fd_sc_hd__xor2_2 _10853_ (.A(_07665_),
    .B(net400),
    .X(_02915_));
 sky130_fd_sc_hd__a22oi_4 _10854_ (.A1(_02902_),
    .A2(_02914_),
    .B1(_02915_),
    .B2(net426),
    .Y(_02916_));
 sky130_fd_sc_hd__xnor2_1 _10855_ (.A(_02900_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__o211ai_4 _10856_ (.A1(_02702_),
    .A2(_02748_),
    .B1(_02766_),
    .C1(net411),
    .Y(_02918_));
 sky130_fd_sc_hd__and2_0 _10857_ (.A(_02772_),
    .B(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__inv_1 _10858_ (.A(_02919_),
    .Y(_02920_));
 sky130_fd_sc_hd__nand2b_1 _10859_ (.A_N(_02770_),
    .B(_02782_),
    .Y(_02921_));
 sky130_fd_sc_hd__nor2_1 _10860_ (.A(_02772_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__o21ai_0 _10861_ (.A1(_02881_),
    .A2(_02903_),
    .B1(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__nor2_1 _10862_ (.A(_02772_),
    .B(_02918_),
    .Y(_02924_));
 sky130_fd_sc_hd__a21oi_1 _10863_ (.A1(_02921_),
    .A2(_02919_),
    .B1(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__a211o_1 _10864_ (.A1(_02816_),
    .A2(_02859_),
    .B1(_02772_),
    .C1(_02921_),
    .X(_02926_));
 sky130_fd_sc_hd__o2111a_1 _10865_ (.A1(net423),
    .A2(_02920_),
    .B1(_02923_),
    .C1(_02925_),
    .D1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__nor3_1 _10866_ (.A(_02881_),
    .B(_02793_),
    .C(_02861_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _10867_ (.A(_02750_),
    .B(_02757_),
    .Y(_02929_));
 sky130_fd_sc_hd__a2111oi_2 _10868_ (.A1(_02881_),
    .A2(_02793_),
    .B1(_02927_),
    .C1(_02928_),
    .D1(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand3b_1 _10869_ (.A_N(_02823_),
    .B(_02845_),
    .C(_02858_),
    .Y(_02931_));
 sky130_fd_sc_hd__nor2_2 _10870_ (.A(_02881_),
    .B(_02903_),
    .Y(_02932_));
 sky130_fd_sc_hd__o21ai_0 _10871_ (.A1(_02811_),
    .A2(_02931_),
    .B1(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__o31ai_1 _10872_ (.A1(_02881_),
    .A2(_02882_),
    .A3(_02806_),
    .B1(_02802_),
    .Y(_02934_));
 sky130_fd_sc_hd__inv_1 _10873_ (.A(_02792_),
    .Y(_02935_));
 sky130_fd_sc_hd__a31oi_2 _10874_ (.A1(_02799_),
    .A2(_02791_),
    .A3(_02935_),
    .B1(_02804_),
    .Y(_02936_));
 sky130_fd_sc_hd__xnor2_2 _10875_ (.A(_02798_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__and4_1 _10876_ (.A(_02816_),
    .B(_02933_),
    .C(_02934_),
    .D(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__inv_1 _10877_ (.A(_07660_),
    .Y(_02939_));
 sky130_fd_sc_hd__xor2_2 _10878_ (.A(_07662_),
    .B(net389),
    .X(_02940_));
 sky130_fd_sc_hd__nor2_1 _10879_ (.A(_02749_),
    .B(_02768_),
    .Y(_02941_));
 sky130_fd_sc_hd__a21oi_1 _10880_ (.A1(_07640_),
    .A2(net18),
    .B1(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__xor2_1 _10881_ (.A(_02782_),
    .B(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__a32oi_4 _10882_ (.A1(_02939_),
    .A2(_02932_),
    .A3(_02902_),
    .B1(_02940_),
    .B2(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_4 _10883_ (.A1(net388),
    .A2(_02766_),
    .B1(_02918_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand4_1 _10884_ (.A(net397),
    .B(net431),
    .C(_07680_),
    .D(_07689_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand4_1 _10885_ (.A(_07669_),
    .B(_07716_),
    .C(_07683_),
    .D(_07686_),
    .Y(_02947_));
 sky130_fd_sc_hd__nor4_1 _10886_ (.A(_02944_),
    .B(_02945_),
    .C(_02946_),
    .D(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand4_1 _10887_ (.A(_02917_),
    .B(_02930_),
    .C(_02938_),
    .D(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__o21ai_2 _10888_ (.A1(_02899_),
    .A2(_02949_),
    .B1(_02858_),
    .Y(_02950_));
 sky130_fd_sc_hd__nor2_2 _10889_ (.A(_02843_),
    .B(_02844_),
    .Y(_02951_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_02829_),
    .B(_02834_),
    .Y(_02952_));
 sky130_fd_sc_hd__nand2_1 _10891_ (.A(_02952_),
    .B(_02839_),
    .Y(_02953_));
 sky130_fd_sc_hd__o2111a_1 _10892_ (.A1(_02811_),
    .A2(_02931_),
    .B1(_02816_),
    .C1(net402),
    .D1(_02807_),
    .X(_02954_));
 sky130_fd_sc_hd__xor2_1 _10893_ (.A(_02823_),
    .B(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__nor2_2 _10894_ (.A(_02953_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__o21a_1 _10895_ (.A1(_07669_),
    .A2(_07670_),
    .B1(_07677_),
    .X(_02957_));
 sky130_fd_sc_hd__o21a_1 _10896_ (.A1(_02957_),
    .A2(_07676_),
    .B1(_07674_),
    .X(_02958_));
 sky130_fd_sc_hd__o21ai_1 _10897_ (.A1(_02958_),
    .A2(_07673_),
    .B1(_07689_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand2b_1 _10898_ (.A_N(_07688_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__a21o_1 _10899_ (.A1(_02960_),
    .A2(_07686_),
    .B1(_07685_),
    .X(_02961_));
 sky130_fd_sc_hd__a21o_1 _10900_ (.A1(_02961_),
    .A2(_07683_),
    .B1(_07682_),
    .X(_02962_));
 sky130_fd_sc_hd__a21oi_4 _10901_ (.A1(_02962_),
    .A2(_07680_),
    .B1(_07679_),
    .Y(_02963_));
 sky130_fd_sc_hd__xnor2_1 _10902_ (.A(_07207_),
    .B(_02916_),
    .Y(_02964_));
 sky130_fd_sc_hd__a221oi_2 _10903_ (.A1(_02902_),
    .A2(_02914_),
    .B1(_02915_),
    .B2(net38),
    .C1(_02049_),
    .Y(_02965_));
 sky130_fd_sc_hd__nor3_1 _10904_ (.A(_02944_),
    .B(_02945_),
    .C(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__o221a_4 _10905_ (.A1(_02919_),
    .A2(_02924_),
    .B1(_02964_),
    .B2(_02963_),
    .C1(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__a21o_1 _10906_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02897_),
    .X(_02968_));
 sky130_fd_sc_hd__nor4_1 _10907_ (.A(_02770_),
    .B(_02783_),
    .C(_02876_),
    .D(net403),
    .Y(_02969_));
 sky130_fd_sc_hd__a21boi_0 _10908_ (.A1(_02784_),
    .A2(net38),
    .B1_N(_02876_),
    .Y(_02970_));
 sky130_fd_sc_hd__nor4b_1 _10909_ (.A(_02789_),
    .B(_02764_),
    .C(_02756_),
    .D_N(_02891_),
    .Y(_02971_));
 sky130_fd_sc_hd__o21ai_1 _10910_ (.A1(_02969_),
    .A2(_02970_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_2 _10911_ (.A1(_02881_),
    .A2(_02793_),
    .B1(_02928_),
    .Y(_02973_));
 sky130_fd_sc_hd__nand2_1 _10912_ (.A(_02932_),
    .B(_02931_),
    .Y(_02974_));
 sky130_fd_sc_hd__and4_1 _10913_ (.A(_02816_),
    .B(_02934_),
    .C(_02937_),
    .D(_02974_),
    .X(_02975_));
 sky130_fd_sc_hd__and4bb_1 _10914_ (.A_N(_02968_),
    .B_N(_02972_),
    .C(_02973_),
    .D(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__nand4_4 _10915_ (.A(_02951_),
    .B(_02956_),
    .C(_02967_),
    .D(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__or2_4 _10916_ (.A(_02950_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__buf_6 _10917_ (.A(_02978_),
    .X(_00552_));
 sky130_fd_sc_hd__xnor2_1 _10918_ (.A(_07680_),
    .B(net408),
    .Y(_02979_));
 sky130_fd_sc_hd__nand2_1 _10919_ (.A(_00552_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__o21ai_0 _10920_ (.A1(_07678_),
    .A2(net35),
    .B1(_02980_),
    .Y(_07691_));
 sky130_fd_sc_hd__nor3_1 _10921_ (.A(_07653_),
    .B(_07655_),
    .C(_02775_),
    .Y(_02981_));
 sky130_fd_sc_hd__or2_0 _10922_ (.A(_02776_),
    .B(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__nor3_1 _10923_ (.A(_07633_),
    .B(_07623_),
    .C(_02615_),
    .Y(_02983_));
 sky130_fd_sc_hd__nor3_1 _10924_ (.A(_07602_),
    .B(_07604_),
    .C(_02487_),
    .Y(_02984_));
 sky130_fd_sc_hd__nor3_1 _10925_ (.A(_07575_),
    .B(_07581_),
    .C(_07574_),
    .Y(_02985_));
 sky130_fd_sc_hd__nor2_1 _10926_ (.A(_02444_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__nor2_4 _10927_ (.A(_07555_),
    .B(_02520_),
    .Y(_07579_));
 sky130_fd_sc_hd__mux2_4 _10928_ (.A0(_02986_),
    .A1(_07579_),
    .S(_02611_),
    .X(_07600_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_02626_),
    .B(_07600_),
    .Y(_02987_));
 sky130_fd_sc_hd__o31ai_1 _10930_ (.A1(_02488_),
    .A2(_02626_),
    .A3(_02984_),
    .B1(_02987_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_1 _10931_ (.A(net18),
    .B(_07631_),
    .Y(_02988_));
 sky130_fd_sc_hd__o31ai_1 _10932_ (.A1(_02616_),
    .A2(net18),
    .A3(_02983_),
    .B1(_02988_),
    .Y(_07651_));
 sky130_fd_sc_hd__nor2_1 _10933_ (.A(net434),
    .B(_07651_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21oi_1 _10934_ (.A1(net434),
    .A2(_02982_),
    .B1(_02989_),
    .Y(_07681_));
 sky130_fd_sc_hd__nor2b_2 _10935_ (.A(_07668_),
    .B_N(net398),
    .Y(_02990_));
 sky130_fd_sc_hd__o21ai_1 _10936_ (.A1(_07676_),
    .A2(_02990_),
    .B1(net432),
    .Y(_02991_));
 sky130_fd_sc_hd__nand2b_1 _10937_ (.A_N(_07673_),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__a21o_1 _10938_ (.A1(_02992_),
    .A2(_07689_),
    .B1(_07688_),
    .X(_02993_));
 sky130_fd_sc_hd__a21o_1 _10939_ (.A1(_02993_),
    .A2(_07686_),
    .B1(_07685_),
    .X(_02994_));
 sky130_fd_sc_hd__xnor2_1 _10940_ (.A(_07683_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__nand2_2 _10941_ (.A(_00552_),
    .B(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__o21ai_1 _10942_ (.A1(net35),
    .A2(_07681_),
    .B1(_02996_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor3_1 _10943_ (.A(_07624_),
    .B(_07626_),
    .C(_02614_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor3_1 _10944_ (.A(_07607_),
    .B(_07605_),
    .C(_07606_),
    .Y(_02998_));
 sky130_fd_sc_hd__nor2_2 _10945_ (.A(_07575_),
    .B(_02611_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand2_1 _10946_ (.A(_02626_),
    .B(_07603_),
    .Y(_02999_));
 sky130_fd_sc_hd__o31ai_4 _10947_ (.A1(_02487_),
    .A2(_02626_),
    .A3(_02998_),
    .B1(_02999_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand2_1 _10948_ (.A(_02866_),
    .B(_07622_),
    .Y(_03000_));
 sky130_fd_sc_hd__o31ai_1 _10949_ (.A1(_02615_),
    .A2(_02866_),
    .A3(_02997_),
    .B1(_03000_),
    .Y(_07654_));
 sky130_fd_sc_hd__nor3_1 _10950_ (.A(_07656_),
    .B(_07658_),
    .C(_02774_),
    .Y(_03001_));
 sky130_fd_sc_hd__o21ai_0 _10951_ (.A1(_02775_),
    .A2(_03001_),
    .B1(_00553_),
    .Y(_03002_));
 sky130_fd_sc_hd__o21a_1 _10952_ (.A1(_00553_),
    .A2(_07654_),
    .B1(_03002_),
    .X(_07684_));
 sky130_fd_sc_hd__xnor2_1 _10953_ (.A(_07686_),
    .B(net409),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_2 _10954_ (.A(_00552_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__o21ai_2 _10955_ (.A1(_00552_),
    .A2(_07684_),
    .B1(_03004_),
    .Y(_07699_));
 sky130_fd_sc_hd__nor3_1 _10956_ (.A(_07627_),
    .B(_07621_),
    .C(_07620_),
    .Y(_03005_));
 sky130_fd_sc_hd__nor2_4 _10957_ (.A(_07607_),
    .B(_02626_),
    .Y(_07625_));
 sky130_fd_sc_hd__nand2_1 _10958_ (.A(_02866_),
    .B(_07625_),
    .Y(_03006_));
 sky130_fd_sc_hd__o31ai_1 _10959_ (.A1(_02614_),
    .A2(_02866_),
    .A3(_03005_),
    .B1(_03006_),
    .Y(_07657_));
 sky130_fd_sc_hd__nor3_1 _10960_ (.A(_07659_),
    .B(_07644_),
    .C(_02773_),
    .Y(_03007_));
 sky130_fd_sc_hd__o21ai_0 _10961_ (.A1(_02774_),
    .A2(_03007_),
    .B1(_02863_),
    .Y(_03008_));
 sky130_fd_sc_hd__o21a_1 _10962_ (.A1(_00553_),
    .A2(_07657_),
    .B1(_03008_),
    .X(_07687_));
 sky130_fd_sc_hd__xnor2_1 _10963_ (.A(_07689_),
    .B(_02992_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2_1 _10964_ (.A(_00552_),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__o21ai_1 _10965_ (.A1(net35),
    .A2(_07687_),
    .B1(_03010_),
    .Y(_07703_));
 sky130_fd_sc_hd__nor2_8 _10966_ (.A(_07621_),
    .B(_02866_),
    .Y(_07643_));
 sky130_fd_sc_hd__nor3_1 _10967_ (.A(_07645_),
    .B(_07647_),
    .C(_07646_),
    .Y(_03011_));
 sky130_fd_sc_hd__o21ai_2 _10968_ (.A1(_02773_),
    .A2(_03011_),
    .B1(_00553_),
    .Y(_03012_));
 sky130_fd_sc_hd__o21a_1 _10969_ (.A1(_00553_),
    .A2(_07643_),
    .B1(_03012_),
    .X(_07672_));
 sky130_fd_sc_hd__nor3_1 _10970_ (.A(net432),
    .B(_07676_),
    .C(net422),
    .Y(_03013_));
 sky130_fd_sc_hd__nor2_1 _10971_ (.A(net416),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__mux2i_1 _10972_ (.A0(net417),
    .A1(_03014_),
    .S(net35),
    .Y(_07707_));
 sky130_fd_sc_hd__nor2_4 _10973_ (.A(\butterfly_count[2] ),
    .B(_02863_),
    .Y(_03015_));
 sky130_fd_sc_hd__a21oi_4 _10974_ (.A1(_02863_),
    .A2(_07647_),
    .B1(_03015_),
    .Y(_07675_));
 sky130_fd_sc_hd__or3_1 _10975_ (.A(_02927_),
    .B(_02950_),
    .C(_02977_),
    .X(_03016_));
 sky130_fd_sc_hd__xnor2_1 _10976_ (.A(_07662_),
    .B(_02780_),
    .Y(_03017_));
 sky130_fd_sc_hd__nor3_1 _10977_ (.A(_02939_),
    .B(_02881_),
    .C(_02903_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_1 _10978_ (.A(_07683_),
    .B(_02994_),
    .Y(_03019_));
 sky130_fd_sc_hd__a221oi_1 _10979_ (.A1(net37),
    .A2(_03017_),
    .B1(_03018_),
    .B2(_02902_),
    .C1(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__o21a_1 _10980_ (.A1(_07682_),
    .A2(_03020_),
    .B1(_07680_),
    .X(_03021_));
 sky130_fd_sc_hd__o21ai_1 _10981_ (.A1(_07679_),
    .A2(_03021_),
    .B1(_02917_),
    .Y(_03022_));
 sky130_fd_sc_hd__and2_0 _10982_ (.A(_02966_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__o31ai_1 _10983_ (.A1(_02881_),
    .A2(_02903_),
    .A3(_02902_),
    .B1(_02934_),
    .Y(_03024_));
 sky130_fd_sc_hd__or4_1 _10984_ (.A(_02881_),
    .B(_02882_),
    .C(_02861_),
    .D(_02886_),
    .X(_03025_));
 sky130_fd_sc_hd__xor2_1 _10985_ (.A(_02937_),
    .B(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__nand3_1 _10986_ (.A(_02879_),
    .B(_02898_),
    .C(_02930_),
    .Y(_03027_));
 sky130_fd_sc_hd__nor4_1 _10987_ (.A(_02967_),
    .B(_03024_),
    .C(_03026_),
    .D(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_02750_),
    .B(_02876_),
    .Y(_03029_));
 sky130_fd_sc_hd__a21oi_1 _10989_ (.A1(net394),
    .A2(net37),
    .B1(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nor2_1 _10990_ (.A(_02969_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2b_1 _10991_ (.A(_03031_),
    .B_N(_02967_),
    .Y(_03032_));
 sky130_fd_sc_hd__a21oi_1 _10992_ (.A1(_03023_),
    .A2(_03028_),
    .B1(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_02977_),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__nor2_1 _10994_ (.A(net405),
    .B(_02940_),
    .Y(_03035_));
 sky130_fd_sc_hd__and2_0 _10995_ (.A(_02902_),
    .B(_03018_),
    .X(_03036_));
 sky130_fd_sc_hd__or3_1 _10996_ (.A(_02965_),
    .B(_03035_),
    .C(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__nor2_1 _10997_ (.A(_02782_),
    .B(_02942_),
    .Y(_03038_));
 sky130_fd_sc_hd__and3_1 _10998_ (.A(_02782_),
    .B(net37),
    .C(_02942_),
    .X(_03039_));
 sky130_fd_sc_hd__mux2i_1 _10999_ (.A0(_03038_),
    .A1(_03039_),
    .S(_02945_),
    .Y(_03040_));
 sky130_fd_sc_hd__nor2_1 _11000_ (.A(_03037_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_1 _11001_ (.A(_02945_),
    .B(_02963_),
    .Y(_03042_));
 sky130_fd_sc_hd__nor4_1 _11002_ (.A(_02965_),
    .B(_03035_),
    .C(_03036_),
    .D(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__nor2_1 _11003_ (.A(_02945_),
    .B(_02963_),
    .Y(_03044_));
 sky130_fd_sc_hd__o221ai_1 _11004_ (.A1(_07679_),
    .A2(_03021_),
    .B1(_03043_),
    .B2(_03044_),
    .C1(_02917_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2b_1 _11005_ (.A_N(_02945_),
    .B(_03037_),
    .Y(_03046_));
 sky130_fd_sc_hd__a211oi_1 _11006_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03038_),
    .C1(_03039_),
    .Y(_03047_));
 sky130_fd_sc_hd__a21oi_1 _11007_ (.A1(_03022_),
    .A2(_03041_),
    .B1(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand2_1 _11008_ (.A(_02966_),
    .B(_03022_),
    .Y(_03049_));
 sky130_fd_sc_hd__nor2_1 _11009_ (.A(_02927_),
    .B(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_02902_),
    .B(_03018_),
    .Y(_03051_));
 sky130_fd_sc_hd__o21ai_1 _11011_ (.A1(net406),
    .A2(_02940_),
    .B1(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2b_1 _11012_ (.A_N(_07682_),
    .B(_03019_),
    .Y(_03053_));
 sky130_fd_sc_hd__a21oi_1 _11013_ (.A1(_07680_),
    .A2(_03053_),
    .B1(_07679_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _11014_ (.A(net37),
    .B(_02940_),
    .Y(_03055_));
 sky130_fd_sc_hd__a31oi_1 _11015_ (.A1(_02939_),
    .A2(_02932_),
    .A3(_02902_),
    .B1(net391),
    .Y(_03056_));
 sky130_fd_sc_hd__a22o_1 _11016_ (.A1(net391),
    .A2(_03051_),
    .B1(_03055_),
    .B2(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__nand2_1 _11017_ (.A(_02963_),
    .B(_03035_),
    .Y(_03058_));
 sky130_fd_sc_hd__a211oi_1 _11018_ (.A1(_03057_),
    .A2(_03058_),
    .B1(_02900_),
    .C1(_03054_),
    .Y(_03059_));
 sky130_fd_sc_hd__a311oi_1 _11019_ (.A1(_02900_),
    .A2(_03052_),
    .A3(_03054_),
    .B1(_03059_),
    .C1(_02916_),
    .Y(_03060_));
 sky130_fd_sc_hd__a21o_1 _11020_ (.A1(_07680_),
    .A2(_03053_),
    .B1(_07679_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _11021_ (.A(_02900_),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_1 _11022_ (.A(_02900_),
    .B(_03054_),
    .Y(_03063_));
 sky130_fd_sc_hd__o22ai_1 _11023_ (.A1(_02963_),
    .A2(_03062_),
    .B1(_03063_),
    .B2(_02049_),
    .Y(_03064_));
 sky130_fd_sc_hd__nor2_1 _11024_ (.A(_03052_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand3_1 _11025_ (.A(_02900_),
    .B(_02963_),
    .C(_03061_),
    .Y(_03066_));
 sky130_fd_sc_hd__o21ai_0 _11026_ (.A1(_02900_),
    .A2(_03061_),
    .B1(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__a21boi_0 _11027_ (.A1(_02049_),
    .A2(_03067_),
    .B1_N(_03052_),
    .Y(_03068_));
 sky130_fd_sc_hd__o21ai_0 _11028_ (.A1(_03065_),
    .A2(_03068_),
    .B1(_02916_),
    .Y(_03069_));
 sky130_fd_sc_hd__nor2_1 _11029_ (.A(_02968_),
    .B(_02972_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand4_1 _11030_ (.A(_02937_),
    .B(_02967_),
    .C(_03070_),
    .D(_02973_),
    .Y(_03071_));
 sky130_fd_sc_hd__nand4b_1 _11031_ (.A_N(_03060_),
    .B(_03069_),
    .C(_03071_),
    .D(_02973_),
    .Y(_03072_));
 sky130_fd_sc_hd__or3_1 _11032_ (.A(_02916_),
    .B(_02944_),
    .C(_02945_),
    .X(_03073_));
 sky130_fd_sc_hd__o32a_1 _11033_ (.A1(_03048_),
    .A2(_03050_),
    .A3(_03072_),
    .B1(_03073_),
    .B2(_02978_),
    .X(_03074_));
 sky130_fd_sc_hd__a31oi_1 _11034_ (.A1(_02796_),
    .A2(_02741_),
    .A3(_02748_),
    .B1(_02830_),
    .Y(_03075_));
 sky130_fd_sc_hd__a31oi_2 _11035_ (.A1(_02796_),
    .A2(_02741_),
    .A3(_02830_),
    .B1(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__or2_1 _11036_ (.A(_02823_),
    .B(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__inv_1 _11037_ (.A(_02954_),
    .Y(_03078_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(_03078_),
    .B(_03076_),
    .Y(_03079_));
 sky130_fd_sc_hd__and4_1 _11039_ (.A(_02879_),
    .B(_02898_),
    .C(_02930_),
    .D(_02938_),
    .X(_03080_));
 sky130_fd_sc_hd__and3_1 _11040_ (.A(_02966_),
    .B(_03022_),
    .C(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__o21ai_0 _11041_ (.A1(_02950_),
    .A2(_02977_),
    .B1(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__mux2i_1 _11042_ (.A0(_03077_),
    .A1(_03079_),
    .S(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__o41ai_1 _11043_ (.A1(_03026_),
    .A2(_03049_),
    .A3(_03027_),
    .A4(_03032_),
    .B1(_03024_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand3_1 _11044_ (.A(_02967_),
    .B(_03070_),
    .C(_02973_),
    .Y(_03085_));
 sky130_fd_sc_hd__a22oi_1 _11045_ (.A1(_02927_),
    .A2(_03049_),
    .B1(_03085_),
    .B2(_03026_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux2i_1 _11046_ (.A0(_02932_),
    .A1(_02974_),
    .S(_02815_),
    .Y(_03087_));
 sky130_fd_sc_hd__nand2_1 _11047_ (.A(_02856_),
    .B(_02731_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor3_1 _11048_ (.A(_02702_),
    .B(_02825_),
    .C(_02830_),
    .Y(_03089_));
 sky130_fd_sc_hd__nand3_1 _11049_ (.A(_03088_),
    .B(_03089_),
    .C(_02828_),
    .Y(_03090_));
 sky130_fd_sc_hd__nand4_2 _11050_ (.A(_07693_),
    .B(_07697_),
    .C(_07701_),
    .D(_07705_),
    .Y(_03091_));
 sky130_fd_sc_hd__a21oi_2 _11051_ (.A1(_07701_),
    .A2(_07704_),
    .B1(_07700_),
    .Y(_03092_));
 sky130_fd_sc_hd__nor2b_2 _11052_ (.A(_03092_),
    .B_N(_07697_),
    .Y(_03093_));
 sky130_fd_sc_hd__o21ai_1 _11053_ (.A1(_03093_),
    .A2(_07696_),
    .B1(_07693_),
    .Y(_03094_));
 sky130_fd_sc_hd__nand2b_1 _11054_ (.A_N(_07692_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a41oi_2 _11055_ (.A1(_07709_),
    .A2(_07715_),
    .A3(_07713_),
    .A4(_07718_),
    .B1(_03091_),
    .Y(_03096_));
 sky130_fd_sc_hd__a21oi_4 _11056_ (.A1(_03095_),
    .A2(_03091_),
    .B1(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__a21oi_2 _11057_ (.A1(_02840_),
    .A2(_03090_),
    .B1(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__or3b_1 _11058_ (.A(_02857_),
    .B(_02847_),
    .C_N(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_02823_),
    .B(_03076_),
    .Y(_03100_));
 sky130_fd_sc_hd__o21ai_0 _11060_ (.A1(_03078_),
    .A2(_03077_),
    .B1(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__or4_4 _11061_ (.A(_02811_),
    .B(_03099_),
    .C(_03101_),
    .D(_03087_),
    .X(_03102_));
 sky130_fd_sc_hd__nand4_1 _11062_ (.A(_02675_),
    .B(net392),
    .C(_02876_),
    .D(net37),
    .Y(_03103_));
 sky130_fd_sc_hd__xor2_1 _11063_ (.A(_02756_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__nor3_1 _11064_ (.A(_02760_),
    .B(_02750_),
    .C(_02756_),
    .Y(_03105_));
 sky130_fd_sc_hd__a21oi_1 _11065_ (.A1(_02750_),
    .A2(_03104_),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nor2b_1 _11066_ (.A(_02967_),
    .B_N(_03031_),
    .Y(_03107_));
 sky130_fd_sc_hd__nor3_1 _11067_ (.A(_02823_),
    .B(_02953_),
    .C(_03078_),
    .Y(_03108_));
 sky130_fd_sc_hd__xor2_1 _11068_ (.A(_02951_),
    .B(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_02956_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nor4_4 _11070_ (.A(_03110_),
    .B(_03106_),
    .C(_03107_),
    .D(_03102_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _11071_ (.A(_02967_),
    .B(_02976_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2b_1 _11072_ (.A_N(_02955_),
    .B(_02951_),
    .Y(_03113_));
 sky130_fd_sc_hd__a21boi_0 _11073_ (.A1(_03112_),
    .A2(_03113_),
    .B1_N(_02898_),
    .Y(_03114_));
 sky130_fd_sc_hd__nand4_2 _11074_ (.A(_03084_),
    .B(_03111_),
    .C(_03086_),
    .D(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__a2111oi_4 _11075_ (.A1(_03016_),
    .A2(_03034_),
    .B1(_03115_),
    .C1(_03083_),
    .D1(_03074_),
    .Y(_03116_));
 sky130_fd_sc_hd__nor3_2 _11076_ (.A(\butterfly_count[1] ),
    .B(_02950_),
    .C(_02977_),
    .Y(_03117_));
 sky130_fd_sc_hd__a21oi_4 _11077_ (.A1(_07669_),
    .A2(net395),
    .B1(_03117_),
    .Y(_05893_));
 sky130_fd_sc_hd__nand3_1 _11078_ (.A(_07709_),
    .B(_07713_),
    .C(_05907_),
    .Y(_03118_));
 sky130_fd_sc_hd__nand2_1 _11079_ (.A(_07715_),
    .B(_07713_),
    .Y(_03119_));
 sky130_fd_sc_hd__o21bai_1 _11080_ (.A1(_07719_),
    .A2(_03119_),
    .B1_N(_07712_),
    .Y(_03120_));
 sky130_fd_sc_hd__a211oi_1 _11081_ (.A1(_07709_),
    .A2(_03120_),
    .B1(_03095_),
    .C1(_07708_),
    .Y(_03121_));
 sky130_fd_sc_hd__o21ai_4 _11082_ (.A1(_05893_),
    .A2(_03118_),
    .B1(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__o2111ai_1 _11083_ (.A1(_02899_),
    .A2(_02949_),
    .B1(_02956_),
    .C1(_02951_),
    .D1(_02858_),
    .Y(_03123_));
 sky130_fd_sc_hd__a31oi_1 _11084_ (.A1(_02967_),
    .A2(_02976_),
    .A3(_03123_),
    .B1(_02954_),
    .Y(_03124_));
 sky130_fd_sc_hd__or2_0 _11085_ (.A(_03089_),
    .B(_02828_),
    .X(_03125_));
 sky130_fd_sc_hd__o211ai_1 _11086_ (.A1(_03077_),
    .A2(_03124_),
    .B1(_03125_),
    .C1(_03090_),
    .Y(_03126_));
 sky130_fd_sc_hd__a211o_1 _11087_ (.A1(_03090_),
    .A2(_03125_),
    .B1(_03124_),
    .C1(_03077_),
    .X(_03127_));
 sky130_fd_sc_hd__nor2_1 _11088_ (.A(_02927_),
    .B(_03029_),
    .Y(_03128_));
 sky130_fd_sc_hd__o211ai_1 _11089_ (.A1(_02950_),
    .A2(_02977_),
    .B1(_03023_),
    .C1(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__xor2_1 _11090_ (.A(_02879_),
    .B(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__a21oi_1 _11091_ (.A1(_03126_),
    .A2(_03127_),
    .B1(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__a211oi_1 _11092_ (.A1(_02846_),
    .A2(_02847_),
    .B1(_02851_),
    .C1(_02855_),
    .Y(_03132_));
 sky130_fd_sc_hd__o211a_1 _11093_ (.A1(_02950_),
    .A2(_02977_),
    .B1(_03081_),
    .C1(_02956_),
    .X(_03133_));
 sky130_fd_sc_hd__o21ai_0 _11094_ (.A1(_03108_),
    .A2(_03133_),
    .B1(_02951_),
    .Y(_03134_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(_03132_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand4_4 _11096_ (.A(_03122_),
    .B(_03116_),
    .C(_03131_),
    .D(_03135_),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_1 _11097_ (.A(\state[0] ),
    .Y(_03136_));
 sky130_fd_sc_hd__buf_4 _11098_ (.A(\state[2] ),
    .X(_03137_));
 sky130_fd_sc_hd__nand2_2 _11099_ (.A(net91),
    .B(_07833_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand2_1 _11100_ (.A(_03137_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__o21ai_0 _11101_ (.A1(_03136_),
    .A2(_00557_),
    .B1(_03139_),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_1 _11102_ (.A(\state[2] ),
    .Y(_03140_));
 sky130_fd_sc_hd__clkbuf_4 _11103_ (.A(\state[1] ),
    .X(_03141_));
 sky130_fd_sc_hd__clkbuf_8 _11104_ (.A(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_03142_),
    .B(_07819_),
    .Y(_03143_));
 sky130_fd_sc_hd__o21ai_0 _11106_ (.A1(_03140_),
    .A2(_03138_),
    .B1(_03143_),
    .Y(_00005_));
 sky130_fd_sc_hd__nor2b_2 _11107_ (.A(\butterfly_count[2] ),
    .B_N(\state[1] ),
    .Y(_03144_));
 sky130_fd_sc_hd__nand3_2 _11108_ (.A(_07819_),
    .B(net354),
    .C(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__inv_8 _11109_ (.A(_03145_),
    .Y(_00007_));
 sky130_fd_sc_hd__buf_6 _11110_ (.A(net519),
    .X(_03146_));
 sky130_fd_sc_hd__buf_6 _11111_ (.A(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__buf_6 _11112_ (.A(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__buf_12 _11113_ (.A(net514),
    .X(_03149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__inv_4 _11115_ (.A(net526),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_8 _11116_ (.A(_03151_),
    .B(net589),
    .Y(_03152_));
 sky130_fd_sc_hd__buf_8 _11117_ (.A(net526),
    .X(_03153_));
 sky130_fd_sc_hd__nand2b_4 _11118_ (.A_N(net520),
    .B(net515),
    .Y(_03154_));
 sky130_fd_sc_hd__buf_6 _11119_ (.A(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__nor2_8 _11120_ (.A(_03155_),
    .B(net633),
    .Y(_03156_));
 sky130_fd_sc_hd__a32oi_2 _11121_ (.A1(\samples_real[5][0] ),
    .A2(_03148_),
    .A3(_03152_),
    .B1(_03156_),
    .B2(\samples_real[2][0] ),
    .Y(_03157_));
 sky130_fd_sc_hd__buf_6 _11122_ (.A(_03151_),
    .X(_03158_));
 sky130_fd_sc_hd__nor2_1 _11123_ (.A(_03158_),
    .B(_03155_),
    .Y(_03159_));
 sky130_fd_sc_hd__nor2_8 _11124_ (.A(net590),
    .B(net572),
    .Y(_03160_));
 sky130_fd_sc_hd__and2_4 _11125_ (.A(_03160_),
    .B(_03146_),
    .X(_03161_));
 sky130_fd_sc_hd__buf_12 clone64 (.A(_05106_),
    .X(net64));
 sky130_fd_sc_hd__a22oi_4 _11127_ (.A1(\samples_real[3][0] ),
    .A2(_03159_),
    .B1(\samples_real[4][0] ),
    .B2(net615),
    .Y(_03163_));
 sky130_fd_sc_hd__buf_12 _11128_ (.A(_03149_),
    .X(_03164_));
 sky130_fd_sc_hd__buf_12 _11129_ (.A(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__buf_6 _11130_ (.A(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__buf_12 _11131_ (.A(_03153_),
    .X(_03167_));
 sky130_fd_sc_hd__mux2_4 _11132_ (.A0(\samples_real[6][0] ),
    .A1(\samples_real[7][0] ),
    .S(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__buf_6 _11133_ (.A(_03147_),
    .X(_03169_));
 sky130_fd_sc_hd__buf_12 _11134_ (.A(_03165_),
    .X(_03170_));
 sky130_fd_sc_hd__nor2_2 _11135_ (.A(_03158_),
    .B(\samples_real[1][0] ),
    .Y(_03171_));
 sky130_fd_sc_hd__nor3_4 _11136_ (.A(_03169_),
    .B(_03170_),
    .C(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__a31oi_4 _11137_ (.A1(_03168_),
    .A2(_03166_),
    .A3(_03148_),
    .B1(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__or3_1 _11138_ (.A(net519),
    .B(net514),
    .C(\idx1[0] ),
    .X(_03174_));
 sky130_fd_sc_hd__buf_6 _11139_ (.A(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_6 _11140_ (.A(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__buf_8 _11141_ (.A(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__nor2_8 _11142_ (.A(\samples_real[0][0] ),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__a31oi_4 _11143_ (.A1(_03157_),
    .A2(_03173_),
    .A3(_03163_),
    .B1(_03178_),
    .Y(_07732_));
 sky130_fd_sc_hd__inv_2 _11144_ (.A(net569),
    .Y(_07734_));
 sky130_fd_sc_hd__clkbuf_2 rebuffer230 (.A(_03170_),
    .X(net601));
 sky130_fd_sc_hd__mux4_2 _11146_ (.A0(\samples_real[0][1] ),
    .A1(\samples_real[2][1] ),
    .A2(\samples_real[1][1] ),
    .A3(\samples_real[3][1] ),
    .S0(net586),
    .S1(net580),
    .X(_03180_));
 sky130_fd_sc_hd__buf_12 _11147_ (.A(_03153_),
    .X(_03181_));
 sky130_fd_sc_hd__buf_8 _11148_ (.A(_03149_),
    .X(_03182_));
 sky130_fd_sc_hd__buf_6 _11149_ (.A(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__mux4_1 _11150_ (.A0(\samples_real[4][1] ),
    .A1(\samples_real[5][1] ),
    .A2(\samples_real[6][1] ),
    .A3(\samples_real[7][1] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__clkbuf_8 _11151_ (.A(_03169_),
    .X(_03185_));
 sky130_fd_sc_hd__mux2_4 _11152_ (.A0(_03180_),
    .A1(_03184_),
    .S(_03185_),
    .X(_05887_));
 sky130_fd_sc_hd__inv_1 _11153_ (.A(_05887_),
    .Y(_05883_));
 sky130_fd_sc_hd__clkinv_8 _11154_ (.A(net53),
    .Y(_05882_));
 sky130_fd_sc_hd__inv_2 _11155_ (.A(_05891_),
    .Y(_05888_));
 sky130_fd_sc_hd__mux2i_1 _11156_ (.A0(_07716_),
    .A1(_07718_),
    .S(_00551_),
    .Y(_00554_));
 sky130_fd_sc_hd__inv_1 _11157_ (.A(_05893_),
    .Y(_03186_));
 sky130_fd_sc_hd__mux2i_1 _11158_ (.A0(_03186_),
    .A1(_05896_),
    .S(_00551_),
    .Y(_00555_));
 sky130_fd_sc_hd__nor2b_1 _11159_ (.A(net399),
    .B_N(_07668_),
    .Y(_03187_));
 sky130_fd_sc_hd__o21ai_0 _11160_ (.A1(_02990_),
    .A2(_03187_),
    .B1(net395),
    .Y(_03188_));
 sky130_fd_sc_hd__o21ai_1 _11161_ (.A1(net395),
    .A2(net427),
    .B1(_03188_),
    .Y(_07711_));
 sky130_fd_sc_hd__xnor2_1 _11162_ (.A(_05895_),
    .B(_07713_),
    .Y(_03189_));
 sky130_fd_sc_hd__mux2i_1 _11163_ (.A0(_07711_),
    .A1(_03189_),
    .S(_00551_),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_4 _11164_ (.A(\stage[1] ),
    .Y(_07804_));
 sky130_fd_sc_hd__mux2i_2 _11165_ (.A0(\butterfly_in_group[0] ),
    .A1(\butterfly_in_group[1] ),
    .S(\stage[0] ),
    .Y(_03190_));
 sky130_fd_sc_hd__inv_8 _11166_ (.A(\stage[0] ),
    .Y(_07803_));
 sky130_fd_sc_hd__nand4_1 _11167_ (.A(_00562_),
    .B(_07803_),
    .C(\butterfly_in_group[2] ),
    .D(_07804_),
    .Y(_03191_));
 sky130_fd_sc_hd__o31ai_4 _11168_ (.A1(_00562_),
    .A2(_07804_),
    .A3(_03190_),
    .B1(_03191_),
    .Y(_05877_));
 sky130_fd_sc_hd__mux2i_4 _11169_ (.A0(\twiddle_idx[0] ),
    .A1(_05877_),
    .S(_00007_),
    .Y(_03192_));
 sky130_fd_sc_hd__inv_1 _11170_ (.A(_03192_),
    .Y(_00000_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\butterfly_in_group[1] ),
    .A1(\butterfly_in_group[2] ),
    .S(\stage[0] ),
    .X(_03193_));
 sky130_fd_sc_hd__nand2_1 _11172_ (.A(\stage[1] ),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nand3_1 _11173_ (.A(\stage[0] ),
    .B(\butterfly_in_group[0] ),
    .C(_07804_),
    .Y(_03195_));
 sky130_fd_sc_hd__a21oi_2 _11174_ (.A1(_03194_),
    .A2(_03195_),
    .B1(_00562_),
    .Y(_05878_));
 sky130_fd_sc_hd__mux2i_4 _11175_ (.A0(\twiddle_idx[1] ),
    .A1(_05878_),
    .S(_00007_),
    .Y(_00002_));
 sky130_fd_sc_hd__nand2_1 _11176_ (.A(_03192_),
    .B(_00002_),
    .Y(_00023_));
 sky130_fd_sc_hd__inv_1 _11177_ (.A(_00023_),
    .Y(_00020_));
 sky130_fd_sc_hd__nor2_1 _11178_ (.A(_03192_),
    .B(_00002_),
    .Y(_00022_));
 sky130_fd_sc_hd__or2_0 _11179_ (.A(_00020_),
    .B(_00022_),
    .X(_00001_));
 sky130_fd_sc_hd__nor3_4 _11180_ (.A(_03146_),
    .B(_03158_),
    .C(_03164_),
    .Y(_03196_));
 sky130_fd_sc_hd__a22oi_4 _11181_ (.A1(net536),
    .A2(\samples_imag[2][0] ),
    .B1(_03196_),
    .B2(\samples_imag[1][0] ),
    .Y(_03197_));
 sky130_fd_sc_hd__and3_2 _11182_ (.A(_03146_),
    .B(net516),
    .C(net65),
    .X(_03198_));
 sky130_fd_sc_hd__a22oi_4 _11183_ (.A1(\samples_imag[4][0] ),
    .A2(net553),
    .B1(_03198_),
    .B2(\samples_imag[7][0] ),
    .Y(_03199_));
 sky130_fd_sc_hd__and3_4 _11184_ (.A(net516),
    .B(net65),
    .C(\samples_imag[3][0] ),
    .X(_03200_));
 sky130_fd_sc_hd__inv_4 _11185_ (.A(_03149_),
    .Y(_03201_));
 sky130_fd_sc_hd__nor2_4 _11186_ (.A(_03201_),
    .B(net575),
    .Y(_03202_));
 sky130_fd_sc_hd__a22oi_1 _11187_ (.A1(\samples_imag[5][0] ),
    .A2(_03152_),
    .B1(_03202_),
    .B2(\samples_imag[6][0] ),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _11188_ (.A(_03147_),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__o31ai_4 _11189_ (.A1(_03146_),
    .A2(_03200_),
    .A3(net555),
    .B1(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_1 _11190_ (.A(\samples_imag[0][0] ),
    .B(_03175_),
    .Y(_03206_));
 sky130_fd_sc_hd__a31oi_4 _11191_ (.A1(_03199_),
    .A2(_03197_),
    .A3(_03205_),
    .B1(_03206_),
    .Y(_07846_));
 sky130_fd_sc_hd__inv_2 _11192_ (.A(net529),
    .Y(_07848_));
 sky130_fd_sc_hd__buf_6 _11193_ (.A(_03176_),
    .X(_03207_));
 sky130_fd_sc_hd__nor2_2 _11194_ (.A(_03146_),
    .B(_03151_),
    .Y(_03208_));
 sky130_fd_sc_hd__buf_8 _11195_ (.A(net591),
    .X(_03209_));
 sky130_fd_sc_hd__nor2b_4 _11196_ (.A(_03209_),
    .B_N(_03147_),
    .Y(_03210_));
 sky130_fd_sc_hd__a22oi_1 _11197_ (.A1(\samples_imag[3][1] ),
    .A2(_03208_),
    .B1(_03210_),
    .B2(\samples_imag[6][1] ),
    .Y(_03211_));
 sky130_fd_sc_hd__nor2_1 _11198_ (.A(_03201_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__buf_12 _11199_ (.A(_03209_),
    .X(_03213_));
 sky130_fd_sc_hd__inv_1 _11200_ (.A(\samples_imag[1][1] ),
    .Y(_03214_));
 sky130_fd_sc_hd__a21oi_4 _11201_ (.A1(_03213_),
    .A2(_03214_),
    .B1(_03169_),
    .Y(_03215_));
 sky130_fd_sc_hd__a21oi_1 _11202_ (.A1(_03158_),
    .A2(\samples_imag[4][1] ),
    .B1(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__mux2_4 _11203_ (.A0(\samples_imag[5][1] ),
    .A1(\samples_imag[7][1] ),
    .S(_03165_),
    .X(_03217_));
 sky130_fd_sc_hd__a32oi_2 _11204_ (.A1(_03185_),
    .A2(_03213_),
    .A3(_03217_),
    .B1(net534),
    .B2(\samples_imag[2][1] ),
    .Y(_03218_));
 sky130_fd_sc_hd__o21ai_1 _11205_ (.A1(_03166_),
    .A2(_03216_),
    .B1(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__o22a_2 _11206_ (.A1(\samples_imag[0][1] ),
    .A2(_03207_),
    .B1(_03212_),
    .B2(_03219_),
    .X(_05902_));
 sky130_fd_sc_hd__inv_2 _11207_ (.A(_05902_),
    .Y(_05898_));
 sky130_fd_sc_hd__inv_6 _11208_ (.A(\temp_imag[0] ),
    .Y(_05897_));
 sky130_fd_sc_hd__inv_2 _11209_ (.A(_05906_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand3_1 _11210_ (.A(_00562_),
    .B(\stage[0] ),
    .C(\stage[1] ),
    .Y(_03220_));
 sky130_fd_sc_hd__and3_1 _11211_ (.A(\group[0] ),
    .B(_02900_),
    .C(_03220_),
    .X(_07913_));
 sky130_fd_sc_hd__and3_1 _11212_ (.A(\group[1] ),
    .B(_02900_),
    .C(_03220_),
    .X(_07915_));
 sky130_fd_sc_hd__and4b_1 _11213_ (.A_N(_07820_),
    .B(_03220_),
    .C(\group[0] ),
    .D(_07807_),
    .X(_07918_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(\group[0] ),
    .B(_07813_),
    .Y(_03221_));
 sky130_fd_sc_hd__nand2_1 _11215_ (.A(\group[1] ),
    .B(_07807_),
    .Y(_03222_));
 sky130_fd_sc_hd__xnor2_1 _11216_ (.A(_03221_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hd__nor2_1 _11217_ (.A(_07820_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(\group[2] ),
    .B(_02900_),
    .Y(_03225_));
 sky130_fd_sc_hd__xnor2_1 _11219_ (.A(_03224_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_03220_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__xor2_1 _11221_ (.A(_07919_),
    .B(_07921_),
    .X(_03228_));
 sky130_fd_sc_hd__xnor2_1 _11222_ (.A(\butterfly_in_group[2] ),
    .B(_07916_),
    .Y(_03229_));
 sky130_fd_sc_hd__xnor2_1 _11223_ (.A(_03228_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__xnor2_1 _11224_ (.A(_03227_),
    .B(_03230_),
    .Y(_00013_));
 sky130_fd_sc_hd__xnor2_1 _11225_ (.A(_05909_),
    .B(_07710_),
    .Y(_03231_));
 sky130_fd_sc_hd__xnor2_1 _11226_ (.A(_00013_),
    .B(_03231_),
    .Y(_00015_));
 sky130_fd_sc_hd__clkbuf_2 clone41 (.A(net474),
    .X(net41));
 sky130_fd_sc_hd__buf_6 _11228_ (.A(net443),
    .X(_03233_));
 sky130_fd_sc_hd__buf_6 _11229_ (.A(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__buf_6 _11230_ (.A(\idx2[0] ),
    .X(_03235_));
 sky130_fd_sc_hd__buf_12 _11231_ (.A(_03235_),
    .X(_03236_));
 sky130_fd_sc_hd__buf_8 _11232_ (.A(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__buf_12 _11233_ (.A(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__mux4_1 _11234_ (.A0(\samples_real[0][12] ),
    .A1(\samples_real[4][12] ),
    .A2(\samples_real[1][12] ),
    .A3(\samples_real[5][12] ),
    .S0(_03234_),
    .S1(net451),
    .X(_03239_));
 sky130_fd_sc_hd__buf_6 _11235_ (.A(_03234_),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_1 _11236_ (.A0(\samples_real[2][12] ),
    .A1(\samples_real[3][12] ),
    .A2(\samples_real[6][12] ),
    .A3(\samples_real[7][12] ),
    .S0(net452),
    .S1(net50),
    .X(_03241_));
 sky130_fd_sc_hd__buf_6 _11237_ (.A(\idx2[1] ),
    .X(_03242_));
 sky130_fd_sc_hd__buf_8 _11238_ (.A(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__buf_4 _11239_ (.A(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__buf_6 _11240_ (.A(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2i_4 _11241_ (.A0(_03239_),
    .A1(_03241_),
    .S(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__buf_4 _11242_ (.A(_00010_),
    .X(_03247_));
 sky130_fd_sc_hd__nand2b_1 _11243_ (.A_N(_03246_),
    .B(_03247_),
    .Y(_05947_));
 sky130_fd_sc_hd__clkinv_8 _11244_ (.A(_00008_),
    .Y(_03248_));
 sky130_fd_sc_hd__clkinv_4 _11245_ (.A(net444),
    .Y(_03249_));
 sky130_fd_sc_hd__nor2_2 _11246_ (.A(_03243_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2b_4 _11247_ (.A(net42),
    .B_N(net46),
    .Y(_03251_));
 sky130_fd_sc_hd__a22o_1 _11248_ (.A1(\samples_imag[5][12] ),
    .A2(_03250_),
    .B1(_03251_),
    .B2(\samples_imag[3][12] ),
    .X(_03252_));
 sky130_fd_sc_hd__inv_1 _11249_ (.A(\samples_imag[4][12] ),
    .Y(_03253_));
 sky130_fd_sc_hd__a21oi_1 _11250_ (.A1(net42),
    .A2(_03253_),
    .B1(net452),
    .Y(_03254_));
 sky130_fd_sc_hd__a21oi_1 _11251_ (.A1(_03249_),
    .A2(\samples_imag[1][12] ),
    .B1(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_4 _11252_ (.A(_03243_),
    .B(net51),
    .Y(_03256_));
 sky130_fd_sc_hd__mux2i_2 _11253_ (.A0(\samples_imag[6][12] ),
    .A1(\samples_imag[7][12] ),
    .S(net452),
    .Y(_03257_));
 sky130_fd_sc_hd__nor2_4 _11254_ (.A(_03235_),
    .B(_03233_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_1 _11255_ (.A(\samples_imag[2][12] ),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__o221ai_4 _11256_ (.A1(_03243_),
    .A2(_03255_),
    .B1(_03256_),
    .B2(_03257_),
    .C1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__a21oi_4 _11257_ (.A1(net451),
    .A2(_03252_),
    .B1(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__or3_4 _11258_ (.A(net493),
    .B(_03235_),
    .C(net443),
    .X(_03262_));
 sky130_fd_sc_hd__buf_6 _11259_ (.A(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__nor2_2 _11260_ (.A(\samples_imag[0][12] ),
    .B(net49),
    .Y(_03264_));
 sky130_fd_sc_hd__nor3_2 _11261_ (.A(_03248_),
    .B(_03261_),
    .C(_03264_),
    .Y(_07938_));
 sky130_fd_sc_hd__buf_8 _11262_ (.A(_03263_),
    .X(_03265_));
 sky130_fd_sc_hd__and3_4 _11263_ (.A(_03242_),
    .B(_03235_),
    .C(_03233_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_4 clone49 (.A(_03262_),
    .X(net49));
 sky130_fd_sc_hd__buf_8 _11265_ (.A(_03266_),
    .X(_03268_));
 sky130_fd_sc_hd__nand2b_4 _11266_ (.A_N(net507),
    .B(net443),
    .Y(_03269_));
 sky130_fd_sc_hd__buf_6 clone51 (.A(_03233_),
    .X(net51));
 sky130_fd_sc_hd__nor2_8 _11268_ (.A(net441),
    .B(net509),
    .Y(_03271_));
 sky130_fd_sc_hd__buf_8 _11269_ (.A(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__a22oi_1 _11270_ (.A1(\samples_real[7][11] ),
    .A2(_03268_),
    .B1(_03272_),
    .B2(\samples_real[4][11] ),
    .Y(_03273_));
 sky130_fd_sc_hd__and2_4 _11271_ (.A(_03242_),
    .B(_03258_),
    .X(_03274_));
 sky130_fd_sc_hd__buf_4 _11272_ (.A(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__nor2_4 _11273_ (.A(_03242_),
    .B(_03233_),
    .Y(_03276_));
 sky130_fd_sc_hd__and2_4 _11274_ (.A(_03276_),
    .B(_03236_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_2 clone43 (.A(_03236_),
    .X(net43));
 sky130_fd_sc_hd__buf_12 _11276_ (.A(_03277_),
    .X(_03279_));
 sky130_fd_sc_hd__a22oi_1 _11277_ (.A1(\samples_real[2][11] ),
    .A2(_03275_),
    .B1(_03279_),
    .B2(\samples_real[1][11] ),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_03273_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__buf_8 _11279_ (.A(_03243_),
    .X(_03282_));
 sky130_fd_sc_hd__buf_12 _11280_ (.A(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__nor2_2 _11281_ (.A(net41),
    .B(_03249_),
    .Y(_03284_));
 sky130_fd_sc_hd__buf_6 _11282_ (.A(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__nor2b_4 _11283_ (.A(net42),
    .B_N(net41),
    .Y(_03286_));
 sky130_fd_sc_hd__clkbuf_8 _11284_ (.A(net510),
    .X(_03287_));
 sky130_fd_sc_hd__a22oi_1 _11285_ (.A1(\samples_real[6][11] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_real[3][11] ),
    .Y(_03288_));
 sky130_fd_sc_hd__and2_2 _11286_ (.A(_03235_),
    .B(_03233_),
    .X(_03289_));
 sky130_fd_sc_hd__buf_6 clone50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_4 _11288_ (.A(_03289_),
    .X(_03291_));
 sky130_fd_sc_hd__buf_4 _11289_ (.A(_03258_),
    .X(_03292_));
 sky130_fd_sc_hd__a211oi_1 _11290_ (.A1(\samples_real[5][11] ),
    .A2(_03291_),
    .B1(_03292_),
    .C1(_03283_),
    .Y(_03293_));
 sky130_fd_sc_hd__a21oi_1 _11291_ (.A1(_03283_),
    .A2(_03288_),
    .B1(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__o22a_4 _11292_ (.A1(\samples_real[0][11] ),
    .A2(_03265_),
    .B1(_03281_),
    .B2(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__nand2_2 _11293_ (.A(_03247_),
    .B(_03295_),
    .Y(_05911_));
 sky130_fd_sc_hd__buf_12 _11294_ (.A(_03283_),
    .X(_03296_));
 sky130_fd_sc_hd__buf_12 _11295_ (.A(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__a22o_1 _11296_ (.A1(\samples_imag[6][11] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_imag[3][11] ),
    .X(_03298_));
 sky130_fd_sc_hd__buf_12 _11297_ (.A(_03238_),
    .X(_03299_));
 sky130_fd_sc_hd__buf_12 _11298_ (.A(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2i_1 _11299_ (.A0(\samples_imag[4][11] ),
    .A1(\samples_imag[5][11] ),
    .S(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand3_1 _11300_ (.A(_03296_),
    .B(net44),
    .C(\samples_imag[7][11] ),
    .Y(_03302_));
 sky130_fd_sc_hd__o21ai_1 _11301_ (.A1(_03296_),
    .A2(_03301_),
    .B1(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__buf_6 _11302_ (.A(_03240_),
    .X(_03304_));
 sky130_fd_sc_hd__inv_1 _11303_ (.A(\samples_imag[1][11] ),
    .Y(_03305_));
 sky130_fd_sc_hd__nand2b_1 _11304_ (.A_N(_03300_),
    .B(\samples_imag[2][11] ),
    .Y(_03306_));
 sky130_fd_sc_hd__a221oi_2 _11305_ (.A1(_03300_),
    .A2(_03305_),
    .B1(_03296_),
    .B2(_03306_),
    .C1(_03304_),
    .Y(_03307_));
 sky130_fd_sc_hd__a221oi_4 _11306_ (.A1(_03297_),
    .A2(_03298_),
    .B1(_03304_),
    .B2(_03303_),
    .C1(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__buf_6 _11307_ (.A(_03265_),
    .X(_03309_));
 sky130_fd_sc_hd__buf_6 _11308_ (.A(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_2 _11309_ (.A(\samples_imag[0][11] ),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__nor3_4 _11310_ (.A(_03248_),
    .B(net497),
    .C(_03311_),
    .Y(_05912_));
 sky130_fd_sc_hd__clkbuf_4 _11311_ (.A(_00008_),
    .X(_03312_));
 sky130_fd_sc_hd__buf_6 _11312_ (.A(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__buf_6 _11313_ (.A(_03309_),
    .X(_03314_));
 sky130_fd_sc_hd__buf_4 _11314_ (.A(_03249_),
    .X(_03315_));
 sky130_fd_sc_hd__and2_2 _11315_ (.A(_03243_),
    .B(net42),
    .X(_03316_));
 sky130_fd_sc_hd__a22oi_2 _11316_ (.A1(_03315_),
    .A2(\samples_imag[2][10] ),
    .B1(_03316_),
    .B2(\samples_imag[6][10] ),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _11317_ (.A1(\samples_imag[5][10] ),
    .A2(_03291_),
    .B1(_03292_),
    .Y(_03318_));
 sky130_fd_sc_hd__and2_4 _11318_ (.A(_03286_),
    .B(net46),
    .X(_03319_));
 sky130_fd_sc_hd__buf_2 clone46 (.A(net493),
    .X(net46));
 sky130_fd_sc_hd__a22o_4 _11320_ (.A1(\samples_imag[1][10] ),
    .A2(_03279_),
    .B1(_03319_),
    .B2(\samples_imag[3][10] ),
    .X(_03321_));
 sky130_fd_sc_hd__a221oi_4 _11321_ (.A1(\samples_imag[7][10] ),
    .A2(_03268_),
    .B1(_03272_),
    .B2(\samples_imag[4][10] ),
    .C1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__o221ai_4 _11322_ (.A1(net44),
    .A2(_03317_),
    .B1(_03318_),
    .B2(_03297_),
    .C1(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__o21ai_4 _11323_ (.A1(_03314_),
    .A2(\samples_imag[0][10] ),
    .B1(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__inv_2 _11324_ (.A(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__nand2_1 _11325_ (.A(_03313_),
    .B(net508),
    .Y(_05921_));
 sky130_fd_sc_hd__inv_1 _11326_ (.A(_05921_),
    .Y(_05913_));
 sky130_fd_sc_hd__a22oi_2 _11327_ (.A1(\samples_imag[7][9] ),
    .A2(_03266_),
    .B1(_03272_),
    .B2(\samples_imag[4][9] ),
    .Y(_03326_));
 sky130_fd_sc_hd__a22oi_1 _11328_ (.A1(\samples_imag[2][9] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\samples_imag[1][9] ),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_03326_),
    .B(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__a22oi_1 _11330_ (.A1(\samples_imag[6][9] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_imag[3][9] ),
    .Y(_03329_));
 sky130_fd_sc_hd__a211oi_1 _11331_ (.A1(\samples_imag[5][9] ),
    .A2(_03289_),
    .B1(_03292_),
    .C1(_03282_),
    .Y(_03330_));
 sky130_fd_sc_hd__a21oi_1 _11332_ (.A1(_03245_),
    .A2(_03329_),
    .B1(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__o22a_4 _11333_ (.A1(\samples_imag[0][9] ),
    .A2(net49),
    .B1(_03328_),
    .B2(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__nand2_2 _11334_ (.A(_00008_),
    .B(_03332_),
    .Y(_05922_));
 sky130_fd_sc_hd__inv_1 _11335_ (.A(_05922_),
    .Y(_05937_));
 sky130_fd_sc_hd__clkbuf_8 _11336_ (.A(_03247_),
    .X(_03333_));
 sky130_fd_sc_hd__nor2_2 _11337_ (.A(\samples_real[0][10] ),
    .B(_03265_),
    .Y(_03334_));
 sky130_fd_sc_hd__buf_4 _11338_ (.A(_03237_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2i_1 _11339_ (.A0(\samples_real[2][10] ),
    .A1(\samples_real[6][10] ),
    .S(_03240_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(\samples_real[7][10] ),
    .B(_03289_),
    .Y(_03337_));
 sky130_fd_sc_hd__o21ai_1 _11341_ (.A1(_03335_),
    .A2(_03336_),
    .B1(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__mux2i_1 _11342_ (.A0(\samples_real[1][10] ),
    .A1(\samples_real[5][10] ),
    .S(_03240_),
    .Y(_03339_));
 sky130_fd_sc_hd__nor2_1 _11343_ (.A(\samples_real[4][10] ),
    .B(net476),
    .Y(_03340_));
 sky130_fd_sc_hd__a211oi_2 _11344_ (.A1(net45),
    .A2(_03339_),
    .B1(_03340_),
    .C1(_03245_),
    .Y(_03341_));
 sky130_fd_sc_hd__a221oi_4 _11345_ (.A1(\samples_real[3][10] ),
    .A2(net465),
    .B1(_03245_),
    .B2(_03338_),
    .C1(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nor2_1 _11346_ (.A(_03334_),
    .B(net462),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_03333_),
    .B(_03343_),
    .Y(_05994_));
 sky130_fd_sc_hd__inv_1 _11348_ (.A(_05994_),
    .Y(_05923_));
 sky130_fd_sc_hd__nor2_2 _11349_ (.A(\samples_imag[0][8] ),
    .B(_03265_),
    .Y(_03344_));
 sky130_fd_sc_hd__nor2b_2 _11350_ (.A(_03243_),
    .B_N(_03289_),
    .Y(_03345_));
 sky130_fd_sc_hd__clkbuf_4 _11351_ (.A(_03345_),
    .X(_03346_));
 sky130_fd_sc_hd__inv_1 _11352_ (.A(\samples_imag[2][8] ),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_1 _11353_ (.A1(_03282_),
    .A2(_03347_),
    .B1(_03335_),
    .Y(_03348_));
 sky130_fd_sc_hd__a31oi_1 _11354_ (.A1(_03282_),
    .A2(_03335_),
    .A3(\samples_imag[3][8] ),
    .B1(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(\samples_imag[6][8] ),
    .A1(\samples_imag[7][8] ),
    .S(_03236_),
    .X(_03350_));
 sky130_fd_sc_hd__nor2_2 _11356_ (.A(_03243_),
    .B(_03237_),
    .Y(_03351_));
 sky130_fd_sc_hd__a221oi_1 _11357_ (.A1(_03282_),
    .A2(_03350_),
    .B1(_03351_),
    .B2(\samples_imag[4][8] ),
    .C1(_03315_),
    .Y(_03352_));
 sky130_fd_sc_hd__a21oi_2 _11358_ (.A1(_03315_),
    .A2(_03349_),
    .B1(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__a221oi_4 _11359_ (.A1(\samples_imag[1][8] ),
    .A2(_03279_),
    .B1(_03346_),
    .B2(\samples_imag[5][8] ),
    .C1(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nor3_4 _11360_ (.A(_03248_),
    .B(_03344_),
    .C(net481),
    .Y(_05938_));
 sky130_fd_sc_hd__a22o_1 _11361_ (.A1(\samples_imag[6][7] ),
    .A2(_03285_),
    .B1(net510),
    .B2(\samples_imag[3][7] ),
    .X(_03355_));
 sky130_fd_sc_hd__mux2i_1 _11362_ (.A0(\samples_imag[4][7] ),
    .A1(\samples_imag[5][7] ),
    .S(_03237_),
    .Y(_03356_));
 sky130_fd_sc_hd__nand3_1 _11363_ (.A(_03244_),
    .B(net469),
    .C(\samples_imag[7][7] ),
    .Y(_03357_));
 sky130_fd_sc_hd__o21ai_2 _11364_ (.A1(_03244_),
    .A2(_03356_),
    .B1(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__inv_1 _11365_ (.A(\samples_imag[1][7] ),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2b_1 _11366_ (.A_N(net452),
    .B(\samples_imag[2][7] ),
    .Y(_03360_));
 sky130_fd_sc_hd__a221oi_2 _11367_ (.A1(net469),
    .A2(_03359_),
    .B1(_03360_),
    .B2(_03244_),
    .C1(net50),
    .Y(_03361_));
 sky130_fd_sc_hd__a221oi_4 _11368_ (.A1(_03355_),
    .A2(_03282_),
    .B1(_03358_),
    .B2(net50),
    .C1(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__nor2_1 _11369_ (.A(\samples_imag[0][7] ),
    .B(_03263_),
    .Y(_03363_));
 sky130_fd_sc_hd__nor2_4 _11370_ (.A(net438),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand2_2 _11371_ (.A(_03312_),
    .B(_03364_),
    .Y(_06069_));
 sky130_fd_sc_hd__inv_1 _11372_ (.A(_06069_),
    .Y(_05980_));
 sky130_fd_sc_hd__a22oi_2 _11373_ (.A1(\samples_imag[7][6] ),
    .A2(_03268_),
    .B1(_03272_),
    .B2(\samples_imag[4][6] ),
    .Y(_03365_));
 sky130_fd_sc_hd__a22oi_1 _11374_ (.A1(\samples_imag[2][6] ),
    .A2(_03275_),
    .B1(_03279_),
    .B2(\samples_imag[1][6] ),
    .Y(_03366_));
 sky130_fd_sc_hd__nand2_1 _11375_ (.A(_03365_),
    .B(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__a22oi_1 _11376_ (.A1(\samples_imag[6][6] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_imag[3][6] ),
    .Y(_03368_));
 sky130_fd_sc_hd__a211oi_2 _11377_ (.A1(\samples_imag[5][6] ),
    .A2(_03291_),
    .B1(_03292_),
    .C1(_03296_),
    .Y(_03369_));
 sky130_fd_sc_hd__a21oi_2 _11378_ (.A1(_03297_),
    .A2(_03368_),
    .B1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o22a_4 _11379_ (.A1(_03309_),
    .A2(\samples_imag[0][6] ),
    .B1(_03367_),
    .B2(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__nand2_2 _11380_ (.A(_03313_),
    .B(_03371_),
    .Y(_06070_));
 sky130_fd_sc_hd__clkinvlp_4 _11381_ (.A(_06070_),
    .Y(_06123_));
 sky130_fd_sc_hd__a22oi_2 _11382_ (.A1(\samples_imag[7][4] ),
    .A2(_03266_),
    .B1(_03272_),
    .B2(\samples_imag[4][4] ),
    .Y(_03372_));
 sky130_fd_sc_hd__a22oi_1 _11383_ (.A1(\samples_imag[2][4] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\samples_imag[1][4] ),
    .Y(_03373_));
 sky130_fd_sc_hd__nand2_1 _11384_ (.A(_03372_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__a22oi_1 _11385_ (.A1(\samples_imag[6][4] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_imag[3][4] ),
    .Y(_03375_));
 sky130_fd_sc_hd__a211oi_1 _11386_ (.A1(\samples_imag[5][4] ),
    .A2(_03289_),
    .B1(_03292_),
    .C1(_03282_),
    .Y(_03376_));
 sky130_fd_sc_hd__a21oi_1 _11387_ (.A1(_03245_),
    .A2(_03375_),
    .B1(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__o22a_4 _11388_ (.A1(\samples_imag[0][4] ),
    .A2(_03265_),
    .B1(_03374_),
    .B2(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__nand2_2 _11389_ (.A(_03312_),
    .B(net483),
    .Y(_07955_));
 sky130_fd_sc_hd__inv_4 _11390_ (.A(_07955_),
    .Y(_06175_));
 sky130_fd_sc_hd__nor2_1 _11391_ (.A(\samples_real[0][9] ),
    .B(_03263_),
    .Y(_03379_));
 sky130_fd_sc_hd__inv_1 _11392_ (.A(\samples_real[2][9] ),
    .Y(_03380_));
 sky130_fd_sc_hd__a21oi_1 _11393_ (.A1(_03243_),
    .A2(_03380_),
    .B1(net43),
    .Y(_03381_));
 sky130_fd_sc_hd__a31oi_1 _11394_ (.A1(_03244_),
    .A2(net43),
    .A3(\samples_real[3][9] ),
    .B1(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(\samples_real[6][9] ),
    .A1(\samples_real[7][9] ),
    .S(_03236_),
    .X(_03383_));
 sky130_fd_sc_hd__a221oi_1 _11396_ (.A1(\samples_real[4][9] ),
    .A2(_03351_),
    .B1(_03383_),
    .B2(_03243_),
    .C1(_03315_),
    .Y(_03384_));
 sky130_fd_sc_hd__a21oi_1 _11397_ (.A1(_03315_),
    .A2(_03382_),
    .B1(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__a221oi_4 _11398_ (.A1(\samples_real[1][9] ),
    .A2(net506),
    .B1(_03345_),
    .B2(\samples_real[5][9] ),
    .C1(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nor2_2 _11399_ (.A(_03379_),
    .B(net504),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_2 _11400_ (.A(_00010_),
    .B(_03387_),
    .Y(_05939_));
 sky130_fd_sc_hd__a22oi_2 _11401_ (.A1(_03249_),
    .A2(\samples_imag[1][5] ),
    .B1(_03289_),
    .B2(\samples_imag[5][5] ),
    .Y(_03388_));
 sky130_fd_sc_hd__a21oi_1 _11402_ (.A1(\samples_imag[6][5] ),
    .A2(_03316_),
    .B1(_03276_),
    .Y(_03389_));
 sky130_fd_sc_hd__a22o_1 _11403_ (.A1(_03271_),
    .A2(\samples_imag[4][5] ),
    .B1(_03274_),
    .B2(\samples_imag[2][5] ),
    .X(_03390_));
 sky130_fd_sc_hd__a221oi_4 _11404_ (.A1(\samples_imag[7][5] ),
    .A2(_03266_),
    .B1(_03319_),
    .B2(\samples_imag[3][5] ),
    .C1(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__o221ai_4 _11405_ (.A1(_03244_),
    .A2(_03388_),
    .B1(_03389_),
    .B2(net451),
    .C1(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__o21ai_4 _11406_ (.A1(\samples_imag[0][5] ),
    .A2(_03263_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_4 _11407_ (.A(_03248_),
    .B(net502),
    .Y(_06124_));
 sky130_fd_sc_hd__mux2i_1 _11408_ (.A0(\samples_imag[6][3] ),
    .A1(\samples_imag[7][3] ),
    .S(_03335_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(\samples_imag[1][3] ),
    .B(_03277_),
    .Y(_03395_));
 sky130_fd_sc_hd__o21ai_1 _11410_ (.A1(_03256_),
    .A2(_03394_),
    .B1(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__a22oi_1 _11411_ (.A1(\samples_imag[5][3] ),
    .A2(_03250_),
    .B1(_03251_),
    .B2(\samples_imag[3][3] ),
    .Y(_03397_));
 sky130_fd_sc_hd__inv_1 _11412_ (.A(\samples_imag[4][3] ),
    .Y(_03398_));
 sky130_fd_sc_hd__a21oi_1 _11413_ (.A1(_03240_),
    .A2(_03398_),
    .B1(_03244_),
    .Y(_03399_));
 sky130_fd_sc_hd__a211oi_1 _11414_ (.A1(_03315_),
    .A2(\samples_imag[2][3] ),
    .B1(_03399_),
    .C1(_03335_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21oi_1 _11415_ (.A1(_03299_),
    .A2(_03397_),
    .B1(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__o22a_4 _11416_ (.A1(\samples_imag[0][3] ),
    .A2(_03265_),
    .B1(_03396_),
    .B2(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_2 _11417_ (.A(_03313_),
    .B(_03402_),
    .Y(_06285_));
 sky130_fd_sc_hd__clkinv_4 _11418_ (.A(_06285_),
    .Y(_06235_));
 sky130_fd_sc_hd__mux4_1 _11419_ (.A0(\samples_imag[2][2] ),
    .A1(\samples_imag[3][2] ),
    .A2(\samples_imag[6][2] ),
    .A3(\samples_imag[7][2] ),
    .S0(_03236_),
    .S1(_03234_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2i_1 _11420_ (.A0(\samples_imag[1][2] ),
    .A1(\samples_imag[5][2] ),
    .S(_03234_),
    .Y(_03404_));
 sky130_fd_sc_hd__nor2_1 _11421_ (.A(\samples_imag[4][2] ),
    .B(net458),
    .Y(_03405_));
 sky130_fd_sc_hd__a211oi_2 _11422_ (.A1(_03237_),
    .A2(_03404_),
    .B1(_03405_),
    .C1(_03244_),
    .Y(_03406_));
 sky130_fd_sc_hd__a21oi_4 _11423_ (.A1(_03282_),
    .A2(_03403_),
    .B1(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__nor2_2 _11424_ (.A(\samples_imag[0][2] ),
    .B(_03263_),
    .Y(_03408_));
 sky130_fd_sc_hd__nor2_1 _11425_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_4 _11426_ (.A(_00008_),
    .B(_03409_),
    .Y(_06286_));
 sky130_fd_sc_hd__inv_2 _11427_ (.A(_06286_),
    .Y(_06501_));
 sky130_fd_sc_hd__mux4_1 _11428_ (.A0(\samples_real[0][8] ),
    .A1(\samples_real[4][8] ),
    .A2(\samples_real[1][8] ),
    .A3(\samples_real[5][8] ),
    .S0(_03234_),
    .S1(_03299_),
    .X(_03410_));
 sky130_fd_sc_hd__mux4_1 _11429_ (.A0(\samples_real[2][8] ),
    .A1(\samples_real[3][8] ),
    .A2(\samples_real[6][8] ),
    .A3(\samples_real[7][8] ),
    .S0(_03238_),
    .S1(_03304_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_4 _11430_ (.A0(_03410_),
    .A1(_03411_),
    .S(_03283_),
    .X(_03412_));
 sky130_fd_sc_hd__and2_2 _11431_ (.A(_03247_),
    .B(_03412_),
    .X(_05958_));
 sky130_fd_sc_hd__inv_1 _11432_ (.A(_05958_),
    .Y(_05981_));
 sky130_fd_sc_hd__mux4_1 _11433_ (.A0(\samples_imag[0][1] ),
    .A1(\samples_imag[4][1] ),
    .A2(\samples_imag[1][1] ),
    .A3(\samples_imag[5][1] ),
    .S0(_03240_),
    .S1(_03299_),
    .X(_03413_));
 sky130_fd_sc_hd__mux4_2 _11434_ (.A0(\samples_imag[2][1] ),
    .A1(\samples_imag[3][1] ),
    .A2(\samples_imag[6][1] ),
    .A3(\samples_imag[7][1] ),
    .S0(net469),
    .S1(_03304_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2i_4 _11435_ (.A0(_03413_),
    .A1(_03414_),
    .S(_03283_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2b_4 _11436_ (.A_N(net499),
    .B(_03312_),
    .Y(_06333_));
 sky130_fd_sc_hd__inv_4 _11437_ (.A(_06333_),
    .Y(_07928_));
 sky130_fd_sc_hd__buf_2 _11438_ (.A(_00009_),
    .X(_03416_));
 sky130_fd_sc_hd__a22oi_2 _11439_ (.A1(\samples_real[7][13] ),
    .A2(_03266_),
    .B1(_03271_),
    .B2(\samples_real[4][13] ),
    .Y(_03417_));
 sky130_fd_sc_hd__a22oi_1 _11440_ (.A1(\samples_real[2][13] ),
    .A2(_03274_),
    .B1(net482),
    .B2(\samples_real[1][13] ),
    .Y(_03418_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(_03417_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__a22oi_1 _11442_ (.A1(\samples_real[6][13] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_real[3][13] ),
    .Y(_03420_));
 sky130_fd_sc_hd__a211oi_1 _11443_ (.A1(\samples_real[5][13] ),
    .A2(_03289_),
    .B1(_03258_),
    .C1(_03244_),
    .Y(_03421_));
 sky130_fd_sc_hd__a21oi_1 _11444_ (.A1(_03282_),
    .A2(_03420_),
    .B1(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__o22a_4 _11445_ (.A1(\samples_real[0][13] ),
    .A2(net49),
    .B1(_03419_),
    .B2(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__and2_0 _11446_ (.A(_03416_),
    .B(_03423_),
    .X(_05954_));
 sky130_fd_sc_hd__a22oi_2 _11447_ (.A1(\samples_real[7][7] ),
    .A2(_03266_),
    .B1(_03272_),
    .B2(\samples_real[4][7] ),
    .Y(_03424_));
 sky130_fd_sc_hd__a22oi_1 _11448_ (.A1(\samples_real[2][7] ),
    .A2(_03275_),
    .B1(net482),
    .B2(\samples_real[1][7] ),
    .Y(_03425_));
 sky130_fd_sc_hd__nand2_1 _11449_ (.A(_03424_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__a22oi_1 _11450_ (.A1(\samples_real[6][7] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_real[3][7] ),
    .Y(_03427_));
 sky130_fd_sc_hd__a211oi_1 _11451_ (.A1(\samples_real[5][7] ),
    .A2(_03291_),
    .B1(_03292_),
    .C1(_03245_),
    .Y(_03428_));
 sky130_fd_sc_hd__a21oi_1 _11452_ (.A1(_03283_),
    .A2(_03427_),
    .B1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o22a_4 _11453_ (.A1(\samples_real[0][7] ),
    .A2(_03265_),
    .B1(_03426_),
    .B2(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_4 _11454_ (.A(_00010_),
    .B(_03430_),
    .Y(_05999_));
 sky130_fd_sc_hd__clkinvlp_4 _11455_ (.A(_05999_),
    .Y(_06002_));
 sky130_fd_sc_hd__clkbuf_4 _11456_ (.A(_00012_),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(_03431_),
    .B(_03295_),
    .Y(_05995_));
 sky130_fd_sc_hd__inv_6 _11458_ (.A(_00010_),
    .Y(_03432_));
 sky130_fd_sc_hd__a22oi_1 _11459_ (.A1(_03315_),
    .A2(\samples_real[1][6] ),
    .B1(_03291_),
    .B2(\samples_real[5][6] ),
    .Y(_03433_));
 sky130_fd_sc_hd__nor2_1 _11460_ (.A(_03297_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__a21oi_1 _11461_ (.A1(\samples_real[6][6] ),
    .A2(_03316_),
    .B1(_03276_),
    .Y(_03435_));
 sky130_fd_sc_hd__nor2_1 _11462_ (.A(net44),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__buf_4 _11463_ (.A(_03275_),
    .X(_03437_));
 sky130_fd_sc_hd__a22oi_1 _11464_ (.A1(\samples_real[4][6] ),
    .A2(_03272_),
    .B1(_03437_),
    .B2(\samples_real[2][6] ),
    .Y(_03438_));
 sky130_fd_sc_hd__buf_6 _11465_ (.A(_03319_),
    .X(_03439_));
 sky130_fd_sc_hd__a22oi_1 _11466_ (.A1(\samples_real[7][6] ),
    .A2(_03268_),
    .B1(_03439_),
    .B2(\samples_real[3][6] ),
    .Y(_03440_));
 sky130_fd_sc_hd__nand2_1 _11467_ (.A(_03438_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__o32ai_4 _11468_ (.A1(_03441_),
    .A2(_03436_),
    .A3(_03434_),
    .B1(_03310_),
    .B2(\samples_real[0][6] ),
    .Y(_03442_));
 sky130_fd_sc_hd__nor2_4 _11469_ (.A(_03432_),
    .B(net455),
    .Y(_05962_));
 sky130_fd_sc_hd__inv_1 _11470_ (.A(_05962_),
    .Y(_06125_));
 sky130_fd_sc_hd__buf_2 _11471_ (.A(_00011_),
    .X(_03443_));
 sky130_fd_sc_hd__mux4_2 _11472_ (.A0(\samples_real[2][5] ),
    .A1(\samples_real[3][5] ),
    .A2(\samples_real[6][5] ),
    .A3(\samples_real[7][5] ),
    .S0(_03299_),
    .S1(_03304_),
    .X(_03444_));
 sky130_fd_sc_hd__mux2i_1 _11473_ (.A0(\samples_real[1][5] ),
    .A1(\samples_real[5][5] ),
    .S(_03304_),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _11474_ (.A(\samples_real[4][5] ),
    .B(net477),
    .Y(_03446_));
 sky130_fd_sc_hd__a211oi_2 _11475_ (.A1(net44),
    .A2(_03445_),
    .B1(_03446_),
    .C1(_03297_),
    .Y(_03447_));
 sky130_fd_sc_hd__a21oi_4 _11476_ (.A1(_03444_),
    .A2(_03297_),
    .B1(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__buf_4 _11477_ (.A(_03309_),
    .X(_03449_));
 sky130_fd_sc_hd__nor2_8 _11478_ (.A(_03449_),
    .B(\samples_real[0][5] ),
    .Y(_03450_));
 sky130_fd_sc_hd__nor2_4 _11479_ (.A(_03450_),
    .B(_03448_),
    .Y(_03451_));
 sky130_fd_sc_hd__and2_4 _11480_ (.A(_03443_),
    .B(_03451_),
    .X(_05963_));
 sky130_fd_sc_hd__mux4_1 _11481_ (.A0(\samples_imag[2][0] ),
    .A1(\samples_imag[3][0] ),
    .A2(\samples_imag[6][0] ),
    .A3(\samples_imag[7][0] ),
    .S0(net475),
    .S1(net446),
    .X(_03452_));
 sky130_fd_sc_hd__nand2_1 _11482_ (.A(net46),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__mux2i_1 _11483_ (.A0(\samples_imag[1][0] ),
    .A1(\samples_imag[5][0] ),
    .S(net447),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _11484_ (.A(\samples_imag[4][0] ),
    .B(_03269_),
    .Y(_03455_));
 sky130_fd_sc_hd__a211o_1 _11485_ (.A1(net41),
    .A2(_03454_),
    .B1(_03455_),
    .C1(net494),
    .X(_03456_));
 sky130_fd_sc_hd__nor2_1 _11486_ (.A(\samples_imag[0][0] ),
    .B(_03262_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21oi_4 _11487_ (.A1(_03453_),
    .A2(_03456_),
    .B1(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_4 _11488_ (.A(_00008_),
    .B(_03458_),
    .Y(_06367_));
 sky130_fd_sc_hd__inv_2 _11489_ (.A(_06367_),
    .Y(_06371_));
 sky130_fd_sc_hd__and2_0 _11490_ (.A(_03416_),
    .B(_03295_),
    .X(_06081_));
 sky130_fd_sc_hd__nor3_4 _11491_ (.A(_03432_),
    .B(_03450_),
    .C(_03448_),
    .Y(_06095_));
 sky130_fd_sc_hd__clkinv_2 _11492_ (.A(_06095_),
    .Y(_06004_));
 sky130_fd_sc_hd__mux4_2 _11493_ (.A0(\samples_real[2][4] ),
    .A1(\samples_real[3][4] ),
    .A2(\samples_real[6][4] ),
    .A3(\samples_real[7][4] ),
    .S0(_03300_),
    .S1(_03304_),
    .X(_03459_));
 sky130_fd_sc_hd__mux2i_1 _11494_ (.A0(\samples_real[1][4] ),
    .A1(\samples_real[5][4] ),
    .S(_03304_),
    .Y(_03460_));
 sky130_fd_sc_hd__nor2_1 _11495_ (.A(\samples_real[4][4] ),
    .B(net477),
    .Y(_03461_));
 sky130_fd_sc_hd__a211oi_2 _11496_ (.A1(_03300_),
    .A2(_03460_),
    .B1(_03297_),
    .C1(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__a21oi_4 _11497_ (.A1(_03459_),
    .A2(_03297_),
    .B1(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_2 _11498_ (.A(\samples_real[0][4] ),
    .B(_03310_),
    .Y(_03464_));
 sky130_fd_sc_hd__nor3_4 _11499_ (.A(_03432_),
    .B(net442),
    .C(_03464_),
    .Y(_06041_));
 sky130_fd_sc_hd__inv_2 _11500_ (.A(_06041_),
    .Y(_06017_));
 sky130_fd_sc_hd__clkbuf_4 _11501_ (.A(_03443_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_4 _11502_ (.A(_03309_),
    .X(_03466_));
 sky130_fd_sc_hd__buf_4 _11503_ (.A(_03272_),
    .X(_03467_));
 sky130_fd_sc_hd__a22oi_4 _11504_ (.A1(\samples_real[7][3] ),
    .A2(_03268_),
    .B1(_03467_),
    .B2(\samples_real[4][3] ),
    .Y(_03468_));
 sky130_fd_sc_hd__clkbuf_4 _11505_ (.A(_03279_),
    .X(_03469_));
 sky130_fd_sc_hd__a22oi_1 _11506_ (.A1(\samples_real[2][3] ),
    .A2(_03437_),
    .B1(_03469_),
    .B2(\samples_real[1][3] ),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _11507_ (.A(_03468_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__a22oi_1 _11508_ (.A1(\samples_real[6][3] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_real[3][3] ),
    .Y(_03472_));
 sky130_fd_sc_hd__a211oi_1 _11509_ (.A1(\samples_real[5][3] ),
    .A2(_03291_),
    .B1(_03292_),
    .C1(_03296_),
    .Y(_03473_));
 sky130_fd_sc_hd__a21oi_1 _11510_ (.A1(_03297_),
    .A2(_03472_),
    .B1(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__o22a_4 _11511_ (.A1(_03466_),
    .A2(\samples_real[0][3] ),
    .B1(_03471_),
    .B2(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__nand2_1 _11512_ (.A(_03465_),
    .B(_03475_),
    .Y(_06018_));
 sky130_fd_sc_hd__inv_1 _11513_ (.A(_06018_),
    .Y(_06031_));
 sky130_fd_sc_hd__mux4_2 _11514_ (.A0(\samples_real[2][2] ),
    .A1(\samples_real[3][2] ),
    .A2(\samples_real[6][2] ),
    .A3(\samples_real[7][2] ),
    .S0(net452),
    .S1(net51),
    .X(_03476_));
 sky130_fd_sc_hd__mux2i_1 _11515_ (.A0(\samples_real[1][2] ),
    .A1(\samples_real[5][2] ),
    .S(_03234_),
    .Y(_03477_));
 sky130_fd_sc_hd__nor2_1 _11516_ (.A(\samples_real[4][2] ),
    .B(net476),
    .Y(_03478_));
 sky130_fd_sc_hd__a211oi_1 _11517_ (.A1(_03335_),
    .A2(_03477_),
    .B1(_03478_),
    .C1(_03282_),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_4 _11518_ (.A1(_03245_),
    .A2(_03476_),
    .B1(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__nor2_1 _11519_ (.A(\samples_real[0][2] ),
    .B(net49),
    .Y(_03481_));
 sky130_fd_sc_hd__nor2_2 _11520_ (.A(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand2_2 _11521_ (.A(_03465_),
    .B(_03482_),
    .Y(_06019_));
 sky130_fd_sc_hd__inv_1 _11522_ (.A(_06019_),
    .Y(_06200_));
 sky130_fd_sc_hd__nand2_4 _11523_ (.A(_03333_),
    .B(_03475_),
    .Y(_06027_));
 sky130_fd_sc_hd__clkinv_2 _11524_ (.A(_06027_),
    .Y(_06199_));
 sky130_fd_sc_hd__a22oi_4 _11525_ (.A1(\samples_real[7][1] ),
    .A2(_03268_),
    .B1(_03467_),
    .B2(\samples_real[4][1] ),
    .Y(_03483_));
 sky130_fd_sc_hd__a22oi_1 _11526_ (.A1(\samples_real[2][1] ),
    .A2(_03275_),
    .B1(_03279_),
    .B2(\samples_real[1][1] ),
    .Y(_03484_));
 sky130_fd_sc_hd__nand2_1 _11527_ (.A(_03483_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__a22oi_1 _11528_ (.A1(\samples_real[6][1] ),
    .A2(_03285_),
    .B1(_03287_),
    .B2(\samples_real[3][1] ),
    .Y(_03486_));
 sky130_fd_sc_hd__a211oi_2 _11529_ (.A1(\samples_real[5][1] ),
    .A2(_03291_),
    .B1(_03292_),
    .C1(_03296_),
    .Y(_03487_));
 sky130_fd_sc_hd__a21oi_1 _11530_ (.A1(_03297_),
    .A2(_03486_),
    .B1(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__o22a_4 _11531_ (.A1(\samples_real[0][1] ),
    .A2(_03449_),
    .B1(_03485_),
    .B2(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_03465_),
    .B(_03489_),
    .Y(_06028_));
 sky130_fd_sc_hd__inv_1 _11533_ (.A(_06028_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand2_1 _11534_ (.A(_03333_),
    .B(_03482_),
    .Y(_06046_));
 sky130_fd_sc_hd__inv_2 _11535_ (.A(_06046_),
    .Y(_06033_));
 sky130_fd_sc_hd__mux4_1 _11536_ (.A0(\samples_real[2][0] ),
    .A1(\samples_real[3][0] ),
    .A2(\samples_real[6][0] ),
    .A3(\samples_real[7][0] ),
    .S0(net41),
    .S1(net42),
    .X(_03490_));
 sky130_fd_sc_hd__inv_1 _11537_ (.A(\samples_real[4][0] ),
    .Y(_03491_));
 sky130_fd_sc_hd__mux2i_1 _11538_ (.A0(\samples_real[1][0] ),
    .A1(\samples_real[5][0] ),
    .S(net445),
    .Y(_03492_));
 sky130_fd_sc_hd__a221oi_2 _11539_ (.A1(_03491_),
    .A2(_03284_),
    .B1(_03492_),
    .B2(net41),
    .C1(net46),
    .Y(_03493_));
 sky130_fd_sc_hd__a21oi_4 _11540_ (.A1(net46),
    .A2(_03490_),
    .B1(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__nor2_4 _11541_ (.A(\samples_real[0][0] ),
    .B(_03262_),
    .Y(_03495_));
 sky130_fd_sc_hd__nor2_1 _11542_ (.A(_03494_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(_03465_),
    .B(_03496_),
    .Y(_06047_));
 sky130_fd_sc_hd__inv_1 _11544_ (.A(_06047_),
    .Y(_06201_));
 sky130_fd_sc_hd__nand2_2 _11545_ (.A(_03333_),
    .B(_03489_),
    .Y(_06434_));
 sky130_fd_sc_hd__clkinv_2 _11546_ (.A(_06434_),
    .Y(_06202_));
 sky130_fd_sc_hd__mux4_1 _11547_ (.A0(\samples_imag[0][13] ),
    .A1(\samples_imag[4][13] ),
    .A2(\samples_imag[1][13] ),
    .A3(\samples_imag[5][13] ),
    .S0(net51),
    .S1(net45),
    .X(_03497_));
 sky130_fd_sc_hd__mux4_1 _11548_ (.A0(\samples_imag[2][13] ),
    .A1(\samples_imag[3][13] ),
    .A2(\samples_imag[6][13] ),
    .A3(\samples_imag[7][13] ),
    .S0(net451),
    .S1(_03304_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2i_4 _11549_ (.A0(_03497_),
    .A1(_03498_),
    .S(_03283_),
    .Y(_03499_));
 sky130_fd_sc_hd__nor2_1 _11550_ (.A(_03248_),
    .B(_03499_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_2 _11551_ (.A(_03333_),
    .B(_03496_),
    .Y(_06465_));
 sky130_fd_sc_hd__inv_2 _11552_ (.A(_06465_),
    .Y(_06382_));
 sky130_fd_sc_hd__clkinvlp_4 _11553_ (.A(_00009_),
    .Y(_03500_));
 sky130_fd_sc_hd__buf_4 _11554_ (.A(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__nor3_1 _11555_ (.A(_03501_),
    .B(_03334_),
    .C(net464),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_1 _11556_ (.A(_03431_),
    .B(_03412_),
    .Y(_06183_));
 sky130_fd_sc_hd__and2_0 _11557_ (.A(_03416_),
    .B(_03412_),
    .X(_06244_));
 sky130_fd_sc_hd__and2_0 _11558_ (.A(_03416_),
    .B(_03430_),
    .X(_06294_));
 sky130_fd_sc_hd__nor2_1 _11559_ (.A(_03501_),
    .B(net456),
    .Y(_06341_));
 sky130_fd_sc_hd__nor2_2 _11560_ (.A(_03463_),
    .B(_03464_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(_03431_),
    .B(_03502_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(_03431_),
    .B(_03482_),
    .Y(_06435_));
 sky130_fd_sc_hd__nor3_1 _11563_ (.A(_03501_),
    .B(net468),
    .C(_03464_),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_1 _11564_ (.A(_03431_),
    .B(_03489_),
    .Y(_06466_));
 sky130_fd_sc_hd__and2_0 _11565_ (.A(_03416_),
    .B(_03489_),
    .X(_08082_));
 sky130_fd_sc_hd__inv_2 _11566_ (.A(_00012_),
    .Y(_03503_));
 sky130_fd_sc_hd__buf_4 _11567_ (.A(_03503_),
    .X(_03504_));
 sky130_fd_sc_hd__nor3_1 _11568_ (.A(_03504_),
    .B(_03494_),
    .C(_03495_),
    .Y(_08083_));
 sky130_fd_sc_hd__and2_0 _11569_ (.A(_08069_),
    .B(_07956_),
    .X(_06471_));
 sky130_fd_sc_hd__nor3_4 _11570_ (.A(_03500_),
    .B(_03494_),
    .C(_03495_),
    .Y(_08120_));
 sky130_fd_sc_hd__inv_1 _11571_ (.A(_08108_),
    .Y(_06331_));
 sky130_fd_sc_hd__nor2b_1 _11572_ (.A(_08108_),
    .B_N(_08112_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_2 _11573_ (.A(_08106_),
    .B(_08124_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand3_1 _11574_ (.A(_08126_),
    .B(_08130_),
    .C(_08116_),
    .Y(_03506_));
 sky130_fd_sc_hd__xnor2_1 _11575_ (.A(_08129_),
    .B(_06367_),
    .Y(_03507_));
 sky130_fd_sc_hd__a21o_1 _11576_ (.A1(_08116_),
    .A2(_08123_),
    .B1(_08115_),
    .X(_03508_));
 sky130_fd_sc_hd__a21oi_4 _11577_ (.A1(_03508_),
    .A2(_08106_),
    .B1(_08105_),
    .Y(_03509_));
 sky130_fd_sc_hd__o41ai_4 _11578_ (.A1(_08120_),
    .A2(_03506_),
    .A3(_03505_),
    .A4(_03507_),
    .B1(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__a21o_1 _11579_ (.A1(_08096_),
    .A2(_03510_),
    .B1(_08095_),
    .X(_03511_));
 sky130_fd_sc_hd__a21oi_2 _11580_ (.A1(_08071_),
    .A2(_03511_),
    .B1(_08070_),
    .Y(_03512_));
 sky130_fd_sc_hd__nor2b_1 _11581_ (.A(_03512_),
    .B_N(_08060_),
    .Y(_03513_));
 sky130_fd_sc_hd__o21ai_1 _11582_ (.A1(_03513_),
    .A2(_08059_),
    .B1(_08047_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2b_1 _11583_ (.A_N(_08046_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21oi_2 _11584_ (.A1(_03515_),
    .A2(_08028_),
    .B1(_08027_),
    .Y(_03516_));
 sky130_fd_sc_hd__nor2b_1 _11585_ (.A(_03516_),
    .B_N(_08013_),
    .Y(_03517_));
 sky130_fd_sc_hd__o21ai_1 _11586_ (.A1(_03517_),
    .A2(_08012_),
    .B1(_08003_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2b_1 _11587_ (.A_N(_08002_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__a21oi_4 _11588_ (.A1(_03519_),
    .A2(_07994_),
    .B1(_07993_),
    .Y(_03520_));
 sky130_fd_sc_hd__o21ai_0 _11589_ (.A1(_03494_),
    .A2(_03495_),
    .B1(_00016_),
    .Y(_03521_));
 sky130_fd_sc_hd__nor2b_1 _11590_ (.A(_03458_),
    .B_N(_00017_),
    .Y(_03522_));
 sky130_fd_sc_hd__xnor2_1 _11591_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__mux2i_1 _11592_ (.A0(\samples_real[6][14] ),
    .A1(\samples_real[7][14] ),
    .S(net43),
    .Y(_03524_));
 sky130_fd_sc_hd__nor2_1 _11593_ (.A(_03256_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__a21oi_1 _11594_ (.A1(\samples_real[1][14] ),
    .A2(net482),
    .B1(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__inv_1 _11595_ (.A(\samples_real[2][14] ),
    .Y(_03527_));
 sky130_fd_sc_hd__nor2_1 _11596_ (.A(_03315_),
    .B(\samples_real[4][14] ),
    .Y(_03528_));
 sky130_fd_sc_hd__o22ai_1 _11597_ (.A1(net51),
    .A2(_03527_),
    .B1(_03528_),
    .B2(_03244_),
    .Y(_03529_));
 sky130_fd_sc_hd__a22oi_1 _11598_ (.A1(\samples_real[5][14] ),
    .A2(_03250_),
    .B1(_03251_),
    .B2(\samples_real[3][14] ),
    .Y(_03530_));
 sky130_fd_sc_hd__nand2_1 _11599_ (.A(_03335_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__o21ai_1 _11600_ (.A1(_03335_),
    .A2(_03529_),
    .B1(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__nor2_1 _11601_ (.A(\samples_real[0][14] ),
    .B(net49),
    .Y(_03533_));
 sky130_fd_sc_hd__a21oi_4 _11602_ (.A1(_03526_),
    .A2(_03532_),
    .B1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_00012_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__xor2_1 _11604_ (.A(_07938_),
    .B(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__xnor2_1 _11605_ (.A(_03523_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__xor2_1 _11606_ (.A(_06124_),
    .B(_06286_),
    .X(_03538_));
 sky130_fd_sc_hd__xnor2_1 _11607_ (.A(_05939_),
    .B(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__xnor2_1 _11608_ (.A(_03537_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__xnor2_1 _11609_ (.A(_05911_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__xor2_1 _11610_ (.A(_03246_),
    .B(_03423_),
    .X(_03542_));
 sky130_fd_sc_hd__xnor2_1 _11611_ (.A(_03343_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_1 _11612_ (.A(_03247_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(_03335_),
    .B(\samples_real[5][15] ),
    .Y(_03545_));
 sky130_fd_sc_hd__mux2_1 _11614_ (.A0(\samples_real[6][15] ),
    .A1(\samples_real[7][15] ),
    .S(net43),
    .X(_03546_));
 sky130_fd_sc_hd__nand2_1 _11615_ (.A(_03245_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__o21ai_1 _11616_ (.A1(_03245_),
    .A2(_03545_),
    .B1(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\samples_real[2][15] ),
    .A1(\samples_real[3][15] ),
    .S(net451),
    .X(_03549_));
 sky130_fd_sc_hd__inv_1 _11618_ (.A(\samples_real[4][15] ),
    .Y(_03550_));
 sky130_fd_sc_hd__a21oi_1 _11619_ (.A1(net50),
    .A2(_03550_),
    .B1(_03335_),
    .Y(_03551_));
 sky130_fd_sc_hd__a21oi_1 _11620_ (.A1(_03315_),
    .A2(\samples_real[1][15] ),
    .B1(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__nor2_1 _11621_ (.A(_03245_),
    .B(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__a221oi_4 _11622_ (.A1(_03304_),
    .A2(_03548_),
    .B1(_03549_),
    .B2(_03251_),
    .C1(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__o21ai_0 _11623_ (.A1(\samples_real[0][15] ),
    .A2(_03265_),
    .B1(_00009_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _11624_ (.A(_03554_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__xor2_2 _11625_ (.A(_00016_),
    .B(_00017_),
    .X(_03557_));
 sky130_fd_sc_hd__xnor2_2 _11626_ (.A(_06212_),
    .B(_05992_),
    .Y(_03558_));
 sky130_fd_sc_hd__xnor2_1 _11627_ (.A(_06109_),
    .B(_06155_),
    .Y(_03559_));
 sky130_fd_sc_hd__xnor2_2 _11628_ (.A(_03559_),
    .B(_03558_),
    .Y(_03560_));
 sky130_fd_sc_hd__xnor2_2 _11629_ (.A(_03557_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__xnor2_1 _11630_ (.A(_03556_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__xnor2_1 _11631_ (.A(_05922_),
    .B(_06069_),
    .Y(_03563_));
 sky130_fd_sc_hd__xnor2_1 _11632_ (.A(_03562_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xnor2_1 _11633_ (.A(_03544_),
    .B(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__xnor2_1 _11634_ (.A(_03565_),
    .B(_03541_),
    .Y(_03566_));
 sky130_fd_sc_hd__xnor2_1 _11635_ (.A(_05928_),
    .B(_05950_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _11636_ (.A(_07987_),
    .B(_07924_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_1 _11637_ (.A(_03567_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__xnor2_1 _11638_ (.A(_06020_),
    .B(_06053_),
    .Y(_03570_));
 sky130_fd_sc_hd__xnor2_1 _11639_ (.A(_07929_),
    .B(_06007_),
    .Y(_03571_));
 sky130_fd_sc_hd__xnor2_1 _11640_ (.A(_03570_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__xnor2_1 _11641_ (.A(_03569_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(_07940_),
    .B(_06015_),
    .Y(_03574_));
 sky130_fd_sc_hd__xnor2_1 _11643_ (.A(_07942_),
    .B(_07945_),
    .Y(_03575_));
 sky130_fd_sc_hd__xnor2_1 _11644_ (.A(_03574_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_1 _11645_ (.A(_03573_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__xnor2_1 _11646_ (.A(_05999_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__xnor2_1 _11647_ (.A(_05932_),
    .B(_05959_),
    .Y(_03579_));
 sky130_fd_sc_hd__xnor2_1 _11648_ (.A(_06035_),
    .B(_05919_),
    .Y(_03580_));
 sky130_fd_sc_hd__xnor2_1 _11649_ (.A(_03579_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__xnor2_1 _11650_ (.A(_07932_),
    .B(_07968_),
    .Y(_03582_));
 sky130_fd_sc_hd__xnor2_1 _11651_ (.A(_05914_),
    .B(_07923_),
    .Y(_03583_));
 sky130_fd_sc_hd__xnor2_1 _11652_ (.A(_03582_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__xnor2_1 _11653_ (.A(_03581_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__xor2_1 _11654_ (.A(_06057_),
    .B(_06089_),
    .X(_03586_));
 sky130_fd_sc_hd__xnor2_1 _11655_ (.A(_06025_),
    .B(_06038_),
    .Y(_03587_));
 sky130_fd_sc_hd__xnor2_1 _11656_ (.A(_03586_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__xnor2_1 _11657_ (.A(_05967_),
    .B(_05971_),
    .Y(_03589_));
 sky130_fd_sc_hd__xnor2_1 _11658_ (.A(_06104_),
    .B(_05964_),
    .Y(_03590_));
 sky130_fd_sc_hd__xnor2_1 _11659_ (.A(_03589_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_1 _11660_ (.A(_03588_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__xnor2_1 _11661_ (.A(_03585_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_03443_),
    .B(_03412_),
    .Y(_03594_));
 sky130_fd_sc_hd__xnor2_1 _11663_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__xnor2_1 _11664_ (.A(_03578_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__a22oi_2 _11665_ (.A1(_03315_),
    .A2(\samples_imag[2][14] ),
    .B1(_03316_),
    .B2(\samples_imag[6][14] ),
    .Y(_03597_));
 sky130_fd_sc_hd__a21oi_1 _11666_ (.A1(\samples_imag[5][14] ),
    .A2(_03291_),
    .B1(_03292_),
    .Y(_03598_));
 sky130_fd_sc_hd__a22o_1 _11667_ (.A1(\samples_imag[4][14] ),
    .A2(_03271_),
    .B1(_03319_),
    .B2(\samples_imag[3][14] ),
    .X(_03599_));
 sky130_fd_sc_hd__a221oi_2 _11668_ (.A1(\samples_imag[7][14] ),
    .A2(_03266_),
    .B1(_03279_),
    .B2(\samples_imag[1][14] ),
    .C1(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__o221ai_4 _11669_ (.A1(net45),
    .A2(_03597_),
    .B1(_03598_),
    .B2(_03283_),
    .C1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__o21ai_2 _11670_ (.A1(\samples_imag[0][14] ),
    .A2(_03265_),
    .B1(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__xor2_1 _11671_ (.A(_03499_),
    .B(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__nand2_1 _11672_ (.A(_03312_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__xnor2_1 _11673_ (.A(_03596_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__xnor2_1 _11674_ (.A(_03605_),
    .B(_03566_),
    .Y(_03606_));
 sky130_fd_sc_hd__xnor2_1 _11675_ (.A(_03520_),
    .B(_03606_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand2_2 _11676_ (.A(_03465_),
    .B(_03458_),
    .Y(_06886_));
 sky130_fd_sc_hd__clkinvlp_4 _11677_ (.A(_06886_),
    .Y(_08131_));
 sky130_fd_sc_hd__and2_1 _11678_ (.A(_00008_),
    .B(_03423_),
    .X(_08132_));
 sky130_fd_sc_hd__nor2b_2 _11679_ (.A(net498),
    .B_N(_03443_),
    .Y(_06531_));
 sky130_fd_sc_hd__inv_1 _11680_ (.A(_06531_),
    .Y(_06829_));
 sky130_fd_sc_hd__nor3_4 _11681_ (.A(_03407_),
    .B(_03408_),
    .C(_03432_),
    .Y(_06713_));
 sky130_fd_sc_hd__nor2_8 _11682_ (.A(net440),
    .B(_03432_),
    .Y(_06526_));
 sky130_fd_sc_hd__clkinv_2 _11683_ (.A(_06526_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_2 _11684_ (.A(_03465_),
    .B(_03409_),
    .Y(_06662_));
 sky130_fd_sc_hd__inv_1 _11685_ (.A(_06662_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand2_2 _11686_ (.A(_03443_),
    .B(_03402_),
    .Y(_06598_));
 sky130_fd_sc_hd__inv_1 _11687_ (.A(_06598_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand2_1 _11688_ (.A(_03465_),
    .B(_03378_),
    .Y(_06563_));
 sky130_fd_sc_hd__inv_2 _11689_ (.A(_03393_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_8 _11690_ (.A(_03247_),
    .B(net461),
    .Y(_06564_));
 sky130_fd_sc_hd__inv_1 _11691_ (.A(_06564_),
    .Y(_06775_));
 sky130_fd_sc_hd__and2_1 _11692_ (.A(_03247_),
    .B(_03378_),
    .X(_06535_));
 sky130_fd_sc_hd__inv_2 _11693_ (.A(_06535_),
    .Y(_06599_));
 sky130_fd_sc_hd__and2_4 _11694_ (.A(_03443_),
    .B(_03607_),
    .X(_06536_));
 sky130_fd_sc_hd__inv_1 _11695_ (.A(_06536_),
    .Y(_06607_));
 sky130_fd_sc_hd__nand2_4 _11696_ (.A(_03333_),
    .B(_03371_),
    .Y(_06608_));
 sky130_fd_sc_hd__inv_4 _11697_ (.A(_06608_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2b_2 _11698_ (.A_N(_03246_),
    .B(_03312_),
    .Y(_06643_));
 sky130_fd_sc_hd__inv_1 _11699_ (.A(_06643_),
    .Y(_06646_));
 sky130_fd_sc_hd__and2_0 _11700_ (.A(_03443_),
    .B(_03371_),
    .X(_08137_));
 sky130_fd_sc_hd__inv_1 _11701_ (.A(_08137_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand2_2 _11702_ (.A(_03333_),
    .B(_03364_),
    .Y(_06577_));
 sky130_fd_sc_hd__inv_1 _11703_ (.A(_06577_),
    .Y(_06721_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_03465_),
    .B(_03364_),
    .Y(_06550_));
 sky130_fd_sc_hd__nor2_1 _11705_ (.A(_03344_),
    .B(net479),
    .Y(_03608_));
 sky130_fd_sc_hd__nand2_2 _11706_ (.A(_03333_),
    .B(_03608_),
    .Y(_06551_));
 sky130_fd_sc_hd__inv_1 _11707_ (.A(_06551_),
    .Y(_06722_));
 sky130_fd_sc_hd__nand2_2 _11708_ (.A(_03333_),
    .B(_03332_),
    .Y(_06552_));
 sky130_fd_sc_hd__inv_1 _11709_ (.A(_06552_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_2 _11710_ (.A(_03247_),
    .B(_03325_),
    .Y(_06610_));
 sky130_fd_sc_hd__inv_2 _11711_ (.A(_06610_),
    .Y(_06546_));
 sky130_fd_sc_hd__nor3_4 _11712_ (.A(_03432_),
    .B(_03311_),
    .C(net495),
    .Y(_06547_));
 sky130_fd_sc_hd__nor3_1 _11713_ (.A(_03432_),
    .B(_03261_),
    .C(_03264_),
    .Y(_06555_));
 sky130_fd_sc_hd__nand2_2 _11714_ (.A(_03313_),
    .B(_03295_),
    .Y(_06630_));
 sky130_fd_sc_hd__inv_1 _11715_ (.A(_06630_),
    .Y(_06693_));
 sky130_fd_sc_hd__nor2_1 _11716_ (.A(_03504_),
    .B(_03499_),
    .Y(_08141_));
 sky130_fd_sc_hd__nor2_1 _11717_ (.A(_03501_),
    .B(_03602_),
    .Y(_08142_));
 sky130_fd_sc_hd__nor3_4 _11718_ (.A(_03480_),
    .B(_03248_),
    .C(_03481_),
    .Y(_06729_));
 sky130_fd_sc_hd__and2_4 _11719_ (.A(_03312_),
    .B(_03489_),
    .X(_06778_));
 sky130_fd_sc_hd__nor3_4 _11720_ (.A(net467),
    .B(_03464_),
    .C(_03248_),
    .Y(_08146_));
 sky130_fd_sc_hd__inv_4 _11721_ (.A(net471),
    .Y(_06853_));
 sky130_fd_sc_hd__nor3_4 _11722_ (.A(net463),
    .B(_03334_),
    .C(_03248_),
    .Y(_06631_));
 sky130_fd_sc_hd__nor3_4 _11723_ (.A(_03248_),
    .B(_03494_),
    .C(_03495_),
    .Y(_06833_));
 sky130_fd_sc_hd__nand2_4 _11724_ (.A(_03313_),
    .B(_03475_),
    .Y(_06903_));
 sky130_fd_sc_hd__clkinv_4 _11725_ (.A(_06903_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand2_4 _11726_ (.A(_03313_),
    .B(_03451_),
    .Y(_06797_));
 sky130_fd_sc_hd__inv_2 _11727_ (.A(_06797_),
    .Y(_06986_));
 sky130_fd_sc_hd__and2_2 _11728_ (.A(_03312_),
    .B(_03430_),
    .X(_08156_));
 sky130_fd_sc_hd__inv_2 _11729_ (.A(_08156_),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_4 _11730_ (.A(_03313_),
    .B(_03412_),
    .Y(_06698_));
 sky130_fd_sc_hd__inv_2 _11731_ (.A(_06698_),
    .Y(_06648_));
 sky130_fd_sc_hd__o32a_4 _11732_ (.A1(_03434_),
    .A2(_03436_),
    .A3(_03441_),
    .B1(_03310_),
    .B2(\samples_real[0][6] ),
    .X(_03609_));
 sky130_fd_sc_hd__nand2_4 _11733_ (.A(_03313_),
    .B(_03609_),
    .Y(_06749_));
 sky130_fd_sc_hd__clkinv_2 _11734_ (.A(_06749_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2_2 _11735_ (.A(_03313_),
    .B(_03387_),
    .Y(_06635_));
 sky130_fd_sc_hd__inv_2 _11736_ (.A(_06635_),
    .Y(_06632_));
 sky130_fd_sc_hd__and2_0 _11737_ (.A(_08335_),
    .B(_06833_),
    .X(_08336_));
 sky130_fd_sc_hd__nand4b_1 _11738_ (.A_N(_07103_),
    .B(_08327_),
    .C(_08329_),
    .D(_08331_),
    .Y(_03610_));
 sky130_fd_sc_hd__a21oi_1 _11739_ (.A1(_08338_),
    .A2(_06833_),
    .B1(_08337_),
    .Y(_03611_));
 sky130_fd_sc_hd__nor2_1 _11740_ (.A(_03610_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__and3_1 _11741_ (.A(_08320_),
    .B(_08266_),
    .C(_08296_),
    .X(_03613_));
 sky130_fd_sc_hd__o2111ai_4 _11742_ (.A1(_08326_),
    .A2(_03612_),
    .B1(_03613_),
    .C1(_08284_),
    .D1(_08313_),
    .Y(_03614_));
 sky130_fd_sc_hd__a21oi_1 _11743_ (.A1(_08319_),
    .A2(_08313_),
    .B1(_08312_),
    .Y(_03615_));
 sky130_fd_sc_hd__nor2b_1 _11744_ (.A(_03615_),
    .B_N(_08296_),
    .Y(_03616_));
 sky130_fd_sc_hd__o21ai_1 _11745_ (.A1(_08295_),
    .A2(_03616_),
    .B1(_08284_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2b_1 _11746_ (.A_N(_08283_),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__a21oi_2 _11747_ (.A1(_08266_),
    .A2(_03618_),
    .B1(_08265_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21boi_0 _11748_ (.A1(_03614_),
    .A2(_03619_),
    .B1_N(_08252_),
    .Y(_03620_));
 sky130_fd_sc_hd__o21ai_1 _11749_ (.A1(_08251_),
    .A2(_03620_),
    .B1(_08238_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2b_1 _11750_ (.A_N(_08237_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__a21oi_2 _11751_ (.A1(_03622_),
    .A2(_08223_),
    .B1(_08222_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _11752_ (.A(_03312_),
    .B(_03534_),
    .Y(_03624_));
 sky130_fd_sc_hd__nor2b_1 _11753_ (.A(_03458_),
    .B_N(_00016_),
    .Y(_03625_));
 sky130_fd_sc_hd__xnor2_1 _11754_ (.A(_03624_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__nor2_1 _11755_ (.A(_03503_),
    .B(_03602_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _11756_ (.A(_03443_),
    .B(_03608_),
    .Y(_03628_));
 sky130_fd_sc_hd__xnor2_1 _11757_ (.A(_03627_),
    .B(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__xnor2_1 _11758_ (.A(_03626_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__xor2_1 _11759_ (.A(_08168_),
    .B(_06702_),
    .X(_03631_));
 sky130_fd_sc_hd__xnor2_1 _11760_ (.A(_06691_),
    .B(_06705_),
    .Y(_03632_));
 sky130_fd_sc_hd__xnor2_1 _11761_ (.A(_03631_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__xnor2_1 _11762_ (.A(_08143_),
    .B(_06628_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_1 _11763_ (.A(_08133_),
    .B(_08136_),
    .Y(_03635_));
 sky130_fd_sc_hd__xnor2_1 _11764_ (.A(_03634_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__xnor2_1 _11765_ (.A(_03633_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__xor2_1 _11766_ (.A(_06587_),
    .B(_06619_),
    .X(_03638_));
 sky130_fd_sc_hd__xnor2_1 _11767_ (.A(_06561_),
    .B(_06574_),
    .Y(_03639_));
 sky130_fd_sc_hd__xnor2_1 _11768_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__xnor2_1 _11769_ (.A(_06529_),
    .B(_08139_),
    .Y(_03641_));
 sky130_fd_sc_hd__xnor2_1 _11770_ (.A(_08197_),
    .B(_06549_),
    .Y(_03642_));
 sky130_fd_sc_hd__xnor2_1 _11771_ (.A(_03641_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__xnor2_1 _11772_ (.A(_03640_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__xnor2_1 _11773_ (.A(_03637_),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xor2_1 _11774_ (.A(_06591_),
    .B(_06556_),
    .X(_03646_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(_06553_),
    .B(_06543_),
    .Y(_03647_));
 sky130_fd_sc_hd__xnor2_1 _11776_ (.A(_03646_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__xnor2_1 _11777_ (.A(_08159_),
    .B(_08158_),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_1 _11778_ (.A(_06583_),
    .B(_06651_),
    .Y(_03650_));
 sky130_fd_sc_hd__xnor2_1 _11779_ (.A(_03649_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__xnor2_1 _11780_ (.A(_03648_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__xnor2_1 _11781_ (.A(_06639_),
    .B(_06644_),
    .Y(_03653_));
 sky130_fd_sc_hd__xnor2_1 _11782_ (.A(_08147_),
    .B(_08161_),
    .Y(_03654_));
 sky130_fd_sc_hd__xnor2_1 _11783_ (.A(_03653_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__xnor2_1 _11784_ (.A(_03652_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__xnor2_1 _11785_ (.A(_03645_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__nor2_1 _11786_ (.A(_03261_),
    .B(_03264_),
    .Y(_03658_));
 sky130_fd_sc_hd__xnor2_1 _11787_ (.A(_03658_),
    .B(_03499_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _11788_ (.A(_03247_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__xnor2_1 _11789_ (.A(_03657_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__xnor2_1 _11790_ (.A(_03630_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__xor2_1 _11791_ (.A(_06713_),
    .B(net487),
    .X(_03663_));
 sky130_fd_sc_hd__o21ai_0 _11792_ (.A1(_03494_),
    .A2(_03495_),
    .B1(_00017_),
    .Y(_03664_));
 sky130_fd_sc_hd__xnor2_1 _11793_ (.A(_08132_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__xnor2_1 _11794_ (.A(_03663_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__xor2_1 _11795_ (.A(net485),
    .B(_03402_),
    .X(_03667_));
 sky130_fd_sc_hd__xnor2_1 _11796_ (.A(net500),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand2_1 _11797_ (.A(_03443_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__xnor2_1 _11798_ (.A(_03666_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__xnor2_1 _11799_ (.A(_03246_),
    .B(_03295_),
    .Y(_03671_));
 sky130_fd_sc_hd__nand2_1 _11800_ (.A(_03312_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__mux2i_1 _11801_ (.A0(\samples_imag[1][15] ),
    .A1(\samples_imag[5][15] ),
    .S(net50),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(net45),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__o21ai_1 _11803_ (.A1(\samples_imag[4][15] ),
    .A2(_03269_),
    .B1(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nor2_8 _11804_ (.A(net43),
    .B(_03256_),
    .Y(_03676_));
 sky130_fd_sc_hd__a22o_1 _11805_ (.A1(\samples_imag[7][15] ),
    .A2(_03266_),
    .B1(_03676_),
    .B2(\samples_imag[6][15] ),
    .X(_03677_));
 sky130_fd_sc_hd__a221oi_2 _11806_ (.A1(\samples_imag[2][15] ),
    .A2(_03275_),
    .B1(net465),
    .B2(\samples_imag[3][15] ),
    .C1(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_4 _11807_ (.A1(_03283_),
    .A2(_03675_),
    .B1(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__o211ai_2 _11808_ (.A1(\samples_imag[0][15] ),
    .A2(_03265_),
    .B1(_03679_),
    .C1(_00009_),
    .Y(_03680_));
 sky130_fd_sc_hd__xor2_2 _11809_ (.A(_06538_),
    .B(_06806_),
    .X(_03681_));
 sky130_fd_sc_hd__xnor2_1 _11810_ (.A(_06633_),
    .B(_06758_),
    .Y(_03682_));
 sky130_fd_sc_hd__xnor2_2 _11811_ (.A(_03682_),
    .B(_03681_),
    .Y(_03683_));
 sky130_fd_sc_hd__xnor2_1 _11812_ (.A(_03683_),
    .B(_03557_),
    .Y(_03684_));
 sky130_fd_sc_hd__xnor2_1 _11813_ (.A(_03684_),
    .B(_03680_),
    .Y(_03685_));
 sky130_fd_sc_hd__xnor2_1 _11814_ (.A(_03685_),
    .B(_06564_),
    .Y(_03686_));
 sky130_fd_sc_hd__xnor2_1 _11815_ (.A(_03686_),
    .B(_03672_),
    .Y(_03687_));
 sky130_fd_sc_hd__xnor2_1 _11816_ (.A(_03687_),
    .B(_03670_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_2 _11817_ (.A(_03688_),
    .B(_03662_),
    .Y(_03689_));
 sky130_fd_sc_hd__xor2_1 _11818_ (.A(_03689_),
    .B(_03623_),
    .X(_00019_));
 sky130_fd_sc_hd__nor2b_1 _11819_ (.A(_07819_),
    .B_N(\state[1] ),
    .Y(_00003_));
 sky130_fd_sc_hd__nand2_1 _11820_ (.A(_03465_),
    .B(_03609_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _11821_ (.A(_03465_),
    .B(_03502_),
    .Y(_06005_));
 sky130_fd_sc_hd__inv_1 _11822_ (.A(_07942_),
    .Y(_06099_));
 sky130_fd_sc_hd__inv_1 _11823_ (.A(_08155_),
    .Y(_06636_));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(_06706_),
    .Y(_06755_));
 sky130_fd_sc_hd__inv_1 _11825_ (.A(_08211_),
    .Y(_06840_));
 sky130_fd_sc_hd__inv_1 _11826_ (.A(_08225_),
    .Y(_06895_));
 sky130_fd_sc_hd__inv_1 _11827_ (.A(_06898_),
    .Y(_06905_));
 sky130_fd_sc_hd__inv_1 _11828_ (.A(_06872_),
    .Y(_06914_));
 sky130_fd_sc_hd__inv_1 _11829_ (.A(_06879_),
    .Y(_06922_));
 sky130_fd_sc_hd__inv_1 _11830_ (.A(_06931_),
    .Y(_06933_));
 sky130_fd_sc_hd__inv_1 _11831_ (.A(_08242_),
    .Y(_06938_));
 sky130_fd_sc_hd__inv_1 _11832_ (.A(net488),
    .Y(_06948_));
 sky130_fd_sc_hd__inv_2 _11833_ (.A(_06713_),
    .Y(_06597_));
 sky130_fd_sc_hd__inv_1 _11834_ (.A(_08256_),
    .Y(_06981_));
 sky130_fd_sc_hd__inv_1 _11835_ (.A(_08274_),
    .Y(_07027_));
 sky130_fd_sc_hd__inv_1 _11836_ (.A(_06930_),
    .Y(_06927_));
 sky130_fd_sc_hd__inv_1 _11837_ (.A(_08276_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand2_1 _11838_ (.A(_03431_),
    .B(_03423_),
    .Y(_05948_));
 sky130_fd_sc_hd__inv_1 _11839_ (.A(_07948_),
    .Y(_06051_));
 sky130_fd_sc_hd__inv_1 _11840_ (.A(_07980_),
    .Y(_06252_));
 sky130_fd_sc_hd__inv_1 _11841_ (.A(_07991_),
    .Y(_06302_));
 sky130_fd_sc_hd__inv_1 _11842_ (.A(_06496_),
    .Y(_06493_));
 sky130_fd_sc_hd__inv_1 _11843_ (.A(_06506_),
    .Y(_06502_));
 sky130_fd_sc_hd__inv_1 _11844_ (.A(_08114_),
    .Y(_06522_));
 sky130_fd_sc_hd__inv_1 _11845_ (.A(_08152_),
    .Y(_06658_));
 sky130_fd_sc_hd__inv_1 _11846_ (.A(_08170_),
    .Y(_06689_));
 sky130_fd_sc_hd__inv_1 _11847_ (.A(_08183_),
    .Y(_06742_));
 sky130_fd_sc_hd__inv_1 _11848_ (.A(_08195_),
    .Y(_06790_));
 sky130_fd_sc_hd__inv_1 _11849_ (.A(_08208_),
    .Y(_06846_));
 sky130_fd_sc_hd__inv_1 _11850_ (.A(_08213_),
    .Y(_06877_));
 sky130_fd_sc_hd__inv_1 _11851_ (.A(_06904_),
    .Y(_06944_));
 sky130_fd_sc_hd__inv_1 _11852_ (.A(_06964_),
    .Y(_06961_));
 sky130_fd_sc_hd__inv_1 _11853_ (.A(_08306_),
    .Y(_07070_));
 sky130_fd_sc_hd__inv_1 _11854_ (.A(_07095_),
    .Y(_07092_));
 sky130_fd_sc_hd__inv_1 _11855_ (.A(_08317_),
    .Y(_07097_));
 sky130_fd_sc_hd__inv_1 _11856_ (.A(_07105_),
    .Y(_07100_));
 sky130_fd_sc_hd__inv_2 _11857_ (.A(_07731_),
    .Y(_05884_));
 sky130_fd_sc_hd__inv_2 _11858_ (.A(_07845_),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _11859_ (.A(_03416_),
    .B(_03534_),
    .Y(_05949_));
 sky130_fd_sc_hd__nand2b_1 _11860_ (.A_N(_03246_),
    .B(_00009_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand2_1 _11861_ (.A(_03416_),
    .B(_03387_),
    .Y(_06184_));
 sky130_fd_sc_hd__inv_1 _11862_ (.A(_07979_),
    .Y(_06253_));
 sky130_fd_sc_hd__inv_1 _11863_ (.A(_07990_),
    .Y(_06303_));
 sky130_fd_sc_hd__nand2_1 _11864_ (.A(_03416_),
    .B(_03451_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_1 _11865_ (.A(_03416_),
    .B(_03475_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(_03416_),
    .B(_03482_),
    .Y(_06467_));
 sky130_fd_sc_hd__inv_1 _11867_ (.A(_06484_),
    .Y(_06494_));
 sky130_fd_sc_hd__inv_1 _11868_ (.A(_06507_),
    .Y(_06503_));
 sky130_fd_sc_hd__inv_1 _11869_ (.A(_08163_),
    .Y(_06638_));
 sky130_fd_sc_hd__inv_1 _11870_ (.A(_08151_),
    .Y(_06659_));
 sky130_fd_sc_hd__inv_1 _11871_ (.A(_08169_),
    .Y(_06690_));
 sky130_fd_sc_hd__inv_1 _11872_ (.A(_08182_),
    .Y(_06743_));
 sky130_fd_sc_hd__inv_1 _11873_ (.A(_08194_),
    .Y(_06791_));
 sky130_fd_sc_hd__inv_1 _11874_ (.A(_08216_),
    .Y(_06842_));
 sky130_fd_sc_hd__inv_1 _11875_ (.A(_08207_),
    .Y(_06847_));
 sky130_fd_sc_hd__inv_1 _11876_ (.A(_08212_),
    .Y(_06878_));
 sky130_fd_sc_hd__inv_1 _11877_ (.A(_08231_),
    .Y(_06897_));
 sky130_fd_sc_hd__inv_1 _11878_ (.A(_06899_),
    .Y(_06924_));
 sky130_fd_sc_hd__inv_1 _11879_ (.A(_08247_),
    .Y(_06940_));
 sky130_fd_sc_hd__inv_1 _11880_ (.A(_06949_),
    .Y(_06945_));
 sky130_fd_sc_hd__nand2_4 _11881_ (.A(_03333_),
    .B(_03402_),
    .Y(_06565_));
 sky130_fd_sc_hd__inv_1 _11882_ (.A(_08261_),
    .Y(_06983_));
 sky130_fd_sc_hd__inv_1 _11883_ (.A(_08281_),
    .Y(_07029_));
 sky130_fd_sc_hd__inv_1 _11884_ (.A(_08287_),
    .Y(_07049_));
 sky130_fd_sc_hd__inv_1 _11885_ (.A(_08316_),
    .Y(_07098_));
 sky130_fd_sc_hd__inv_1 _11886_ (.A(_05910_),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_1 _11887_ (.A(_05956_),
    .Y(_07936_));
 sky130_fd_sc_hd__inv_1 _11888_ (.A(_05968_),
    .Y(_05991_));
 sky130_fd_sc_hd__inv_1 _11889_ (.A(_05993_),
    .Y(_06013_));
 sky130_fd_sc_hd__inv_1 _11890_ (.A(_06049_),
    .Y(_06100_));
 sky130_fd_sc_hd__inv_1 _11891_ (.A(_06083_),
    .Y(_07963_));
 sky130_fd_sc_hd__inv_1 _11892_ (.A(_06087_),
    .Y(_06130_));
 sky130_fd_sc_hd__inv_1 _11893_ (.A(_06136_),
    .Y(_07972_));
 sky130_fd_sc_hd__inv_1 _11894_ (.A(_06139_),
    .Y(_06180_));
 sky130_fd_sc_hd__inv_1 _11895_ (.A(_06190_),
    .Y(_06240_));
 sky130_fd_sc_hd__inv_1 _11896_ (.A(_06194_),
    .Y(_06206_));
 sky130_fd_sc_hd__inv_1 _11897_ (.A(_06197_),
    .Y(_06251_));
 sky130_fd_sc_hd__inv_1 _11898_ (.A(_06246_),
    .Y(_07995_));
 sky130_fd_sc_hd__inv_1 _11899_ (.A(_06250_),
    .Y(_06290_));
 sky130_fd_sc_hd__inv_1 _11900_ (.A(_06280_),
    .Y(_08004_));
 sky130_fd_sc_hd__inv_1 _11901_ (.A(_06296_),
    .Y(_08006_));
 sky130_fd_sc_hd__inv_1 _11902_ (.A(_06300_),
    .Y(_06337_));
 sky130_fd_sc_hd__inv_1 _11903_ (.A(_06328_),
    .Y(_08014_));
 sky130_fd_sc_hd__inv_1 _11904_ (.A(_06332_),
    .Y(_08016_));
 sky130_fd_sc_hd__inv_2 _11905_ (.A(_06343_),
    .Y(_08019_));
 sky130_fd_sc_hd__inv_1 _11906_ (.A(_06347_),
    .Y(_06375_));
 sky130_fd_sc_hd__inv_1 _11907_ (.A(_06370_),
    .Y(_08048_));
 sky130_fd_sc_hd__inv_2 _11908_ (.A(_06408_),
    .Y(_08037_));
 sky130_fd_sc_hd__inv_1 _11909_ (.A(_06431_),
    .Y(_08052_));
 sky130_fd_sc_hd__inv_1 _11910_ (.A(_06455_),
    .Y(_08072_));
 sky130_fd_sc_hd__inv_1 _11911_ (.A(_06462_),
    .Y(_08063_));
 sky130_fd_sc_hd__inv_1 _11912_ (.A(_06530_),
    .Y(_08135_));
 sky130_fd_sc_hd__inv_2 _11913_ (.A(_06539_),
    .Y(_06541_));
 sky130_fd_sc_hd__inv_2 _11914_ (.A(_06562_),
    .Y(_06589_));
 sky130_fd_sc_hd__inv_1 _11915_ (.A(_06575_),
    .Y(_06581_));
 sky130_fd_sc_hd__inv_1 _11916_ (.A(_06596_),
    .Y(_06653_));
 sky130_fd_sc_hd__inv_1 _11917_ (.A(_06616_),
    .Y(_06655_));
 sky130_fd_sc_hd__inv_1 _11918_ (.A(_06620_),
    .Y(_06626_));
 sky130_fd_sc_hd__inv_1 _11919_ (.A(_06634_),
    .Y(_06641_));
 sky130_fd_sc_hd__inv_1 _11920_ (.A(_06679_),
    .Y(_06685_));
 sky130_fd_sc_hd__inv_1 _11921_ (.A(_06712_),
    .Y(_06763_));
 sky130_fd_sc_hd__inv_1 _11922_ (.A(_06732_),
    .Y(_06737_));
 sky130_fd_sc_hd__inv_1 _11923_ (.A(_06769_),
    .Y(_06815_));
 sky130_fd_sc_hd__inv_1 _11924_ (.A(_06788_),
    .Y(_06817_));
 sky130_fd_sc_hd__inv_1 _11925_ (.A(_06823_),
    .Y(_06873_));
 sky130_fd_sc_hd__inv_1 _11926_ (.A(_06835_),
    .Y(_06841_));
 sky130_fd_sc_hd__inv_1 _11927_ (.A(_06860_),
    .Y(_06871_));
 sky130_fd_sc_hd__inv_1 _11928_ (.A(_06909_),
    .Y(_06920_));
 sky130_fd_sc_hd__inv_1 _11929_ (.A(_06926_),
    .Y(_06965_));
 sky130_fd_sc_hd__inv_1 _11930_ (.A(_06955_),
    .Y(_06967_));
 sky130_fd_sc_hd__inv_1 _11931_ (.A(_06973_),
    .Y(_07007_));
 sky130_fd_sc_hd__inv_1 _11932_ (.A(_06992_),
    .Y(_07021_));
 sky130_fd_sc_hd__inv_1 _11933_ (.A(_06997_),
    .Y(_07009_));
 sky130_fd_sc_hd__inv_1 _11934_ (.A(_07068_),
    .Y(_07071_));
 sky130_fd_sc_hd__inv_1 _11935_ (.A(_05955_),
    .Y(_07931_));
 sky130_fd_sc_hd__inv_1 _11936_ (.A(_06029_),
    .Y(_06024_));
 sky130_fd_sc_hd__inv_1 _11937_ (.A(_06011_),
    .Y(_06008_));
 sky130_fd_sc_hd__inv_1 _11938_ (.A(_06048_),
    .Y(_06044_));
 sky130_fd_sc_hd__inv_1 _11939_ (.A(_06082_),
    .Y(_07950_));
 sky130_fd_sc_hd__inv_1 _11940_ (.A(_06135_),
    .Y(_07964_));
 sky130_fd_sc_hd__inv_1 _11941_ (.A(_06245_),
    .Y(_07984_));
 sky130_fd_sc_hd__inv_1 _11942_ (.A(_06295_),
    .Y(_07996_));
 sky130_fd_sc_hd__inv_1 _11943_ (.A(_06327_),
    .Y(_08005_));
 sky130_fd_sc_hd__inv_1 _11944_ (.A(_06342_),
    .Y(_08007_));
 sky130_fd_sc_hd__inv_1 _11945_ (.A(_06369_),
    .Y(_08017_));
 sky130_fd_sc_hd__inv_1 _11946_ (.A(_06407_),
    .Y(_08022_));
 sky130_fd_sc_hd__inv_1 _11947_ (.A(_06430_),
    .Y(_08038_));
 sky130_fd_sc_hd__inv_1 _11948_ (.A(_06454_),
    .Y(_08049_));
 sky130_fd_sc_hd__inv_1 _11949_ (.A(_06461_),
    .Y(_08053_));
 sky130_fd_sc_hd__inv_1 _11950_ (.A(_06533_),
    .Y(_06540_));
 sky130_fd_sc_hd__inv_1 _11951_ (.A(_06570_),
    .Y(_06580_));
 sky130_fd_sc_hd__inv_1 _11952_ (.A(_06595_),
    .Y(_06590_));
 sky130_fd_sc_hd__inv_1 _11953_ (.A(_06604_),
    .Y(_06582_));
 sky130_fd_sc_hd__inv_1 _11954_ (.A(_06615_),
    .Y(_06625_));
 sky130_fd_sc_hd__inv_1 _11955_ (.A(_06647_),
    .Y(_06642_));
 sky130_fd_sc_hd__inv_1 _11956_ (.A(_06674_),
    .Y(_06684_));
 sky130_fd_sc_hd__inv_1 _11957_ (.A(_06678_),
    .Y(_06627_));
 sky130_fd_sc_hd__inv_1 _11958_ (.A(_06711_),
    .Y(_06707_));
 sky130_fd_sc_hd__inv_1 _11959_ (.A(_06727_),
    .Y(_06736_));
 sky130_fd_sc_hd__inv_1 _11960_ (.A(_06731_),
    .Y(_06686_));
 sky130_fd_sc_hd__inv_1 _11961_ (.A(_06768_),
    .Y(_06764_));
 sky130_fd_sc_hd__inv_1 _11962_ (.A(_06780_),
    .Y(_06738_));
 sky130_fd_sc_hd__inv_1 _11963_ (.A(_06787_),
    .Y(_06800_));
 sky130_fd_sc_hd__inv_1 _11964_ (.A(_06822_),
    .Y(_06816_));
 sky130_fd_sc_hd__inv_1 _11965_ (.A(_06925_),
    .Y(_06919_));
 sky130_fd_sc_hd__inv_1 _11966_ (.A(_06972_),
    .Y(_06966_));
 sky130_fd_sc_hd__inv_1 _11967_ (.A(_07014_),
    .Y(_07008_));
 sky130_fd_sc_hd__inv_1 _11968_ (.A(_07025_),
    .Y(_07022_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(\samples_real[6][14] ),
    .A1(\samples_real[7][14] ),
    .S(_03181_),
    .X(_03690_));
 sky130_fd_sc_hd__a22o_1 _11970_ (.A1(\samples_real[3][14] ),
    .A2(_03208_),
    .B1(_03690_),
    .B2(_03169_),
    .X(_03691_));
 sky130_fd_sc_hd__inv_1 _11971_ (.A(\samples_real[1][14] ),
    .Y(_03692_));
 sky130_fd_sc_hd__a21oi_1 _11972_ (.A1(net580),
    .A2(_03692_),
    .B1(_03183_),
    .Y(_03693_));
 sky130_fd_sc_hd__a21oi_1 _11973_ (.A1(_03158_),
    .A2(\samples_real[2][14] ),
    .B1(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__buf_12 _11974_ (.A(_03209_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2i_1 _11975_ (.A0(\samples_real[4][14] ),
    .A1(\samples_real[5][14] ),
    .S(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_03147_),
    .B(_03201_),
    .Y(_03697_));
 sky130_fd_sc_hd__o22ai_1 _11977_ (.A1(_03148_),
    .A2(_03694_),
    .B1(_03696_),
    .B2(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__a21oi_1 _11978_ (.A1(_03166_),
    .A2(_03691_),
    .B1(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__nor2_1 _11979_ (.A(\samples_real[0][14] ),
    .B(_03207_),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_1 _11980_ (.A(_03699_),
    .B(_03700_),
    .Y(_07721_));
 sky130_fd_sc_hd__mux4_1 _11981_ (.A0(\samples_real[0][13] ),
    .A1(\samples_real[2][13] ),
    .A2(\samples_real[1][13] ),
    .A3(\samples_real[3][13] ),
    .S0(net56),
    .S1(net580),
    .X(_03701_));
 sky130_fd_sc_hd__mux4_1 _11982_ (.A0(\samples_real[4][13] ),
    .A1(\samples_real[5][13] ),
    .A2(\samples_real[6][13] ),
    .A3(\samples_real[7][13] ),
    .S0(net582),
    .S1(_03183_),
    .X(_03702_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(_03701_),
    .A1(_03702_),
    .S(_03185_),
    .X(_07726_));
 sky130_fd_sc_hd__mux4_1 _11984_ (.A0(\samples_real[0][15] ),
    .A1(\samples_real[2][15] ),
    .A2(\samples_real[1][15] ),
    .A3(\samples_real[3][15] ),
    .S0(net517),
    .S1(net67),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_1 _11985_ (.A0(\samples_real[4][15] ),
    .A1(\samples_real[5][15] ),
    .A2(\samples_real[6][15] ),
    .A3(\samples_real[7][15] ),
    .S0(net67),
    .S1(net636),
    .X(_03704_));
 sky130_fd_sc_hd__mux2_2 _11986_ (.A0(_03703_),
    .A1(_03704_),
    .S(net522),
    .X(_07736_));
 sky130_fd_sc_hd__mux4_1 _11987_ (.A0(\samples_real[0][12] ),
    .A1(\samples_real[2][12] ),
    .A2(\samples_real[1][12] ),
    .A3(\samples_real[3][12] ),
    .S0(net56),
    .S1(net580),
    .X(_03705_));
 sky130_fd_sc_hd__mux4_1 _11988_ (.A0(\samples_real[4][12] ),
    .A1(\samples_real[5][12] ),
    .A2(\samples_real[6][12] ),
    .A3(\samples_real[7][12] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03706_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(_03705_),
    .A1(_03706_),
    .S(_03148_),
    .X(_07740_));
 sky130_fd_sc_hd__mux4_1 _11990_ (.A0(\samples_real[0][11] ),
    .A1(\samples_real[2][11] ),
    .A2(\samples_real[1][11] ),
    .A3(\samples_real[3][11] ),
    .S0(net56),
    .S1(net580),
    .X(_03707_));
 sky130_fd_sc_hd__mux4_1 _11991_ (.A0(\samples_real[4][11] ),
    .A1(\samples_real[5][11] ),
    .A2(\samples_real[6][11] ),
    .A3(\samples_real[7][11] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03708_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(_03707_),
    .A1(_03708_),
    .S(_03185_),
    .X(_07745_));
 sky130_fd_sc_hd__a22oi_2 _11993_ (.A1(\samples_real[2][10] ),
    .A2(net535),
    .B1(_03198_),
    .B2(\samples_real[7][10] ),
    .Y(_03709_));
 sky130_fd_sc_hd__a22oi_2 _11994_ (.A1(\samples_real[4][10] ),
    .A2(net552),
    .B1(net547),
    .B2(\samples_real[1][10] ),
    .Y(_03710_));
 sky130_fd_sc_hd__and3_1 _11995_ (.A(_03183_),
    .B(net643),
    .C(\samples_real[3][10] ),
    .X(_03711_));
 sky130_fd_sc_hd__a22oi_1 _11996_ (.A1(\samples_real[5][10] ),
    .A2(net562),
    .B1(net613),
    .B2(\samples_real[6][10] ),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_03185_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__o31ai_2 _11998_ (.A1(_03148_),
    .A2(net556),
    .A3(_03711_),
    .B1(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__clkbuf_4 _11999_ (.A(_03176_),
    .X(_03715_));
 sky130_fd_sc_hd__nor2_1 _12000_ (.A(\samples_real[0][10] ),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__a31oi_4 _12001_ (.A1(_03709_),
    .A2(_03710_),
    .A3(_03714_),
    .B1(_03716_),
    .Y(_07750_));
 sky130_fd_sc_hd__a22o_1 _12002_ (.A1(\samples_real[3][9] ),
    .A2(_03208_),
    .B1(_03210_),
    .B2(\samples_real[6][9] ),
    .X(_03717_));
 sky130_fd_sc_hd__nand2_1 _12003_ (.A(_03166_),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__o21ai_0 _12004_ (.A1(_03158_),
    .A2(\samples_real[1][9] ),
    .B1(_03201_),
    .Y(_03719_));
 sky130_fd_sc_hd__o21ai_0 _12005_ (.A1(_03213_),
    .A2(_03380_),
    .B1(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__mux2i_1 _12006_ (.A0(\samples_real[4][9] ),
    .A1(\samples_real[5][9] ),
    .S(net643),
    .Y(_03721_));
 sky130_fd_sc_hd__nand3_1 _12007_ (.A(_03166_),
    .B(_03213_),
    .C(\samples_real[7][9] ),
    .Y(_03722_));
 sky130_fd_sc_hd__o211ai_1 _12008_ (.A1(_03166_),
    .A2(_03721_),
    .B1(_03722_),
    .C1(_03148_),
    .Y(_03723_));
 sky130_fd_sc_hd__o21ai_0 _12009_ (.A1(_03185_),
    .A2(_03720_),
    .B1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_1 _12010_ (.A(\samples_real[0][9] ),
    .B(_03715_),
    .Y(_03725_));
 sky130_fd_sc_hd__a21oi_2 _12011_ (.A1(_03718_),
    .A2(_03724_),
    .B1(_03725_),
    .Y(_07755_));
 sky130_fd_sc_hd__mux4_1 _12012_ (.A0(\samples_real[0][8] ),
    .A1(\samples_real[2][8] ),
    .A2(\samples_real[1][8] ),
    .A3(\samples_real[3][8] ),
    .S0(net606),
    .S1(_03213_),
    .X(_03726_));
 sky130_fd_sc_hd__mux4_1 _12013_ (.A0(\samples_real[4][8] ),
    .A1(\samples_real[5][8] ),
    .A2(\samples_real[6][8] ),
    .A3(\samples_real[7][8] ),
    .S0(_03209_),
    .S1(_03166_),
    .X(_03727_));
 sky130_fd_sc_hd__buf_6 _12014_ (.A(_03169_),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _12015_ (.A0(_03726_),
    .A1(_03727_),
    .S(_03728_),
    .X(_07760_));
 sky130_fd_sc_hd__mux4_1 _12016_ (.A0(\samples_real[0][7] ),
    .A1(\samples_real[2][7] ),
    .A2(\samples_real[1][7] ),
    .A3(\samples_real[3][7] ),
    .S0(net587),
    .S1(net580),
    .X(_03729_));
 sky130_fd_sc_hd__mux4_1 _12017_ (.A0(\samples_real[4][7] ),
    .A1(\samples_real[5][7] ),
    .A2(\samples_real[6][7] ),
    .A3(\samples_real[7][7] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(_03729_),
    .A1(_03730_),
    .S(_03148_),
    .X(_07765_));
 sky130_fd_sc_hd__mux2i_1 _12019_ (.A0(\samples_real[6][6] ),
    .A1(\samples_real[7][6] ),
    .S(_03695_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(\samples_real[5][6] ),
    .B(net561),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ai_0 _12021_ (.A1(_03201_),
    .A2(_03731_),
    .B1(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__inv_1 _12022_ (.A(\samples_real[2][6] ),
    .Y(_03734_));
 sky130_fd_sc_hd__a21oi_1 _12023_ (.A1(net66),
    .A2(_03734_),
    .B1(_03169_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21oi_1 _12024_ (.A1(_03201_),
    .A2(\samples_real[4][6] ),
    .B1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__mux2i_1 _12025_ (.A0(\samples_real[1][6] ),
    .A1(\samples_real[3][6] ),
    .S(_03166_),
    .Y(_03737_));
 sky130_fd_sc_hd__nand2b_1 _12026_ (.A_N(_03169_),
    .B(net643),
    .Y(_03738_));
 sky130_fd_sc_hd__o22ai_1 _12027_ (.A1(_03213_),
    .A2(_03736_),
    .B1(_03737_),
    .B2(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__a21oi_1 _12028_ (.A1(_03728_),
    .A2(_03733_),
    .B1(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__nor2_1 _12029_ (.A(\samples_real[0][6] ),
    .B(_03207_),
    .Y(_03741_));
 sky130_fd_sc_hd__nor2_2 _12030_ (.A(_03740_),
    .B(_03741_),
    .Y(_07770_));
 sky130_fd_sc_hd__mux4_1 _12031_ (.A0(\samples_real[0][5] ),
    .A1(\samples_real[2][5] ),
    .A2(\samples_real[1][5] ),
    .A3(\samples_real[3][5] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03742_));
 sky130_fd_sc_hd__mux4_1 _12032_ (.A0(\samples_real[4][5] ),
    .A1(\samples_real[5][5] ),
    .A2(\samples_real[6][5] ),
    .A3(\samples_real[7][5] ),
    .S0(net583),
    .S1(net66),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _12033_ (.A0(_03742_),
    .A1(_03743_),
    .S(_03185_),
    .X(_07775_));
 sky130_fd_sc_hd__mux4_1 _12034_ (.A0(\samples_real[0][4] ),
    .A1(\samples_real[2][4] ),
    .A2(\samples_real[1][4] ),
    .A3(\samples_real[3][4] ),
    .S0(net586),
    .S1(net580),
    .X(_03744_));
 sky130_fd_sc_hd__mux4_1 _12035_ (.A0(\samples_real[4][4] ),
    .A1(\samples_real[5][4] ),
    .A2(\samples_real[6][4] ),
    .A3(\samples_real[7][4] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(_03744_),
    .A1(_03745_),
    .S(_03185_),
    .X(_07780_));
 sky130_fd_sc_hd__mux4_2 _12037_ (.A0(\samples_real[0][3] ),
    .A1(\samples_real[2][3] ),
    .A2(\samples_real[1][3] ),
    .A3(\samples_real[3][3] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03746_));
 sky130_fd_sc_hd__mux4_1 _12038_ (.A0(\samples_real[4][3] ),
    .A1(\samples_real[5][3] ),
    .A2(\samples_real[6][3] ),
    .A3(\samples_real[7][3] ),
    .S0(net582),
    .S1(net601),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_2 _12039_ (.A0(_03746_),
    .A1(_03747_),
    .S(_03728_),
    .X(_07785_));
 sky130_fd_sc_hd__mux4_1 _12040_ (.A0(\samples_real[0][2] ),
    .A1(\samples_real[2][2] ),
    .A2(\samples_real[1][2] ),
    .A3(\samples_real[3][2] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03748_));
 sky130_fd_sc_hd__mux4_1 _12041_ (.A0(\samples_real[4][2] ),
    .A1(\samples_real[5][2] ),
    .A2(\samples_real[6][2] ),
    .A3(\samples_real[7][2] ),
    .S0(net582),
    .S1(net600),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_4 _12042_ (.A0(_03748_),
    .A1(_03749_),
    .S(_03728_),
    .X(_07790_));
 sky130_fd_sc_hd__inv_1 _12043_ (.A(\sample_count[0] ),
    .Y(_07827_));
 sky130_fd_sc_hd__mux4_1 _12044_ (.A0(\samples_imag[1][14] ),
    .A1(\samples_imag[3][14] ),
    .A2(\samples_imag[5][14] ),
    .A3(\samples_imag[7][14] ),
    .S0(net55),
    .S1(_03169_),
    .X(_03750_));
 sky130_fd_sc_hd__mux2i_1 _12045_ (.A0(\samples_imag[4][14] ),
    .A1(\samples_imag[6][14] ),
    .S(net66),
    .Y(_03751_));
 sky130_fd_sc_hd__nor2_1 _12046_ (.A(\samples_imag[2][14] ),
    .B(_03155_),
    .Y(_03752_));
 sky130_fd_sc_hd__a211oi_1 _12047_ (.A1(_03728_),
    .A2(_03751_),
    .B1(_03752_),
    .C1(_03213_),
    .Y(_03753_));
 sky130_fd_sc_hd__a21oi_1 _12048_ (.A1(_03213_),
    .A2(_03750_),
    .B1(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__nor2_1 _12049_ (.A(\samples_imag[0][14] ),
    .B(_03207_),
    .Y(_03755_));
 sky130_fd_sc_hd__nor2_1 _12050_ (.A(_03754_),
    .B(_03755_),
    .Y(_07835_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(\samples_imag[0][13] ),
    .B(net584),
    .Y(_03756_));
 sky130_fd_sc_hd__mux2i_1 _12052_ (.A0(\samples_imag[6][13] ),
    .A1(\samples_imag[7][13] ),
    .S(net546),
    .Y(_03757_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(\samples_imag[5][13] ),
    .B(net559),
    .Y(_03758_));
 sky130_fd_sc_hd__o21ai_0 _12054_ (.A1(_03201_),
    .A2(_03757_),
    .B1(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__mux2i_1 _12055_ (.A0(\samples_imag[2][13] ),
    .A1(\samples_imag[3][13] ),
    .S(_03181_),
    .Y(_03760_));
 sky130_fd_sc_hd__inv_1 _12056_ (.A(\samples_imag[1][13] ),
    .Y(_03761_));
 sky130_fd_sc_hd__a21oi_1 _12057_ (.A1(net546),
    .A2(_03761_),
    .B1(_03146_),
    .Y(_03762_));
 sky130_fd_sc_hd__a21oi_1 _12058_ (.A1(_03158_),
    .A2(\samples_imag[4][13] ),
    .B1(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__o22ai_1 _12059_ (.A1(net539),
    .A2(_03760_),
    .B1(_03763_),
    .B2(net55),
    .Y(_03764_));
 sky130_fd_sc_hd__a21oi_1 _12060_ (.A1(_03147_),
    .A2(_03759_),
    .B1(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_2 _12061_ (.A(_03756_),
    .B(_03765_),
    .Y(_07840_));
 sky130_fd_sc_hd__mux4_1 _12062_ (.A0(\samples_imag[1][15] ),
    .A1(\samples_imag[3][15] ),
    .A2(\samples_imag[5][15] ),
    .A3(\samples_imag[7][15] ),
    .S0(net634),
    .S1(net521),
    .X(_03766_));
 sky130_fd_sc_hd__mux2i_1 _12063_ (.A0(\samples_imag[4][15] ),
    .A1(\samples_imag[6][15] ),
    .S(net635),
    .Y(_03767_));
 sky130_fd_sc_hd__nor2_1 _12064_ (.A(\samples_imag[2][15] ),
    .B(net539),
    .Y(_03768_));
 sky130_fd_sc_hd__a211oi_1 _12065_ (.A1(net521),
    .A2(_03767_),
    .B1(_03768_),
    .C1(net67),
    .Y(_03769_));
 sky130_fd_sc_hd__a21oi_1 _12066_ (.A1(net67),
    .A2(_03766_),
    .B1(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__nor2_1 _12067_ (.A(\samples_imag[0][15] ),
    .B(net584),
    .Y(_03771_));
 sky130_fd_sc_hd__nor2_4 _12068_ (.A(_03770_),
    .B(_03771_),
    .Y(_07850_));
 sky130_fd_sc_hd__inv_1 _12069_ (.A(\samples_imag[5][12] ),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_4 _12070_ (.A(_03147_),
    .B(net560),
    .Y(_03773_));
 sky130_fd_sc_hd__a2bb2oi_1 _12071_ (.A1_N(_03772_),
    .A2_N(_03773_),
    .B1(net548),
    .B2(\samples_imag[1][12] ),
    .Y(_03774_));
 sky130_fd_sc_hd__mux2i_1 _12072_ (.A0(\samples_imag[4][12] ),
    .A1(\samples_imag[6][12] ),
    .S(net55),
    .Y(_03775_));
 sky130_fd_sc_hd__o21ai_0 _12073_ (.A1(\samples_imag[2][12] ),
    .A2(net538),
    .B1(_03158_),
    .Y(_03776_));
 sky130_fd_sc_hd__a21oi_1 _12074_ (.A1(_03148_),
    .A2(_03775_),
    .B1(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__a221oi_1 _12075_ (.A1(\samples_imag[3][12] ),
    .A2(_03159_),
    .B1(_03198_),
    .B2(\samples_imag[7][12] ),
    .C1(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__nor2_2 _12076_ (.A(\samples_imag[0][12] ),
    .B(_03207_),
    .Y(_03779_));
 sky130_fd_sc_hd__a21oi_2 _12077_ (.A1(_03774_),
    .A2(_03778_),
    .B1(_03779_),
    .Y(_07854_));
 sky130_fd_sc_hd__mux4_1 _12078_ (.A0(\samples_imag[1][11] ),
    .A1(\samples_imag[3][11] ),
    .A2(\samples_imag[5][11] ),
    .A3(\samples_imag[7][11] ),
    .S0(_03182_),
    .S1(_03169_),
    .X(_03780_));
 sky130_fd_sc_hd__mux2i_1 _12079_ (.A0(\samples_imag[4][11] ),
    .A1(\samples_imag[6][11] ),
    .S(net55),
    .Y(_03781_));
 sky130_fd_sc_hd__nor2_1 _12080_ (.A(\samples_imag[2][11] ),
    .B(_03155_),
    .Y(_03782_));
 sky130_fd_sc_hd__a211oi_1 _12081_ (.A1(_03148_),
    .A2(_03781_),
    .B1(_03782_),
    .C1(_03213_),
    .Y(_03783_));
 sky130_fd_sc_hd__a21oi_1 _12082_ (.A1(_03213_),
    .A2(_03780_),
    .B1(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__nor2_1 _12083_ (.A(\samples_imag[0][11] ),
    .B(_03207_),
    .Y(_03785_));
 sky130_fd_sc_hd__nor2_1 _12084_ (.A(_03784_),
    .B(_03785_),
    .Y(_07859_));
 sky130_fd_sc_hd__mux4_1 _12085_ (.A0(\samples_imag[0][10] ),
    .A1(\samples_imag[2][10] ),
    .A2(\samples_imag[1][10] ),
    .A3(\samples_imag[3][10] ),
    .S0(net56),
    .S1(net580),
    .X(_03786_));
 sky130_fd_sc_hd__mux4_1 _12086_ (.A0(\samples_imag[4][10] ),
    .A1(\samples_imag[5][10] ),
    .A2(\samples_imag[6][10] ),
    .A3(\samples_imag[7][10] ),
    .S0(_03181_),
    .S1(net604),
    .X(_03787_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(_03786_),
    .A1(_03787_),
    .S(_03148_),
    .X(_07864_));
 sky130_fd_sc_hd__mux4_1 _12088_ (.A0(\samples_imag[2][9] ),
    .A1(\samples_imag[3][9] ),
    .A2(\samples_imag[6][9] ),
    .A3(\samples_imag[7][9] ),
    .S0(net640),
    .S1(_03169_),
    .X(_03788_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_03166_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__mux2i_1 _12090_ (.A0(\samples_imag[4][9] ),
    .A1(\samples_imag[5][9] ),
    .S(_03695_),
    .Y(_03790_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_03728_),
    .B(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__o211ai_1 _12092_ (.A1(\samples_imag[1][9] ),
    .A2(_03738_),
    .B1(_03791_),
    .C1(_03201_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(\samples_imag[0][9] ),
    .B(_03207_),
    .Y(_03793_));
 sky130_fd_sc_hd__a21oi_2 _12094_ (.A1(_03789_),
    .A2(_03792_),
    .B1(_03793_),
    .Y(_07869_));
 sky130_fd_sc_hd__mux4_1 _12095_ (.A0(\samples_imag[0][8] ),
    .A1(\samples_imag[2][8] ),
    .A2(\samples_imag[1][8] ),
    .A3(\samples_imag[3][8] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03794_));
 sky130_fd_sc_hd__mux4_1 _12096_ (.A0(\samples_imag[4][8] ),
    .A1(\samples_imag[5][8] ),
    .A2(\samples_imag[6][8] ),
    .A3(\samples_imag[7][8] ),
    .S0(net574),
    .S1(net66),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_2 _12097_ (.A0(_03794_),
    .A1(_03795_),
    .S(_03728_),
    .X(_07874_));
 sky130_fd_sc_hd__mux4_1 _12098_ (.A0(\samples_imag[0][7] ),
    .A1(\samples_imag[2][7] ),
    .A2(\samples_imag[1][7] ),
    .A3(\samples_imag[3][7] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03796_));
 sky130_fd_sc_hd__mux4_1 _12099_ (.A0(\samples_imag[4][7] ),
    .A1(\samples_imag[5][7] ),
    .A2(\samples_imag[6][7] ),
    .A3(\samples_imag[7][7] ),
    .S0(net574),
    .S1(net66),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_2 _12100_ (.A0(_03796_),
    .A1(_03797_),
    .S(_03728_),
    .X(_07879_));
 sky130_fd_sc_hd__mux4_1 _12101_ (.A0(\samples_imag[0][6] ),
    .A1(\samples_imag[2][6] ),
    .A2(\samples_imag[1][6] ),
    .A3(\samples_imag[3][6] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03798_));
 sky130_fd_sc_hd__mux4_1 _12102_ (.A0(\samples_imag[4][6] ),
    .A1(\samples_imag[5][6] ),
    .A2(\samples_imag[6][6] ),
    .A3(\samples_imag[7][6] ),
    .S0(net640),
    .S1(_03166_),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _12103_ (.A0(_03798_),
    .A1(_03799_),
    .S(_03728_),
    .X(_07884_));
 sky130_fd_sc_hd__mux4_1 _12104_ (.A0(\samples_imag[0][5] ),
    .A1(\samples_imag[2][5] ),
    .A2(\samples_imag[1][5] ),
    .A3(\samples_imag[3][5] ),
    .S0(net607),
    .S1(net580),
    .X(_03800_));
 sky130_fd_sc_hd__mux4_1 _12105_ (.A0(\samples_imag[4][5] ),
    .A1(\samples_imag[5][5] ),
    .A2(\samples_imag[6][5] ),
    .A3(\samples_imag[7][5] ),
    .S0(_03181_),
    .S1(_03183_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _12106_ (.A0(_03800_),
    .A1(_03801_),
    .S(_03185_),
    .X(_07889_));
 sky130_fd_sc_hd__mux4_1 _12107_ (.A0(\samples_imag[0][4] ),
    .A1(\samples_imag[2][4] ),
    .A2(\samples_imag[1][4] ),
    .A3(\samples_imag[3][4] ),
    .S0(_03182_),
    .S1(net580),
    .X(_03802_));
 sky130_fd_sc_hd__mux4_1 _12108_ (.A0(\samples_imag[4][4] ),
    .A1(\samples_imag[5][4] ),
    .A2(\samples_imag[6][4] ),
    .A3(\samples_imag[7][4] ),
    .S0(net574),
    .S1(net603),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_2 _12109_ (.A0(_03802_),
    .A1(_03803_),
    .S(_03185_),
    .X(_07894_));
 sky130_fd_sc_hd__mux4_1 _12110_ (.A0(\samples_imag[0][3] ),
    .A1(\samples_imag[2][3] ),
    .A2(\samples_imag[1][3] ),
    .A3(\samples_imag[3][3] ),
    .S0(_03182_),
    .S1(_03695_),
    .X(_03804_));
 sky130_fd_sc_hd__mux4_2 _12111_ (.A0(\samples_imag[4][3] ),
    .A1(\samples_imag[5][3] ),
    .A2(\samples_imag[6][3] ),
    .A3(\samples_imag[7][3] ),
    .S0(net574),
    .S1(net601),
    .X(_03805_));
 sky130_fd_sc_hd__mux2_4 _12112_ (.A0(_03804_),
    .A1(_03805_),
    .S(_03728_),
    .X(_07899_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(\samples_imag[6][2] ),
    .A1(\samples_imag[7][2] ),
    .S(net576),
    .X(_03806_));
 sky130_fd_sc_hd__a22o_1 _12114_ (.A1(\samples_imag[3][2] ),
    .A2(_03208_),
    .B1(_03806_),
    .B2(_03146_),
    .X(_03807_));
 sky130_fd_sc_hd__o21ai_0 _12115_ (.A1(_03151_),
    .A2(\samples_imag[1][2] ),
    .B1(_03201_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21boi_0 _12116_ (.A1(_03158_),
    .A2(\samples_imag[2][2] ),
    .B1_N(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__mux2i_2 _12117_ (.A0(\samples_imag[4][2] ),
    .A1(\samples_imag[5][2] ),
    .S(_03181_),
    .Y(_03810_));
 sky130_fd_sc_hd__o22ai_1 _12118_ (.A1(_03147_),
    .A2(_03809_),
    .B1(_03810_),
    .B2(_03697_),
    .Y(_03811_));
 sky130_fd_sc_hd__a21oi_2 _12119_ (.A1(_03807_),
    .A2(_03183_),
    .B1(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__nor2_1 _12120_ (.A(\samples_imag[0][2] ),
    .B(_03175_),
    .Y(_03813_));
 sky130_fd_sc_hd__nor2_4 _12121_ (.A(_03813_),
    .B(_03812_),
    .Y(_07904_));
 sky130_fd_sc_hd__inv_1 _12122_ (.A(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__inv_1 _12123_ (.A(_05929_),
    .Y(_05931_));
 sky130_fd_sc_hd__inv_1 _12124_ (.A(_05941_),
    .Y(_05976_));
 sky130_fd_sc_hd__inv_1 _12125_ (.A(_05911_),
    .Y(_05952_));
 sky130_fd_sc_hd__and2_0 _12126_ (.A(_03443_),
    .B(_03430_),
    .X(_05961_));
 sky130_fd_sc_hd__inv_1 _12127_ (.A(_07933_),
    .Y(_05989_));
 sky130_fd_sc_hd__inv_1 _12128_ (.A(_05946_),
    .Y(_05974_));
 sky130_fd_sc_hd__inv_1 _12129_ (.A(_05983_),
    .Y(_06065_));
 sky130_fd_sc_hd__inv_1 _12130_ (.A(_05939_),
    .Y(_05957_));
 sky130_fd_sc_hd__inv_1 _12131_ (.A(_06006_),
    .Y(_06022_));
 sky130_fd_sc_hd__inv_1 _12132_ (.A(_06009_),
    .Y(_06036_));
 sky130_fd_sc_hd__inv_1 _12133_ (.A(_07941_),
    .Y(_07944_));
 sky130_fd_sc_hd__inv_1 _12134_ (.A(_06016_),
    .Y(_06056_));
 sky130_fd_sc_hd__inv_1 _12135_ (.A(_05988_),
    .Y(_06063_));
 sky130_fd_sc_hd__inv_1 _12136_ (.A(_06043_),
    .Y(_06085_));
 sky130_fd_sc_hd__inv_1 _12137_ (.A(_06106_),
    .Y(_06102_));
 sky130_fd_sc_hd__inv_1 _12138_ (.A(_06094_),
    .Y(_06092_));
 sky130_fd_sc_hd__inv_1 _12139_ (.A(_07947_),
    .Y(_07951_));
 sky130_fd_sc_hd__inv_1 _12140_ (.A(_06105_),
    .Y(_06108_));
 sky130_fd_sc_hd__inv_1 _12141_ (.A(_06114_),
    .Y(_06112_));
 sky130_fd_sc_hd__inv_1 _12142_ (.A(_06076_),
    .Y(_06118_));
 sky130_fd_sc_hd__inv_1 _12143_ (.A(_06127_),
    .Y(_06171_));
 sky130_fd_sc_hd__inv_1 _12144_ (.A(_06152_),
    .Y(_06148_));
 sky130_fd_sc_hd__inv_1 _12145_ (.A(_06147_),
    .Y(_06187_));
 sky130_fd_sc_hd__inv_1 _12146_ (.A(_07923_),
    .Y(_07965_));
 sky130_fd_sc_hd__inv_1 _12147_ (.A(_06151_),
    .Y(_06158_));
 sky130_fd_sc_hd__inv_1 _12148_ (.A(_06163_),
    .Y(_06161_));
 sky130_fd_sc_hd__inv_1 _12149_ (.A(_06167_),
    .Y(_06165_));
 sky130_fd_sc_hd__inv_1 _12150_ (.A(_06177_),
    .Y(_06231_));
 sky130_fd_sc_hd__inv_1 _12151_ (.A(_06198_),
    .Y(_06247_));
 sky130_fd_sc_hd__inv_1 _12152_ (.A(_07987_),
    .Y(_07976_));
 sky130_fd_sc_hd__inv_1 _12153_ (.A(_06208_),
    .Y(_07981_));
 sky130_fd_sc_hd__inv_1 _12154_ (.A(_06209_),
    .Y(_06218_));
 sky130_fd_sc_hd__inv_1 _12155_ (.A(_06223_),
    .Y(_06221_));
 sky130_fd_sc_hd__inv_1 _12156_ (.A(_06227_),
    .Y(_06225_));
 sky130_fd_sc_hd__inv_1 _12157_ (.A(_06237_),
    .Y(_06281_));
 sky130_fd_sc_hd__inv_1 _12158_ (.A(_07997_),
    .Y(_05925_));
 sky130_fd_sc_hd__inv_1 _12159_ (.A(_06258_),
    .Y(_07992_));
 sky130_fd_sc_hd__inv_1 _12160_ (.A(_06259_),
    .Y(_06268_));
 sky130_fd_sc_hd__inv_1 _12161_ (.A(_06273_),
    .Y(_06271_));
 sky130_fd_sc_hd__inv_1 _12162_ (.A(_06277_),
    .Y(_06275_));
 sky130_fd_sc_hd__inv_1 _12163_ (.A(_06310_),
    .Y(_06305_));
 sky130_fd_sc_hd__inv_1 _12164_ (.A(_05942_),
    .Y(_07927_));
 sky130_fd_sc_hd__inv_1 _12165_ (.A(_06324_),
    .Y(_06321_));
 sky130_fd_sc_hd__inv_1 _12166_ (.A(_08008_),
    .Y(_06348_));
 sky130_fd_sc_hd__inv_1 _12167_ (.A(_05984_),
    .Y(_07934_));
 sky130_fd_sc_hd__inv_1 _12168_ (.A(_06456_),
    .Y(_06452_));
 sky130_fd_sc_hd__inv_2 _12169_ (.A(_06409_),
    .Y(_06404_));
 sky130_fd_sc_hd__inv_1 _12170_ (.A(_08023_),
    .Y(_06384_));
 sky130_fd_sc_hd__inv_1 _12171_ (.A(_08041_),
    .Y(_06072_));
 sky130_fd_sc_hd__inv_1 _12172_ (.A(_06366_),
    .Y(_06396_));
 sky130_fd_sc_hd__inv_1 _12173_ (.A(_06432_),
    .Y(_06427_));
 sky130_fd_sc_hd__inv_1 _12174_ (.A(_08039_),
    .Y(_06411_));
 sky130_fd_sc_hd__inv_1 _12175_ (.A(_07958_),
    .Y(_08043_));
 sky130_fd_sc_hd__inv_1 _12176_ (.A(_06403_),
    .Y(_06423_));
 sky130_fd_sc_hd__inv_1 _12177_ (.A(_06463_),
    .Y(_06458_));
 sky130_fd_sc_hd__inv_1 _12178_ (.A(_08054_),
    .Y(_08057_));
 sky130_fd_sc_hd__inv_2 _12179_ (.A(_06450_),
    .Y(_06447_));
 sky130_fd_sc_hd__inv_1 _12180_ (.A(_08065_),
    .Y(_08067_));
 sky130_fd_sc_hd__inv_1 _12181_ (.A(_08061_),
    .Y(_06477_));
 sky130_fd_sc_hd__mux2_1 _12182_ (.A0(_03402_),
    .A1(_08065_),
    .S(net484),
    .X(_03814_));
 sky130_fd_sc_hd__nand2_1 _12183_ (.A(_03313_),
    .B(_03814_),
    .Y(_06475_));
 sky130_fd_sc_hd__inv_1 _12184_ (.A(_08062_),
    .Y(_08075_));
 sky130_fd_sc_hd__inv_1 _12185_ (.A(_08088_),
    .Y(_06482_));
 sky130_fd_sc_hd__inv_1 _12186_ (.A(_08081_),
    .Y(_08100_));
 sky130_fd_sc_hd__inv_1 _12187_ (.A(_06329_),
    .Y(_06326_));
 sky130_fd_sc_hd__inv_1 _12188_ (.A(_06495_),
    .Y(_06512_));
 sky130_fd_sc_hd__inv_1 _12189_ (.A(_06504_),
    .Y(_06509_));
 sky130_fd_sc_hd__inv_1 _12190_ (.A(_06505_),
    .Y(_06514_));
 sky130_fd_sc_hd__inv_1 _12191_ (.A(_08111_),
    .Y(_08109_));
 sky130_fd_sc_hd__inv_1 _12192_ (.A(_06554_),
    .Y(_06572_));
 sky130_fd_sc_hd__inv_2 _12193_ (.A(_06544_),
    .Y(_06560_));
 sky130_fd_sc_hd__inv_1 _12194_ (.A(_06579_),
    .Y(_06602_));
 sky130_fd_sc_hd__nor3_1 _12195_ (.A(_03504_),
    .B(_03261_),
    .C(_03264_),
    .Y(_08144_));
 sky130_fd_sc_hd__inv_1 _12196_ (.A(_06611_),
    .Y(_06621_));
 sky130_fd_sc_hd__inv_1 _12197_ (.A(_06601_),
    .Y(_08149_));
 sky130_fd_sc_hd__inv_1 _12198_ (.A(_06609_),
    .Y(_06665_));
 sky130_fd_sc_hd__nor3_1 _12199_ (.A(_03504_),
    .B(net495),
    .C(_03311_),
    .Y(_08153_));
 sky130_fd_sc_hd__inv_1 _12200_ (.A(_06670_),
    .Y(_06680_));
 sky130_fd_sc_hd__inv_1 _12201_ (.A(_06645_),
    .Y(_08167_));
 sky130_fd_sc_hd__inv_1 _12202_ (.A(_06664_),
    .Y(_08171_));
 sky130_fd_sc_hd__inv_1 _12203_ (.A(_06669_),
    .Y(_06716_));
 sky130_fd_sc_hd__inv_1 _12204_ (.A(_06660_),
    .Y(_06709_));
 sky130_fd_sc_hd__nor2_1 _12205_ (.A(_03504_),
    .B(_03324_),
    .Y(_08174_));
 sky130_fd_sc_hd__inv_1 _12206_ (.A(_06700_),
    .Y(_06745_));
 sky130_fd_sc_hd__inv_1 _12207_ (.A(_06720_),
    .Y(_06770_));
 sky130_fd_sc_hd__and2_0 _12208_ (.A(_03431_),
    .B(_03332_),
    .X(_08186_));
 sky130_fd_sc_hd__inv_1 _12209_ (.A(_06751_),
    .Y(_06793_));
 sky130_fd_sc_hd__inv_1 _12210_ (.A(_06753_),
    .Y(_08196_));
 sky130_fd_sc_hd__inv_1 _12211_ (.A(_06774_),
    .Y(_06824_));
 sky130_fd_sc_hd__nor3_1 _12212_ (.A(_03504_),
    .B(_03344_),
    .C(net480),
    .Y(_08199_));
 sky130_fd_sc_hd__inv_1 _12213_ (.A(_06831_),
    .Y(_06836_));
 sky130_fd_sc_hd__inv_1 _12214_ (.A(_06799_),
    .Y(_06849_));
 sky130_fd_sc_hd__inv_1 _12215_ (.A(_06802_),
    .Y(_08209_));
 sky130_fd_sc_hd__inv_1 _12216_ (.A(_06762_),
    .Y(_06808_));
 sky130_fd_sc_hd__inv_1 _12217_ (.A(_06830_),
    .Y(_06880_));
 sky130_fd_sc_hd__nor3_1 _12218_ (.A(_03503_),
    .B(net438),
    .C(_03363_),
    .Y(_08214_));
 sky130_fd_sc_hd__inv_1 _12219_ (.A(_06888_),
    .Y(_06890_));
 sky130_fd_sc_hd__inv_1 _12220_ (.A(_06843_),
    .Y(_06856_));
 sky130_fd_sc_hd__inv_1 _12221_ (.A(_06814_),
    .Y(_06865_));
 sky130_fd_sc_hd__inv_1 _12222_ (.A(_06832_),
    .Y(_06882_));
 sky130_fd_sc_hd__and2_0 _12223_ (.A(_03431_),
    .B(_03371_),
    .X(_08229_));
 sky130_fd_sc_hd__inv_1 _12224_ (.A(_06902_),
    .Y(_08232_));
 sky130_fd_sc_hd__inv_1 _12225_ (.A(_06929_),
    .Y(_08240_));
 sky130_fd_sc_hd__nor2_1 _12226_ (.A(_03504_),
    .B(net503),
    .Y(_08245_));
 sky130_fd_sc_hd__inv_1 _12227_ (.A(_06974_),
    .Y(_06976_));
 sky130_fd_sc_hd__inv_1 _12228_ (.A(_06941_),
    .Y(_06951_));
 sky130_fd_sc_hd__inv_1 _12229_ (.A(_06950_),
    .Y(_06987_));
 sky130_fd_sc_hd__inv_1 _12230_ (.A(_06921_),
    .Y(_06960_));
 sky130_fd_sc_hd__inv_1 _12231_ (.A(_06942_),
    .Y(_06971_));
 sky130_fd_sc_hd__inv_1 _12232_ (.A(_06932_),
    .Y(_08253_));
 sky130_fd_sc_hd__and2_0 _12233_ (.A(_03431_),
    .B(net483),
    .X(_08259_));
 sky130_fd_sc_hd__inv_1 _12234_ (.A(_06984_),
    .Y(_06993_));
 sky130_fd_sc_hd__inv_1 _12235_ (.A(_06968_),
    .Y(_07002_));
 sky130_fd_sc_hd__inv_1 _12236_ (.A(_06985_),
    .Y(_07013_));
 sky130_fd_sc_hd__and2_0 _12237_ (.A(_00012_),
    .B(_03402_),
    .X(_08270_));
 sky130_fd_sc_hd__inv_1 _12238_ (.A(_07024_),
    .Y(_08278_));
 sky130_fd_sc_hd__inv_1 _12239_ (.A(_07030_),
    .Y(_08282_));
 sky130_fd_sc_hd__inv_1 _12240_ (.A(_07010_),
    .Y(_07036_));
 sky130_fd_sc_hd__inv_1 _12241_ (.A(_07031_),
    .Y(_07041_));
 sky130_fd_sc_hd__nor3_1 _12242_ (.A(_03503_),
    .B(_03407_),
    .C(_03408_),
    .Y(_08288_));
 sky130_fd_sc_hd__inv_1 _12243_ (.A(_07051_),
    .Y(_08297_));
 sky130_fd_sc_hd__nor2_1 _12244_ (.A(_03504_),
    .B(net501),
    .Y(_08302_));
 sky130_fd_sc_hd__inv_1 _12245_ (.A(_07072_),
    .Y(_07079_));
 sky130_fd_sc_hd__inv_1 _12246_ (.A(_07073_),
    .Y(_07082_));
 sky130_fd_sc_hd__and2_0 _12247_ (.A(_00012_),
    .B(_03458_),
    .X(_08333_));
 sky130_fd_sc_hd__o21a_1 _12248_ (.A1(_07113_),
    .A2(_00640_),
    .B1(_00644_),
    .X(_07122_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_00686_),
    .B(_00689_),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_00627_),
    .B(_00649_),
    .Y(_07134_));
 sky130_fd_sc_hd__a21bo_1 _12251_ (.A1(_00648_),
    .A2(_07125_),
    .B1_N(_00693_),
    .X(_07137_));
 sky130_fd_sc_hd__clkinv_2 _12252_ (.A(_00767_),
    .Y(_07140_));
 sky130_fd_sc_hd__inv_1 _12253_ (.A(_00870_),
    .Y(_07143_));
 sky130_fd_sc_hd__inv_1 _12254_ (.A(_07134_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand2_1 _12255_ (.A(_00674_),
    .B(net6),
    .Y(_03816_));
 sky130_fd_sc_hd__o21ai_2 _12256_ (.A1(net6),
    .A2(_03815_),
    .B1(_03816_),
    .Y(_07154_));
 sky130_fd_sc_hd__nor2_4 _12257_ (.A(_00690_),
    .B(_00697_),
    .Y(_03817_));
 sky130_fd_sc_hd__inv_2 _12258_ (.A(_03817_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand2_1 _12259_ (.A(_00675_),
    .B(_00772_),
    .Y(_03818_));
 sky130_fd_sc_hd__o21ai_0 _12260_ (.A1(_00675_),
    .A2(_00767_),
    .B1(_03818_),
    .Y(_07160_));
 sky130_fd_sc_hd__o211ai_1 _12261_ (.A1(_03815_),
    .A2(_00739_),
    .B1(_00676_),
    .C1(_00681_),
    .Y(_07167_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_00660_),
    .B(_00717_),
    .Y(_03819_));
 sky130_fd_sc_hd__o21ai_2 _12263_ (.A1(_00660_),
    .A2(_03817_),
    .B1(_03819_),
    .Y(_07170_));
 sky130_fd_sc_hd__nor2_1 _12264_ (.A(_00660_),
    .B(_07163_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_1 _12265_ (.A1(net36),
    .A2(_00876_),
    .B1(_03820_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(_00710_),
    .A2(_07170_),
    .B1(_00716_),
    .X(_07187_));
 sky130_fd_sc_hd__nor2_1 _12267_ (.A(_00698_),
    .B(_07173_),
    .Y(_03821_));
 sky130_fd_sc_hd__nor2_1 _12268_ (.A(_00775_),
    .B(_03821_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_00709_),
    .B(_00726_),
    .Y(_03822_));
 sky130_fd_sc_hd__a22o_1 _12270_ (.A1(_00683_),
    .A2(_03822_),
    .B1(_00842_),
    .B2(_00752_),
    .X(_07208_));
 sky130_fd_sc_hd__o22ai_1 _12271_ (.A1(_00797_),
    .A2(_00788_),
    .B1(_00824_),
    .B2(_00786_),
    .Y(_07211_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(_00869_),
    .B(_00825_),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(_03823_),
    .B(_00912_),
    .Y(_07214_));
 sky130_fd_sc_hd__inv_1 _12274_ (.A(_01227_),
    .Y(_07311_));
 sky130_fd_sc_hd__inv_1 _12275_ (.A(_02107_),
    .Y(_07491_));
 sky130_fd_sc_hd__nor2_1 _12276_ (.A(_07532_),
    .B(_02307_),
    .Y(_07551_));
 sky130_fd_sc_hd__inv_1 _12277_ (.A(_02688_),
    .Y(_07585_));
 sky130_fd_sc_hd__nor4_1 _12278_ (.A(_05887_),
    .B(_07726_),
    .C(_07736_),
    .D(_07760_),
    .Y(_03824_));
 sky130_fd_sc_hd__nor4_1 _12279_ (.A(_07740_),
    .B(_07745_),
    .C(_07775_),
    .D(_07790_),
    .Y(_03825_));
 sky130_fd_sc_hd__nor4_1 _12280_ (.A(_07755_),
    .B(_07765_),
    .C(_07780_),
    .D(_07785_),
    .Y(_03826_));
 sky130_fd_sc_hd__nor4_1 _12281_ (.A(_07732_),
    .B(_07721_),
    .C(_07750_),
    .D(_07770_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand4_1 _12282_ (.A(_03824_),
    .B(_03825_),
    .C(_03826_),
    .D(_03827_),
    .Y(_07737_));
 sky130_fd_sc_hd__inv_1 _12283_ (.A(_07815_),
    .Y(_07818_));
 sky130_fd_sc_hd__inv_1 _12284_ (.A(\sample_count[1] ),
    .Y(_07828_));
 sky130_fd_sc_hd__inv_1 _12285_ (.A(_07717_),
    .Y(_05894_));
 sky130_fd_sc_hd__or4_1 _12286_ (.A(net637),
    .B(_07840_),
    .C(_07850_),
    .D(_07904_),
    .X(_03828_));
 sky130_fd_sc_hd__nor4_1 _12287_ (.A(_07854_),
    .B(_07859_),
    .C(_07869_),
    .D(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__nor4_1 _12288_ (.A(_07864_),
    .B(_07889_),
    .C(_07894_),
    .D(_07899_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor2_1 _12289_ (.A(_05902_),
    .B(_07835_),
    .Y(_03831_));
 sky130_fd_sc_hd__nor3_1 _12290_ (.A(_07874_),
    .B(_07879_),
    .C(_07884_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand4_1 _12291_ (.A(_03829_),
    .B(_03830_),
    .C(_03831_),
    .D(_03832_),
    .Y(_07851_));
 sky130_fd_sc_hd__inv_1 _12292_ (.A(_05940_),
    .Y(_05934_));
 sky130_fd_sc_hd__inv_1 _12293_ (.A(_07925_),
    .Y(_05926_));
 sky130_fd_sc_hd__inv_1 _12294_ (.A(_07926_),
    .Y(_05927_));
 sky130_fd_sc_hd__inv_1 _12295_ (.A(_05982_),
    .Y(_05977_));
 sky130_fd_sc_hd__nor2_1 _12296_ (.A(_03504_),
    .B(_03246_),
    .Y(_05953_));
 sky130_fd_sc_hd__inv_1 _12297_ (.A(_06000_),
    .Y(_05966_));
 sky130_fd_sc_hd__inv_1 _12298_ (.A(_07937_),
    .Y(_05990_));
 sky130_fd_sc_hd__nor3_1 _12299_ (.A(_03503_),
    .B(_03334_),
    .C(net464),
    .Y(_06080_));
 sky130_fd_sc_hd__inv_1 _12300_ (.A(_06021_),
    .Y(_06023_));
 sky130_fd_sc_hd__inv_1 _12301_ (.A(_06045_),
    .Y(_06091_));
 sky130_fd_sc_hd__inv_1 _12302_ (.A(_06126_),
    .Y(_06120_));
 sky130_fd_sc_hd__inv_1 _12303_ (.A(_07949_),
    .Y(_06073_));
 sky130_fd_sc_hd__inv_1 _12304_ (.A(_07960_),
    .Y(_06074_));
 sky130_fd_sc_hd__nor3_1 _12305_ (.A(_03503_),
    .B(_03379_),
    .C(net505),
    .Y(_06133_));
 sky130_fd_sc_hd__inv_1 _12306_ (.A(_06140_),
    .Y(_06137_));
 sky130_fd_sc_hd__inv_1 _12307_ (.A(_06101_),
    .Y(_06144_));
 sky130_fd_sc_hd__inv_1 _12308_ (.A(_07922_),
    .Y(_07953_));
 sky130_fd_sc_hd__inv_1 _12309_ (.A(_06176_),
    .Y(_06172_));
 sky130_fd_sc_hd__inv_1 _12310_ (.A(_06191_),
    .Y(_06188_));
 sky130_fd_sc_hd__inv_1 _12311_ (.A(_07974_),
    .Y(_07966_));
 sky130_fd_sc_hd__inv_1 _12312_ (.A(_06236_),
    .Y(_06232_));
 sky130_fd_sc_hd__and2_0 _12313_ (.A(_00012_),
    .B(_03430_),
    .X(_06243_));
 sky130_fd_sc_hd__inv_1 _12314_ (.A(_07975_),
    .Y(_07977_));
 sky130_fd_sc_hd__nor2_1 _12315_ (.A(_03504_),
    .B(net456),
    .Y(_06293_));
 sky130_fd_sc_hd__inv_1 _12316_ (.A(_07988_),
    .Y(_05918_));
 sky130_fd_sc_hd__nor3_1 _12317_ (.A(_03503_),
    .B(_03448_),
    .C(_03450_),
    .Y(_06340_));
 sky130_fd_sc_hd__inv_1 _12318_ (.A(_06323_),
    .Y(_06320_));
 sky130_fd_sc_hd__inv_1 _12319_ (.A(_06304_),
    .Y(_06306_));
 sky130_fd_sc_hd__inv_1 _12320_ (.A(_07998_),
    .Y(_05935_));
 sky130_fd_sc_hd__inv_1 _12321_ (.A(_06372_),
    .Y(_06368_));
 sky130_fd_sc_hd__inv_1 _12322_ (.A(_08009_),
    .Y(_05978_));
 sky130_fd_sc_hd__inv_1 _12323_ (.A(_06362_),
    .Y(_06360_));
 sky130_fd_sc_hd__inv_1 _12324_ (.A(_06457_),
    .Y(_06453_));
 sky130_fd_sc_hd__inv_1 _12325_ (.A(_06410_),
    .Y(_06405_));
 sky130_fd_sc_hd__inv_1 _12326_ (.A(_08024_),
    .Y(_06067_));
 sky130_fd_sc_hd__inv_1 _12327_ (.A(_06399_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _12328_ (.A(_03431_),
    .B(_03475_),
    .Y(_08032_));
 sky130_fd_sc_hd__inv_1 _12329_ (.A(_06433_),
    .Y(_06428_));
 sky130_fd_sc_hd__inv_1 _12330_ (.A(_08042_),
    .Y(_06121_));
 sky130_fd_sc_hd__inv_1 _12331_ (.A(_06426_),
    .Y(_06424_));
 sky130_fd_sc_hd__inv_1 _12332_ (.A(_06464_),
    .Y(_06459_));
 sky130_fd_sc_hd__inv_1 _12333_ (.A(_06451_),
    .Y(_06448_));
 sky130_fd_sc_hd__inv_1 _12334_ (.A(_08077_),
    .Y(_08064_));
 sky130_fd_sc_hd__inv_1 _12335_ (.A(_07955_),
    .Y(_08068_));
 sky130_fd_sc_hd__inv_1 _12336_ (.A(_08073_),
    .Y(_06478_));
 sky130_fd_sc_hd__inv_1 _12337_ (.A(_08080_),
    .Y(_08076_));
 sky130_fd_sc_hd__inv_1 _12338_ (.A(_08084_),
    .Y(_08079_));
 sky130_fd_sc_hd__inv_1 _12339_ (.A(_08101_),
    .Y(_08087_));
 sky130_fd_sc_hd__inv_1 _12340_ (.A(_07982_),
    .Y(_06481_));
 sky130_fd_sc_hd__inv_1 _12341_ (.A(_06491_),
    .Y(_06489_));
 sky130_fd_sc_hd__inv_1 _12342_ (.A(_08089_),
    .Y(_08098_));
 sky130_fd_sc_hd__inv_1 _12343_ (.A(_06498_),
    .Y(_06283_));
 sky130_fd_sc_hd__inv_1 _12344_ (.A(_06516_),
    .Y(_06513_));
 sky130_fd_sc_hd__inv_1 _12345_ (.A(_06524_),
    .Y(_06517_));
 sky130_fd_sc_hd__inv_1 _12346_ (.A(_08110_),
    .Y(_08117_));
 sky130_fd_sc_hd__a21o_1 _12347_ (.A1(_08118_),
    .A2(_06367_),
    .B1(_08128_),
    .X(_08125_));
 sky130_fd_sc_hd__and2_4 _12348_ (.A(_03247_),
    .B(_03458_),
    .X(_06532_));
 sky130_fd_sc_hd__inv_1 _12349_ (.A(_06578_),
    .Y(_06573_));
 sky130_fd_sc_hd__inv_1 _12350_ (.A(_06566_),
    .Y(_06568_));
 sky130_fd_sc_hd__inv_1 _12351_ (.A(_06600_),
    .Y(_06569_));
 sky130_fd_sc_hd__inv_1 _12352_ (.A(_06606_),
    .Y(_06603_));
 sky130_fd_sc_hd__nor2_1 _12353_ (.A(_03501_),
    .B(_03499_),
    .Y(_08145_));
 sky130_fd_sc_hd__inv_1 _12354_ (.A(_06663_),
    .Y(_08150_));
 sky130_fd_sc_hd__inv_1 _12355_ (.A(_06668_),
    .Y(_06666_));
 sky130_fd_sc_hd__nor3_1 _12356_ (.A(_03501_),
    .B(_03261_),
    .C(_03264_),
    .Y(_08154_));
 sky130_fd_sc_hd__inv_1 _12357_ (.A(_06699_),
    .Y(_06694_));
 sky130_fd_sc_hd__inv_1 _12358_ (.A(_06719_),
    .Y(_06717_));
 sky130_fd_sc_hd__nor3_1 _12359_ (.A(_03501_),
    .B(net496),
    .C(_03311_),
    .Y(_08175_));
 sky130_fd_sc_hd__inv_1 _12360_ (.A(_06750_),
    .Y(_06746_));
 sky130_fd_sc_hd__inv_1 _12361_ (.A(_06773_),
    .Y(_06771_));
 sky130_fd_sc_hd__nor2_1 _12362_ (.A(_03501_),
    .B(net478),
    .Y(_08187_));
 sky130_fd_sc_hd__inv_1 _12363_ (.A(_06798_),
    .Y(_06794_));
 sky130_fd_sc_hd__inv_1 _12364_ (.A(_06760_),
    .Y(_06756_));
 sky130_fd_sc_hd__inv_1 _12365_ (.A(_06828_),
    .Y(_06825_));
 sky130_fd_sc_hd__and2_0 _12366_ (.A(_00009_),
    .B(_03332_),
    .X(_08200_));
 sky130_fd_sc_hd__inv_1 _12367_ (.A(_06854_),
    .Y(_06850_));
 sky130_fd_sc_hd__inv_1 _12368_ (.A(_06812_),
    .Y(_06809_));
 sky130_fd_sc_hd__inv_1 _12369_ (.A(_06885_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor3_1 _12370_ (.A(_03500_),
    .B(_03344_),
    .C(net480),
    .Y(_08215_));
 sky130_fd_sc_hd__inv_1 _12371_ (.A(_06848_),
    .Y(_06857_));
 sky130_fd_sc_hd__inv_1 _12372_ (.A(_06901_),
    .Y(_08217_));
 sky130_fd_sc_hd__inv_1 _12373_ (.A(_06869_),
    .Y(_06866_));
 sky130_fd_sc_hd__inv_1 _12374_ (.A(_06928_),
    .Y(_08224_));
 sky130_fd_sc_hd__nor3_1 _12375_ (.A(_03500_),
    .B(net439),
    .C(_03363_),
    .Y(_08230_));
 sky130_fd_sc_hd__inv_1 _12376_ (.A(_06918_),
    .Y(_06915_));
 sky130_fd_sc_hd__and2_0 _12377_ (.A(_00009_),
    .B(_03371_),
    .X(_08246_));
 sky130_fd_sc_hd__nor2_1 _12378_ (.A(_03501_),
    .B(net502),
    .Y(_08260_));
 sky130_fd_sc_hd__inv_1 _12379_ (.A(_07023_),
    .Y(_08262_));
 sky130_fd_sc_hd__inv_1 _12380_ (.A(_07006_),
    .Y(_07003_));
 sky130_fd_sc_hd__inv_1 _12381_ (.A(_06975_),
    .Y(_08267_));
 sky130_fd_sc_hd__and2_0 _12382_ (.A(_00009_),
    .B(net483),
    .X(_08271_));
 sky130_fd_sc_hd__inv_1 _12383_ (.A(_07050_),
    .Y(_08285_));
 sky130_fd_sc_hd__and2_0 _12384_ (.A(_00009_),
    .B(_03402_),
    .X(_08289_));
 sky130_fd_sc_hd__nor3_1 _12385_ (.A(_03500_),
    .B(_03407_),
    .C(_03408_),
    .Y(_08303_));
 sky130_fd_sc_hd__inv_1 _12386_ (.A(_07102_),
    .Y(_08330_));
 sky130_fd_sc_hd__nor2_1 _12387_ (.A(_03501_),
    .B(net499),
    .Y(_08334_));
 sky130_fd_sc_hd__inv_1 _12388_ (.A(_08074_),
    .Y(_08097_));
 sky130_fd_sc_hd__inv_1 _12389_ (.A(_08099_),
    .Y(_08107_));
 sky130_fd_sc_hd__inv_1 _12390_ (.A(_08148_),
    .Y(_06657_));
 sky130_fd_sc_hd__inv_1 _12391_ (.A(_08162_),
    .Y(_06637_));
 sky130_fd_sc_hd__inv_1 _12392_ (.A(_08177_),
    .Y(_06741_));
 sky130_fd_sc_hd__inv_1 _12393_ (.A(_08189_),
    .Y(_06789_));
 sky130_fd_sc_hd__inv_1 _12394_ (.A(_08202_),
    .Y(_06845_));
 sky130_fd_sc_hd__inv_1 _12395_ (.A(_08210_),
    .Y(_06876_));
 sky130_fd_sc_hd__inv_1 _12396_ (.A(_08275_),
    .Y(_07028_));
 sky130_fd_sc_hd__inv_1 _12397_ (.A(_08314_),
    .Y(_07096_));
 sky130_fd_sc_hd__inv_1 _12398_ (.A(_07930_),
    .Y(_05970_));
 sky130_fd_sc_hd__inv_1 _12399_ (.A(_07935_),
    .Y(_06060_));
 sky130_fd_sc_hd__inv_1 _12400_ (.A(_07946_),
    .Y(_06050_));
 sky130_fd_sc_hd__inv_1 _12401_ (.A(_07957_),
    .Y(_06173_));
 sky130_fd_sc_hd__inv_1 _12402_ (.A(_07962_),
    .Y(_06169_));
 sky130_fd_sc_hd__inv_1 _12403_ (.A(_07970_),
    .Y(_06233_));
 sky130_fd_sc_hd__inv_1 _12404_ (.A(_07971_),
    .Y(_06229_));
 sky130_fd_sc_hd__inv_1 _12405_ (.A(_07983_),
    .Y(_06279_));
 sky130_fd_sc_hd__inv_1 _12406_ (.A(_07985_),
    .Y(_06301_));
 sky130_fd_sc_hd__inv_1 _12407_ (.A(_08078_),
    .Y(_08086_));
 sky130_fd_sc_hd__inv_1 _12408_ (.A(_08085_),
    .Y(_08119_));
 sky130_fd_sc_hd__inv_1 _12409_ (.A(_08102_),
    .Y(_06497_));
 sky130_fd_sc_hd__inv_1 _12410_ (.A(_08228_),
    .Y(_06896_));
 sky130_fd_sc_hd__inv_1 _12411_ (.A(_08244_),
    .Y(_06939_));
 sky130_fd_sc_hd__inv_1 _12412_ (.A(_08258_),
    .Y(_06982_));
 sky130_fd_sc_hd__inv_1 _12413_ (.A(_07104_),
    .Y(_07101_));
 sky130_fd_sc_hd__inv_1 _12414_ (.A(_08272_),
    .Y(_07048_));
 sky130_fd_sc_hd__inv_1 _12415_ (.A(\sample_count[2] ),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _12416_ (.A(_03137_),
    .B(net91),
    .Y(_03834_));
 sky130_fd_sc_hd__clkbuf_2 _12417_ (.A(\bit_rev_idx[0] ),
    .X(_03835_));
 sky130_fd_sc_hd__nand2_1 _12418_ (.A(_03835_),
    .B(_03834_),
    .Y(_03836_));
 sky130_fd_sc_hd__o21ai_0 _12419_ (.A1(_03833_),
    .A2(_03834_),
    .B1(_03836_),
    .Y(_00024_));
 sky130_fd_sc_hd__clkbuf_2 _12420_ (.A(\bit_rev_idx[1] ),
    .X(_03837_));
 sky130_fd_sc_hd__nand2_1 _12421_ (.A(_03837_),
    .B(_03834_),
    .Y(_03838_));
 sky130_fd_sc_hd__o21ai_0 _12422_ (.A1(_07828_),
    .A2(_03834_),
    .B1(_03838_),
    .Y(_00025_));
 sky130_fd_sc_hd__clkbuf_2 _12423_ (.A(\bit_rev_idx[2] ),
    .X(_03839_));
 sky130_fd_sc_hd__nand2_1 _12424_ (.A(_03839_),
    .B(_03834_),
    .Y(_03840_));
 sky130_fd_sc_hd__o21ai_0 _12425_ (.A1(_07827_),
    .A2(_03834_),
    .B1(_03840_),
    .Y(_00026_));
 sky130_fd_sc_hd__inv_1 _12426_ (.A(net94),
    .Y(_03841_));
 sky130_fd_sc_hd__nor2_1 _12427_ (.A(_00557_),
    .B(_00559_),
    .Y(_03842_));
 sky130_fd_sc_hd__nor2_1 _12428_ (.A(net93),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__o21ai_0 _12429_ (.A1(_03842_),
    .A2(_03843_),
    .B1(\state[0] ),
    .Y(_03844_));
 sky130_fd_sc_hd__o21ai_0 _12430_ (.A1(_00560_),
    .A2(_03841_),
    .B1(_03844_),
    .Y(_00027_));
 sky130_fd_sc_hd__nor2_2 _12431_ (.A(_03137_),
    .B(\state[1] ),
    .Y(_03845_));
 sky130_fd_sc_hd__a211oi_4 _12432_ (.A1(_03137_),
    .A2(_03138_),
    .B1(_00003_),
    .C1(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand3_1 _12433_ (.A(_07716_),
    .B(_03144_),
    .C(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__o21ai_0 _12434_ (.A1(_07716_),
    .A2(_03846_),
    .B1(_03847_),
    .Y(_00028_));
 sky130_fd_sc_hd__nand3_1 _12435_ (.A(_07800_),
    .B(_03144_),
    .C(_03846_),
    .Y(_03848_));
 sky130_fd_sc_hd__o21ai_0 _12436_ (.A1(_07666_),
    .A2(_03846_),
    .B1(_03848_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand3_1 _12437_ (.A(_07801_),
    .B(_03144_),
    .C(_03846_),
    .Y(_03849_));
 sky130_fd_sc_hd__o21ai_0 _12438_ (.A1(_00811_),
    .A2(_03846_),
    .B1(_03849_),
    .Y(_00030_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(net95),
    .A1(\samples_imag[0][0] ),
    .S(_00560_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _12440_ (.A0(net96),
    .A1(\samples_imag[6][4] ),
    .S(_00560_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(net97),
    .A1(\samples_imag[6][5] ),
    .S(_00560_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _12442_ (.A0(net98),
    .A1(\samples_imag[6][6] ),
    .S(_00560_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(net99),
    .A1(\samples_imag[6][7] ),
    .S(_00560_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(net100),
    .A1(\samples_imag[6][8] ),
    .S(_00560_),
    .X(_00036_));
 sky130_fd_sc_hd__buf_6 _12445_ (.A(_00559_),
    .X(_03850_));
 sky130_fd_sc_hd__mux2_1 _12446_ (.A0(net101),
    .A1(\samples_imag[6][9] ),
    .S(_03850_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(net102),
    .A1(\samples_imag[6][10] ),
    .S(_03850_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _12448_ (.A0(net103),
    .A1(\samples_imag[6][11] ),
    .S(_03850_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(net104),
    .A1(\samples_imag[6][12] ),
    .S(_03850_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _12450_ (.A0(net105),
    .A1(\samples_imag[6][13] ),
    .S(_03850_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(net106),
    .A1(\samples_imag[0][10] ),
    .S(_03850_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _12452_ (.A0(net107),
    .A1(\samples_imag[6][14] ),
    .S(_03850_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(net108),
    .A1(\samples_imag[6][15] ),
    .S(_03850_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _12454_ (.A0(net109),
    .A1(\samples_imag[7][0] ),
    .S(_03850_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(net110),
    .A1(\samples_imag[7][1] ),
    .S(_03850_),
    .X(_00046_));
 sky130_fd_sc_hd__clkbuf_4 _12456_ (.A(_00559_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(net111),
    .A1(\samples_imag[7][2] ),
    .S(_03851_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _12458_ (.A0(net112),
    .A1(\samples_imag[7][3] ),
    .S(_03851_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(net113),
    .A1(\samples_imag[7][4] ),
    .S(_03851_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _12460_ (.A0(net114),
    .A1(\samples_imag[7][5] ),
    .S(_03851_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _12461_ (.A0(net115),
    .A1(\samples_imag[7][6] ),
    .S(_03851_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(net116),
    .A1(\samples_imag[7][7] ),
    .S(_03851_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(net117),
    .A1(\samples_imag[0][11] ),
    .S(_03851_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(net118),
    .A1(\samples_imag[7][8] ),
    .S(_03851_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _12465_ (.A0(net119),
    .A1(\samples_imag[7][9] ),
    .S(_03851_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(net120),
    .A1(\samples_imag[7][10] ),
    .S(_03851_),
    .X(_00056_));
 sky130_fd_sc_hd__buf_4 _12467_ (.A(_00559_),
    .X(_03852_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(net121),
    .A1(\samples_imag[7][11] ),
    .S(_03852_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(net122),
    .A1(\samples_imag[7][12] ),
    .S(_03852_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(net123),
    .A1(\samples_imag[7][13] ),
    .S(_03852_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(net124),
    .A1(\samples_imag[7][14] ),
    .S(_03852_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(net125),
    .A1(\samples_imag[7][15] ),
    .S(_03852_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _12473_ (.A0(net126),
    .A1(\samples_imag[0][12] ),
    .S(_03852_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(net127),
    .A1(\samples_imag[0][13] ),
    .S(_03852_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _12475_ (.A0(net128),
    .A1(\samples_imag[0][14] ),
    .S(_03852_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(net129),
    .A1(\samples_imag[0][15] ),
    .S(_03852_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _12477_ (.A0(net130),
    .A1(\samples_imag[1][0] ),
    .S(_03852_),
    .X(_00066_));
 sky130_fd_sc_hd__buf_6 _12478_ (.A(_00559_),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _12479_ (.A0(net131),
    .A1(\samples_imag[1][1] ),
    .S(_03853_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(net132),
    .A1(\samples_imag[1][2] ),
    .S(_03853_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(net133),
    .A1(\samples_imag[1][3] ),
    .S(_03853_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _12482_ (.A0(net134),
    .A1(\samples_imag[0][1] ),
    .S(_03853_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(net135),
    .A1(\samples_imag[1][4] ),
    .S(_03853_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(net136),
    .A1(\samples_imag[1][5] ),
    .S(_03853_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(net137),
    .A1(\samples_imag[1][6] ),
    .S(_03853_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _12486_ (.A0(net138),
    .A1(\samples_imag[1][7] ),
    .S(_03853_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(net139),
    .A1(\samples_imag[1][8] ),
    .S(_03853_),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(net140),
    .A1(\samples_imag[1][9] ),
    .S(_03853_),
    .X(_00076_));
 sky130_fd_sc_hd__clkbuf_8 _12489_ (.A(_00559_),
    .X(_03854_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(net141),
    .A1(\samples_imag[1][10] ),
    .S(_03854_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(net142),
    .A1(\samples_imag[1][11] ),
    .S(_03854_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(net143),
    .A1(\samples_imag[1][12] ),
    .S(_03854_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(net144),
    .A1(\samples_imag[1][13] ),
    .S(_03854_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _12494_ (.A0(net145),
    .A1(\samples_imag[0][2] ),
    .S(_03854_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(net146),
    .A1(\samples_imag[1][14] ),
    .S(_03854_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(net147),
    .A1(\samples_imag[1][15] ),
    .S(_03854_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(net148),
    .A1(\samples_imag[2][0] ),
    .S(_03854_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(net149),
    .A1(\samples_imag[2][1] ),
    .S(_03854_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(net150),
    .A1(\samples_imag[2][2] ),
    .S(_03854_),
    .X(_00086_));
 sky130_fd_sc_hd__buf_6 _12500_ (.A(_00559_),
    .X(_03855_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(net151),
    .A1(\samples_imag[2][3] ),
    .S(_03855_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _12502_ (.A0(net152),
    .A1(\samples_imag[2][4] ),
    .S(_03855_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _12503_ (.A0(net153),
    .A1(\samples_imag[2][5] ),
    .S(_03855_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(net154),
    .A1(\samples_imag[2][6] ),
    .S(_03855_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(net155),
    .A1(\samples_imag[2][7] ),
    .S(_03855_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(net156),
    .A1(\samples_imag[0][3] ),
    .S(_03855_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _12507_ (.A0(net157),
    .A1(\samples_imag[2][8] ),
    .S(_03855_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _12508_ (.A0(net158),
    .A1(\samples_imag[2][9] ),
    .S(_03855_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(net159),
    .A1(\samples_imag[2][10] ),
    .S(_03855_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(net160),
    .A1(\samples_imag[2][11] ),
    .S(_03855_),
    .X(_00096_));
 sky130_fd_sc_hd__buf_4 _12511_ (.A(_00559_),
    .X(_03856_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(net161),
    .A1(\samples_imag[2][12] ),
    .S(_03856_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(net162),
    .A1(\samples_imag[2][13] ),
    .S(_03856_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(net163),
    .A1(\samples_imag[2][14] ),
    .S(_03856_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(net164),
    .A1(\samples_imag[2][15] ),
    .S(_03856_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(net165),
    .A1(\samples_imag[3][0] ),
    .S(_03856_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(net166),
    .A1(\samples_imag[3][1] ),
    .S(_03856_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(net167),
    .A1(\samples_imag[0][4] ),
    .S(_03856_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(net168),
    .A1(\samples_imag[3][2] ),
    .S(_03856_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(net169),
    .A1(\samples_imag[3][3] ),
    .S(_03856_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _12521_ (.A0(net170),
    .A1(\samples_imag[3][4] ),
    .S(_03856_),
    .X(_00106_));
 sky130_fd_sc_hd__buf_6 _12522_ (.A(_00559_),
    .X(_03857_));
 sky130_fd_sc_hd__mux2_1 _12523_ (.A0(net171),
    .A1(\samples_imag[3][5] ),
    .S(_03857_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(net172),
    .A1(\samples_imag[3][6] ),
    .S(_03857_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(net173),
    .A1(\samples_imag[3][7] ),
    .S(_03857_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _12526_ (.A0(net174),
    .A1(\samples_imag[3][8] ),
    .S(_03857_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _12527_ (.A0(net175),
    .A1(\samples_imag[3][9] ),
    .S(_03857_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _12528_ (.A0(net176),
    .A1(\samples_imag[3][10] ),
    .S(_03857_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _12529_ (.A0(net177),
    .A1(\samples_imag[3][11] ),
    .S(_03857_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _12530_ (.A0(net178),
    .A1(\samples_imag[0][5] ),
    .S(_03857_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _12531_ (.A0(net179),
    .A1(\samples_imag[3][12] ),
    .S(_03857_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _12532_ (.A0(net180),
    .A1(\samples_imag[3][13] ),
    .S(_03857_),
    .X(_00116_));
 sky130_fd_sc_hd__buf_6 _12533_ (.A(_00558_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_4 _12534_ (.A(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(net181),
    .A1(\samples_imag[3][14] ),
    .S(_03859_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _12536_ (.A0(net182),
    .A1(\samples_imag[3][15] ),
    .S(_03859_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(net183),
    .A1(\samples_imag[4][0] ),
    .S(_03859_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(net184),
    .A1(\samples_imag[4][1] ),
    .S(_03859_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(net185),
    .A1(\samples_imag[4][2] ),
    .S(_03859_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _12540_ (.A0(net186),
    .A1(\samples_imag[4][3] ),
    .S(_03859_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(net187),
    .A1(\samples_imag[4][4] ),
    .S(_03859_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _12542_ (.A0(net188),
    .A1(\samples_imag[4][5] ),
    .S(_03859_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(net189),
    .A1(\samples_imag[0][6] ),
    .S(_03859_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(net190),
    .A1(\samples_imag[4][6] ),
    .S(_03859_),
    .X(_00126_));
 sky130_fd_sc_hd__clkbuf_4 _12545_ (.A(_03858_),
    .X(_03860_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(net191),
    .A1(\samples_imag[4][7] ),
    .S(_03860_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(net192),
    .A1(\samples_imag[4][8] ),
    .S(_03860_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(net193),
    .A1(\samples_imag[4][9] ),
    .S(_03860_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(net194),
    .A1(\samples_imag[4][10] ),
    .S(_03860_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(net195),
    .A1(\samples_imag[4][11] ),
    .S(_03860_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(net196),
    .A1(\samples_imag[4][12] ),
    .S(_03860_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(net197),
    .A1(\samples_imag[4][13] ),
    .S(_03860_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(net198),
    .A1(\samples_imag[4][14] ),
    .S(_03860_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(net199),
    .A1(\samples_imag[4][15] ),
    .S(_03860_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(net200),
    .A1(\samples_imag[0][7] ),
    .S(_03860_),
    .X(_00136_));
 sky130_fd_sc_hd__clkbuf_4 _12556_ (.A(_03858_),
    .X(_03861_));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(net201),
    .A1(\samples_imag[5][0] ),
    .S(_03861_),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(net202),
    .A1(\samples_imag[5][1] ),
    .S(_03861_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(net203),
    .A1(\samples_imag[5][2] ),
    .S(_03861_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(net204),
    .A1(\samples_imag[5][3] ),
    .S(_03861_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(net205),
    .A1(\samples_imag[5][4] ),
    .S(_03861_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(net206),
    .A1(\samples_imag[5][5] ),
    .S(_03861_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(net207),
    .A1(\samples_imag[5][6] ),
    .S(_03861_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(net208),
    .A1(\samples_imag[5][7] ),
    .S(_03861_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(net209),
    .A1(\samples_imag[5][8] ),
    .S(_03861_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(net210),
    .A1(\samples_imag[5][9] ),
    .S(_03861_),
    .X(_00146_));
 sky130_fd_sc_hd__buf_4 _12567_ (.A(_03858_),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_1 _12568_ (.A0(net211),
    .A1(\samples_imag[0][8] ),
    .S(_03862_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(net212),
    .A1(\samples_imag[5][10] ),
    .S(_03862_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(net213),
    .A1(\samples_imag[5][11] ),
    .S(_03862_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(net214),
    .A1(\samples_imag[5][12] ),
    .S(_03862_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(net215),
    .A1(\samples_imag[5][13] ),
    .S(_03862_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(net216),
    .A1(\samples_imag[5][14] ),
    .S(_03862_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(net217),
    .A1(\samples_imag[5][15] ),
    .S(_03862_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(net218),
    .A1(\samples_imag[6][0] ),
    .S(_03862_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(net219),
    .A1(\samples_imag[6][1] ),
    .S(_03862_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(net220),
    .A1(\samples_imag[6][2] ),
    .S(_03862_),
    .X(_00156_));
 sky130_fd_sc_hd__buf_4 _12578_ (.A(_03858_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(net221),
    .A1(\samples_imag[6][3] ),
    .S(_03863_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(net222),
    .A1(\samples_imag[0][9] ),
    .S(_03863_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(net223),
    .A1(\samples_real[0][0] ),
    .S(_03863_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(net224),
    .A1(\samples_real[6][4] ),
    .S(_03863_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(net225),
    .A1(\samples_real[6][5] ),
    .S(_03863_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(net226),
    .A1(\samples_real[6][6] ),
    .S(_03863_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(net227),
    .A1(\samples_real[6][7] ),
    .S(_03863_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(net228),
    .A1(\samples_real[6][8] ),
    .S(_03863_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(net229),
    .A1(\samples_real[6][9] ),
    .S(_03863_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(net230),
    .A1(\samples_real[6][10] ),
    .S(_03863_),
    .X(_00166_));
 sky130_fd_sc_hd__buf_4 _12589_ (.A(_03858_),
    .X(_03864_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(net231),
    .A1(\samples_real[6][11] ),
    .S(_03864_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(net232),
    .A1(\samples_real[6][12] ),
    .S(_03864_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(net233),
    .A1(\samples_real[6][13] ),
    .S(_03864_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(net234),
    .A1(\samples_real[0][10] ),
    .S(_03864_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(net235),
    .A1(\samples_real[6][14] ),
    .S(_03864_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(net236),
    .A1(\samples_real[6][15] ),
    .S(_03864_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(net237),
    .A1(\samples_real[7][0] ),
    .S(_03864_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(net238),
    .A1(\samples_real[7][1] ),
    .S(_03864_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(net239),
    .A1(\samples_real[7][2] ),
    .S(_03864_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _12599_ (.A0(net240),
    .A1(\samples_real[7][3] ),
    .S(_03864_),
    .X(_00176_));
 sky130_fd_sc_hd__buf_4 _12600_ (.A(_03858_),
    .X(_03865_));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(net241),
    .A1(\samples_real[7][4] ),
    .S(_03865_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(net242),
    .A1(\samples_real[7][5] ),
    .S(_03865_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(net243),
    .A1(\samples_real[7][6] ),
    .S(_03865_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(net244),
    .A1(\samples_real[7][7] ),
    .S(_03865_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(net245),
    .A1(\samples_real[0][11] ),
    .S(_03865_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(net246),
    .A1(\samples_real[7][8] ),
    .S(_03865_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(net247),
    .A1(\samples_real[7][9] ),
    .S(_03865_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(net248),
    .A1(\samples_real[7][10] ),
    .S(_03865_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(net249),
    .A1(\samples_real[7][11] ),
    .S(_03865_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _12610_ (.A0(net250),
    .A1(\samples_real[7][12] ),
    .S(_03865_),
    .X(_00186_));
 sky130_fd_sc_hd__buf_6 _12611_ (.A(_03858_),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(net251),
    .A1(\samples_real[7][13] ),
    .S(_03866_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _12613_ (.A0(net252),
    .A1(\samples_real[7][14] ),
    .S(_03866_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _12614_ (.A0(net253),
    .A1(\samples_real[7][15] ),
    .S(_03866_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(net254),
    .A1(\samples_real[0][12] ),
    .S(_03866_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _12616_ (.A0(net255),
    .A1(\samples_real[0][13] ),
    .S(_03866_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(net256),
    .A1(\samples_real[0][14] ),
    .S(_03866_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _12618_ (.A0(net257),
    .A1(\samples_real[0][15] ),
    .S(_03866_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(net258),
    .A1(\samples_real[1][0] ),
    .S(_03866_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _12620_ (.A0(net259),
    .A1(\samples_real[1][1] ),
    .S(_03866_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(net260),
    .A1(\samples_real[1][2] ),
    .S(_03866_),
    .X(_00196_));
 sky130_fd_sc_hd__clkbuf_4 _12622_ (.A(_03858_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _12623_ (.A0(net261),
    .A1(\samples_real[1][3] ),
    .S(_03867_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _12624_ (.A0(net262),
    .A1(\samples_real[0][1] ),
    .S(_03867_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(net263),
    .A1(\samples_real[1][4] ),
    .S(_03867_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _12626_ (.A0(net264),
    .A1(\samples_real[1][5] ),
    .S(_03867_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(net265),
    .A1(\samples_real[1][6] ),
    .S(_03867_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _12628_ (.A0(net266),
    .A1(\samples_real[1][7] ),
    .S(_03867_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _12629_ (.A0(net267),
    .A1(\samples_real[1][8] ),
    .S(_03867_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(net268),
    .A1(\samples_real[1][9] ),
    .S(_03867_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(net269),
    .A1(\samples_real[1][10] ),
    .S(_03867_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(net270),
    .A1(\samples_real[1][11] ),
    .S(_03867_),
    .X(_00206_));
 sky130_fd_sc_hd__buf_4 _12633_ (.A(_03858_),
    .X(_03868_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(net271),
    .A1(\samples_real[1][12] ),
    .S(_03868_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _12635_ (.A0(net272),
    .A1(\samples_real[1][13] ),
    .S(_03868_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(net273),
    .A1(\samples_real[0][2] ),
    .S(_03868_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _12637_ (.A0(net274),
    .A1(\samples_real[1][14] ),
    .S(_03868_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(net275),
    .A1(\samples_real[1][15] ),
    .S(_03868_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _12639_ (.A0(net276),
    .A1(\samples_real[2][0] ),
    .S(_03868_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(net277),
    .A1(\samples_real[2][1] ),
    .S(_03868_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(net278),
    .A1(\samples_real[2][2] ),
    .S(_03868_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _12642_ (.A0(net279),
    .A1(\samples_real[2][3] ),
    .S(_03868_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(net280),
    .A1(\samples_real[2][4] ),
    .S(_03868_),
    .X(_00216_));
 sky130_fd_sc_hd__clkbuf_4 _12644_ (.A(_00558_),
    .X(_03869_));
 sky130_fd_sc_hd__mux2_1 _12645_ (.A0(net281),
    .A1(\samples_real[2][5] ),
    .S(_03869_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(net282),
    .A1(\samples_real[2][6] ),
    .S(_03869_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _12647_ (.A0(net283),
    .A1(\samples_real[2][7] ),
    .S(_03869_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(net284),
    .A1(\samples_real[0][3] ),
    .S(_03869_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _12649_ (.A0(net285),
    .A1(\samples_real[2][8] ),
    .S(_03869_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _12650_ (.A0(net286),
    .A1(\samples_real[2][9] ),
    .S(_03869_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _12651_ (.A0(net287),
    .A1(\samples_real[2][10] ),
    .S(_03869_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(net288),
    .A1(\samples_real[2][11] ),
    .S(_03869_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _12653_ (.A0(net289),
    .A1(\samples_real[2][12] ),
    .S(_03869_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(net290),
    .A1(\samples_real[2][13] ),
    .S(_03869_),
    .X(_00226_));
 sky130_fd_sc_hd__buf_4 _12655_ (.A(_00558_),
    .X(_03870_));
 sky130_fd_sc_hd__mux2_1 _12656_ (.A0(net291),
    .A1(\samples_real[2][14] ),
    .S(_03870_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _12657_ (.A0(net292),
    .A1(\samples_real[2][15] ),
    .S(_03870_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(net293),
    .A1(\samples_real[3][0] ),
    .S(_03870_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(net294),
    .A1(\samples_real[3][1] ),
    .S(_03870_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(net295),
    .A1(\samples_real[0][4] ),
    .S(_03870_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(net296),
    .A1(\samples_real[3][2] ),
    .S(_03870_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(net297),
    .A1(\samples_real[3][3] ),
    .S(_03870_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _12663_ (.A0(net298),
    .A1(\samples_real[3][4] ),
    .S(_03870_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _12664_ (.A0(net299),
    .A1(\samples_real[3][5] ),
    .S(_03870_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _12665_ (.A0(net300),
    .A1(\samples_real[3][6] ),
    .S(_03870_),
    .X(_00236_));
 sky130_fd_sc_hd__clkbuf_4 _12666_ (.A(_00558_),
    .X(_03871_));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(net301),
    .A1(\samples_real[3][7] ),
    .S(_03871_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(net302),
    .A1(\samples_real[3][8] ),
    .S(_03871_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _12669_ (.A0(net303),
    .A1(\samples_real[3][9] ),
    .S(_03871_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(net304),
    .A1(\samples_real[3][10] ),
    .S(_03871_),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(net305),
    .A1(\samples_real[3][11] ),
    .S(_03871_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _12672_ (.A0(net306),
    .A1(\samples_real[0][5] ),
    .S(_03871_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(net307),
    .A1(\samples_real[3][12] ),
    .S(_03871_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _12674_ (.A0(net308),
    .A1(\samples_real[3][13] ),
    .S(_03871_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(net309),
    .A1(\samples_real[3][14] ),
    .S(_03871_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _12676_ (.A0(net310),
    .A1(\samples_real[3][15] ),
    .S(_03871_),
    .X(_00246_));
 sky130_fd_sc_hd__buf_4 _12677_ (.A(_00558_),
    .X(_03872_));
 sky130_fd_sc_hd__mux2_1 _12678_ (.A0(net311),
    .A1(\samples_real[4][0] ),
    .S(_03872_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _12679_ (.A0(net312),
    .A1(\samples_real[4][1] ),
    .S(_03872_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _12680_ (.A0(net313),
    .A1(\samples_real[4][2] ),
    .S(_03872_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _12681_ (.A0(net314),
    .A1(\samples_real[4][3] ),
    .S(_03872_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(net315),
    .A1(\samples_real[4][4] ),
    .S(_03872_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(net316),
    .A1(\samples_real[4][5] ),
    .S(_03872_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(net317),
    .A1(\samples_real[0][6] ),
    .S(_03872_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(net318),
    .A1(\samples_real[4][6] ),
    .S(_03872_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(net319),
    .A1(\samples_real[4][7] ),
    .S(_03872_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _12687_ (.A0(net320),
    .A1(\samples_real[4][8] ),
    .S(_03872_),
    .X(_00256_));
 sky130_fd_sc_hd__clkbuf_4 _12688_ (.A(_00558_),
    .X(_03873_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(net321),
    .A1(\samples_real[4][9] ),
    .S(_03873_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(net322),
    .A1(\samples_real[4][10] ),
    .S(_03873_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(net323),
    .A1(\samples_real[4][11] ),
    .S(_03873_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(net324),
    .A1(\samples_real[4][12] ),
    .S(_03873_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(net325),
    .A1(\samples_real[4][13] ),
    .S(_03873_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(net326),
    .A1(\samples_real[4][14] ),
    .S(_03873_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(net327),
    .A1(\samples_real[4][15] ),
    .S(_03873_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(net328),
    .A1(\samples_real[0][7] ),
    .S(_03873_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(net329),
    .A1(\samples_real[5][0] ),
    .S(_03873_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(net330),
    .A1(\samples_real[5][1] ),
    .S(_03873_),
    .X(_00266_));
 sky130_fd_sc_hd__clkbuf_4 _12699_ (.A(_00558_),
    .X(_03874_));
 sky130_fd_sc_hd__mux2_1 _12700_ (.A0(net331),
    .A1(\samples_real[5][2] ),
    .S(_03874_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(net332),
    .A1(\samples_real[5][3] ),
    .S(_03874_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _12702_ (.A0(net333),
    .A1(\samples_real[5][4] ),
    .S(_03874_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(net334),
    .A1(\samples_real[5][5] ),
    .S(_03874_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _12704_ (.A0(net335),
    .A1(\samples_real[5][6] ),
    .S(_03874_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(net336),
    .A1(\samples_real[5][7] ),
    .S(_03874_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(net337),
    .A1(\samples_real[5][8] ),
    .S(_03874_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(net338),
    .A1(\samples_real[5][9] ),
    .S(_03874_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _12708_ (.A0(net339),
    .A1(\samples_real[0][8] ),
    .S(_03874_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(net340),
    .A1(\samples_real[5][10] ),
    .S(_03874_),
    .X(_00276_));
 sky130_fd_sc_hd__buf_4 _12710_ (.A(_00558_),
    .X(_03875_));
 sky130_fd_sc_hd__mux2_1 _12711_ (.A0(net341),
    .A1(\samples_real[5][11] ),
    .S(_03875_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(net342),
    .A1(\samples_real[5][12] ),
    .S(_03875_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(net343),
    .A1(\samples_real[5][13] ),
    .S(_03875_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(net344),
    .A1(\samples_real[5][14] ),
    .S(_03875_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(net345),
    .A1(\samples_real[5][15] ),
    .S(_03875_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(net346),
    .A1(\samples_real[6][0] ),
    .S(_03875_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(net347),
    .A1(\samples_real[6][1] ),
    .S(_03875_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(net348),
    .A1(\samples_real[6][2] ),
    .S(_03875_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _12719_ (.A0(net349),
    .A1(\samples_real[6][3] ),
    .S(_03875_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(net350),
    .A1(\samples_real[0][9] ),
    .S(_03875_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2i_1 _12721_ (.A0(_03140_),
    .A1(net351),
    .S(_00557_),
    .Y(_03876_));
 sky130_fd_sc_hd__a21oi_1 _12722_ (.A1(_03136_),
    .A2(_00560_),
    .B1(net351),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _12723_ (.A(net351),
    .B(_03138_),
    .Y(_03878_));
 sky130_fd_sc_hd__o221ai_1 _12724_ (.A1(_03136_),
    .A2(_03876_),
    .B1(_03877_),
    .B2(_03137_),
    .C1(_03878_),
    .Y(_00287_));
 sky130_fd_sc_hd__o21bai_1 _12725_ (.A1(net93),
    .A2(net352),
    .B1_N(_03842_),
    .Y(_03879_));
 sky130_fd_sc_hd__nor2_1 _12726_ (.A(_00560_),
    .B(net352),
    .Y(_03880_));
 sky130_fd_sc_hd__a21oi_1 _12727_ (.A1(\state[0] ),
    .A2(_03879_),
    .B1(_03880_),
    .Y(_00288_));
 sky130_fd_sc_hd__nor2_1 _12728_ (.A(_03140_),
    .B(net91),
    .Y(_03881_));
 sky130_fd_sc_hd__o21ai_0 _12729_ (.A1(_03136_),
    .A2(net93),
    .B1(_03143_),
    .Y(_03882_));
 sky130_fd_sc_hd__a211oi_2 _12730_ (.A1(_03136_),
    .A2(_03845_),
    .B1(_03881_),
    .C1(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__nand4b_1 _12731_ (.A_N(_07833_),
    .B(_07827_),
    .C(_03883_),
    .D(_03137_),
    .Y(_03884_));
 sky130_fd_sc_hd__o21ai_0 _12732_ (.A1(_07827_),
    .A2(_03883_),
    .B1(_03884_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand4b_1 _12733_ (.A_N(_07833_),
    .B(_07830_),
    .C(_03883_),
    .D(_03137_),
    .Y(_03885_));
 sky130_fd_sc_hd__o21ai_0 _12734_ (.A1(_07828_),
    .A2(_03883_),
    .B1(_03885_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand3_1 _12735_ (.A(_03137_),
    .B(_07834_),
    .C(_03883_),
    .Y(_03886_));
 sky130_fd_sc_hd__o21ai_0 _12736_ (.A1(_03833_),
    .A2(_03883_),
    .B1(_03886_),
    .Y(_00291_));
 sky130_fd_sc_hd__nor2b_2 _12737_ (.A(\sample_count[2] ),
    .B_N(_07829_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2b_4 _12738_ (.A_N(_03887_),
    .B(_03137_),
    .Y(_03888_));
 sky130_fd_sc_hd__nor3_1 _12739_ (.A(_03837_),
    .B(_03835_),
    .C(_03839_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2b_1 _12740_ (.A_N(\butterfly_count[2] ),
    .B(_07819_),
    .Y(_03890_));
 sky130_fd_sc_hd__a211oi_4 _12741_ (.A1(\state[1] ),
    .A2(_03890_),
    .B1(_03881_),
    .C1(_03845_),
    .Y(_03891_));
 sky130_fd_sc_hd__o21ai_4 _12742_ (.A1(_03888_),
    .A2(_03889_),
    .B1(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__buf_2 _12743_ (.A(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__clkbuf_4 _12744_ (.A(_03309_),
    .X(_03894_));
 sky130_fd_sc_hd__xnor2_4 _12745_ (.A(\temp_imag[0] ),
    .B(_07850_),
    .Y(_03895_));
 sky130_fd_sc_hd__clkbuf_2 _12746_ (.A(_07842_),
    .X(_03896_));
 sky130_fd_sc_hd__inv_1 _12747_ (.A(_07856_),
    .Y(_03897_));
 sky130_fd_sc_hd__clkbuf_2 _12748_ (.A(_07861_),
    .X(_03898_));
 sky130_fd_sc_hd__inv_1 _12749_ (.A(_07866_),
    .Y(_03899_));
 sky130_fd_sc_hd__clkbuf_2 _12750_ (.A(_07871_),
    .X(_03900_));
 sky130_fd_sc_hd__inv_1 _12751_ (.A(_07876_),
    .Y(_03901_));
 sky130_fd_sc_hd__clkbuf_2 _12752_ (.A(_07881_),
    .X(_03902_));
 sky130_fd_sc_hd__inv_1 _12753_ (.A(_07886_),
    .Y(_03903_));
 sky130_fd_sc_hd__clkbuf_2 _12754_ (.A(_07891_),
    .X(_03904_));
 sky130_fd_sc_hd__clkbuf_2 _12755_ (.A(_07896_),
    .X(_03905_));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer167 (.A(_03156_),
    .X(net534));
 sky130_fd_sc_hd__buf_6 _12757_ (.A(_07906_),
    .X(_03907_));
 sky130_fd_sc_hd__a21o_1 _12758_ (.A1(_05903_),
    .A2(_07910_),
    .B1(_07909_),
    .X(_03908_));
 sky130_fd_sc_hd__a21o_1 _12759_ (.A1(_03908_),
    .A2(_03907_),
    .B1(_07905_),
    .X(_03909_));
 sky130_fd_sc_hd__a21o_1 _12760_ (.A1(_03909_),
    .A2(_07901_),
    .B1(_07900_),
    .X(_03910_));
 sky130_fd_sc_hd__a21o_1 _12761_ (.A1(_03910_),
    .A2(_03905_),
    .B1(_07895_),
    .X(_03911_));
 sky130_fd_sc_hd__a21oi_2 _12762_ (.A1(_03911_),
    .A2(_03904_),
    .B1(_07890_),
    .Y(_03912_));
 sky130_fd_sc_hd__o21bai_2 _12763_ (.A1(_03912_),
    .A2(_03903_),
    .B1_N(_07885_),
    .Y(_03913_));
 sky130_fd_sc_hd__a21oi_2 _12764_ (.A1(_03913_),
    .A2(_03902_),
    .B1(_07880_),
    .Y(_03914_));
 sky130_fd_sc_hd__o21bai_2 _12765_ (.A1(_03914_),
    .A2(_03901_),
    .B1_N(_07875_),
    .Y(_03915_));
 sky130_fd_sc_hd__a21oi_2 _12766_ (.A1(_03915_),
    .A2(_03900_),
    .B1(_07870_),
    .Y(_03916_));
 sky130_fd_sc_hd__o21bai_2 _12767_ (.A1(_03916_),
    .A2(_03899_),
    .B1_N(_07865_),
    .Y(_03917_));
 sky130_fd_sc_hd__a21oi_2 _12768_ (.A1(_03917_),
    .A2(_03898_),
    .B1(_07860_),
    .Y(_03918_));
 sky130_fd_sc_hd__o21bai_2 _12769_ (.A1(_03918_),
    .A2(_03897_),
    .B1_N(_07855_),
    .Y(_03919_));
 sky130_fd_sc_hd__a21o_1 _12770_ (.A1(_03919_),
    .A2(_03896_),
    .B1(_07841_),
    .X(_03920_));
 sky130_fd_sc_hd__a21oi_4 _12771_ (.A1(_07837_),
    .A2(_03920_),
    .B1(_07836_),
    .Y(_03921_));
 sky130_fd_sc_hd__xnor2_4 _12772_ (.A(_03895_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__and3_4 _12773_ (.A(\temp_imag[0] ),
    .B(_07853_),
    .C(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__xnor2_4 clone54 (.A(net523),
    .B(_03895_),
    .Y(net54));
 sky130_fd_sc_hd__nand2b_4 _12775_ (.A_N(_03923_),
    .B(_07847_),
    .Y(_03925_));
 sky130_fd_sc_hd__buf_1 rebuffer164 (.A(_03921_),
    .X(net531));
 sky130_fd_sc_hd__inv_1 _12777_ (.A(_07910_),
    .Y(_03927_));
 sky130_fd_sc_hd__a21oi_1 _12778_ (.A1(_03927_),
    .A2(_07845_),
    .B1(_07911_),
    .Y(_03928_));
 sky130_fd_sc_hd__nor2_1 _12779_ (.A(_03907_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nor2_1 _12780_ (.A(_07907_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__nor2_1 _12781_ (.A(_07901_),
    .B(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__nor2_1 _12782_ (.A(_07902_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__nor2_1 _12783_ (.A(_03905_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__nor2_1 _12784_ (.A(_07897_),
    .B(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__o21bai_1 _12785_ (.A1(_03904_),
    .A2(_03934_),
    .B1_N(_07892_),
    .Y(_03935_));
 sky130_fd_sc_hd__a21oi_2 _12786_ (.A1(_03903_),
    .A2(_03935_),
    .B1(_07887_),
    .Y(_03936_));
 sky130_fd_sc_hd__o21bai_1 _12787_ (.A1(_03902_),
    .A2(_03936_),
    .B1_N(_07882_),
    .Y(_03937_));
 sky130_fd_sc_hd__a21oi_2 _12788_ (.A1(_03937_),
    .A2(_03901_),
    .B1(_07877_),
    .Y(_03938_));
 sky130_fd_sc_hd__o21bai_1 _12789_ (.A1(_03900_),
    .A2(_03938_),
    .B1_N(_07872_),
    .Y(_03939_));
 sky130_fd_sc_hd__a21oi_2 _12790_ (.A1(_03939_),
    .A2(_03899_),
    .B1(_07867_),
    .Y(_03940_));
 sky130_fd_sc_hd__o21bai_1 _12791_ (.A1(_03898_),
    .A2(_03940_),
    .B1_N(_07862_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21oi_2 _12792_ (.A1(_03897_),
    .A2(_03941_),
    .B1(_07857_),
    .Y(_03942_));
 sky130_fd_sc_hd__nor2_1 _12793_ (.A(_03896_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__nor2_1 _12794_ (.A(_07843_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__nor2_1 _12795_ (.A(_07837_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__nor2_1 _12796_ (.A(_03945_),
    .B(_07838_),
    .Y(_03946_));
 sky130_fd_sc_hd__xor2_2 _12797_ (.A(_03895_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__nor2_1 _12798_ (.A(_03907_),
    .B(_05900_),
    .Y(_03948_));
 sky130_fd_sc_hd__nor2_1 _12799_ (.A(_07907_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__nor2_1 _12800_ (.A(_07901_),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__nor2_1 _12801_ (.A(_03950_),
    .B(_07902_),
    .Y(_03951_));
 sky130_fd_sc_hd__nor2_1 _12802_ (.A(_03905_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__nor2_1 _12803_ (.A(_07897_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__nor2_1 _12804_ (.A(_03904_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__nor2_1 _12805_ (.A(_03954_),
    .B(_07892_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_1 _12806_ (.A(_07886_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__nor2_1 _12807_ (.A(_07887_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__nor2_2 _12808_ (.A(_03957_),
    .B(_03902_),
    .Y(_03958_));
 sky130_fd_sc_hd__nor2_2 _12809_ (.A(_07882_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nor2_1 _12810_ (.A(_07876_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nor2_1 _12811_ (.A(_07877_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__nor2_1 _12812_ (.A(_03900_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__nor2_1 _12813_ (.A(_03962_),
    .B(_07872_),
    .Y(_03963_));
 sky130_fd_sc_hd__nor2_1 _12814_ (.A(_07866_),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__nor2_1 _12815_ (.A(_07867_),
    .B(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hd__nor2_1 _12816_ (.A(_03898_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__nor2_1 _12817_ (.A(_07862_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__nor2_1 _12818_ (.A(_07856_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__nor2_1 _12819_ (.A(_07857_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__nor2_1 _12820_ (.A(_03896_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__nor2_1 _12821_ (.A(_07843_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__xnor2_1 _12822_ (.A(_03971_),
    .B(_07837_),
    .Y(_03972_));
 sky130_fd_sc_hd__xnor2_1 _12823_ (.A(_03896_),
    .B(_03942_),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_1 _12824_ (.A(_07856_),
    .B(net616),
    .Y(_03974_));
 sky130_fd_sc_hd__xnor2_1 _12825_ (.A(_07886_),
    .B(net557),
    .Y(_03975_));
 sky130_fd_sc_hd__xnor2_1 _12826_ (.A(_03904_),
    .B(net638),
    .Y(_03976_));
 sky130_fd_sc_hd__xnor2_1 _12827_ (.A(_07901_),
    .B(net644),
    .Y(_03977_));
 sky130_fd_sc_hd__xnor2_1 _12828_ (.A(_03907_),
    .B(_05900_),
    .Y(_03978_));
 sky130_fd_sc_hd__xnor2_1 _12829_ (.A(_03905_),
    .B(net554),
    .Y(_03979_));
 sky130_fd_sc_hd__and4b_1 _12830_ (.A_N(_07847_),
    .B(_03978_),
    .C(_03979_),
    .D(_05901_),
    .X(_03980_));
 sky130_fd_sc_hd__nand4_1 _12831_ (.A(_03975_),
    .B(_03976_),
    .C(_03977_),
    .D(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__xnor2_1 _12832_ (.A(_07876_),
    .B(net641),
    .Y(_03982_));
 sky130_fd_sc_hd__xnor2_1 _12833_ (.A(_03902_),
    .B(_03936_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _12834_ (.A(_03982_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__nor2_1 _12835_ (.A(_03981_),
    .B(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__xnor2_1 _12836_ (.A(_03900_),
    .B(_03938_),
    .Y(_03986_));
 sky130_fd_sc_hd__xnor2_1 _12837_ (.A(_07866_),
    .B(net563),
    .Y(_03987_));
 sky130_fd_sc_hd__xnor2_1 _12838_ (.A(_03898_),
    .B(_03940_),
    .Y(_03988_));
 sky130_fd_sc_hd__and4_1 _12839_ (.A(_03985_),
    .B(_03986_),
    .C(_03987_),
    .D(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__nand4_2 _12840_ (.A(_03989_),
    .B(_03973_),
    .C(_03974_),
    .D(_03972_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand3_4 _12841_ (.A(\temp_imag[0] ),
    .B(_03990_),
    .C(_07852_),
    .Y(_03991_));
 sky130_fd_sc_hd__nor2_8 _12842_ (.A(_03947_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__nor2b_4 _12843_ (.A(_03992_),
    .B_N(_07847_),
    .Y(_03993_));
 sky130_fd_sc_hd__buf_6 _12844_ (.A(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__nor2_1 _12845_ (.A(_03176_),
    .B(_03892_),
    .Y(_03995_));
 sky130_fd_sc_hd__a22o_1 _12846_ (.A1(\samples_imag[0][0] ),
    .A2(_03176_),
    .B1(_03994_),
    .B2(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(_03449_),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__o31ai_2 _12848_ (.A1(_03894_),
    .A2(_03893_),
    .A3(_03925_),
    .B1(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__buf_6 _12849_ (.A(_03142_),
    .X(_03999_));
 sky130_fd_sc_hd__nand2b_1 _12850_ (.A_N(_03141_),
    .B(net34),
    .Y(_04000_));
 sky130_fd_sc_hd__buf_4 _12851_ (.A(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__nor2_1 _12852_ (.A(_03893_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__a221o_1 _12853_ (.A1(\samples_imag[0][0] ),
    .A2(_03893_),
    .B1(_03998_),
    .B2(_03999_),
    .C1(_04002_),
    .X(_00292_));
 sky130_fd_sc_hd__clkbuf_4 _12854_ (.A(_03893_),
    .X(_04003_));
 sky130_fd_sc_hd__buf_6 _12855_ (.A(_03142_),
    .X(_04004_));
 sky130_fd_sc_hd__buf_6 _12856_ (.A(_03992_),
    .X(_04005_));
 sky130_fd_sc_hd__or2_4 _12857_ (.A(_04005_),
    .B(_03987_),
    .X(_04006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__nor2_1 _12859_ (.A(_03177_),
    .B(_04006_),
    .Y(_04008_));
 sky130_fd_sc_hd__a21oi_1 _12860_ (.A1(\samples_imag[0][10] ),
    .A2(_03207_),
    .B1(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__buf_12 _12861_ (.A(_03923_),
    .X(_04010_));
 sky130_fd_sc_hd__a21o_1 _12862_ (.A1(_03907_),
    .A2(_05904_),
    .B1(_07905_),
    .X(_04011_));
 sky130_fd_sc_hd__a21o_1 _12863_ (.A1(_07901_),
    .A2(_04011_),
    .B1(_07900_),
    .X(_04012_));
 sky130_fd_sc_hd__a21o_1 _12864_ (.A1(_03905_),
    .A2(_04012_),
    .B1(_07895_),
    .X(_04013_));
 sky130_fd_sc_hd__a21oi_2 _12865_ (.A1(_03904_),
    .A2(_04013_),
    .B1(_07890_),
    .Y(_04014_));
 sky130_fd_sc_hd__o21bai_1 _12866_ (.A1(_03903_),
    .A2(_04014_),
    .B1_N(_07885_),
    .Y(_04015_));
 sky130_fd_sc_hd__a21oi_2 _12867_ (.A1(_04015_),
    .A2(_03902_),
    .B1(_07880_),
    .Y(_04016_));
 sky130_fd_sc_hd__o21bai_1 _12868_ (.A1(_03901_),
    .A2(_04016_),
    .B1_N(_07875_),
    .Y(_04017_));
 sky130_fd_sc_hd__a21oi_2 _12869_ (.A1(_03900_),
    .A2(_04017_),
    .B1(_07870_),
    .Y(_04018_));
 sky130_fd_sc_hd__xnor2_2 _12870_ (.A(_03899_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__nor2_8 _12871_ (.A(net62),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__nor2_1 _12872_ (.A(_03314_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21oi_1 _12873_ (.A1(_04009_),
    .A2(_03310_),
    .B1(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__buf_2 _12874_ (.A(\state[1] ),
    .X(_04023_));
 sky130_fd_sc_hd__nor2b_1 _12875_ (.A(_04023_),
    .B_N(net40),
    .Y(_04024_));
 sky130_fd_sc_hd__buf_4 _12876_ (.A(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__a21oi_1 _12877_ (.A1(_04004_),
    .A2(_04022_),
    .B1(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__buf_2 _12878_ (.A(_03893_),
    .X(_04027_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(\samples_imag[0][10] ),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__o21ai_1 _12880_ (.A1(_04003_),
    .A2(_04026_),
    .B1(_04028_),
    .Y(_00293_));
 sky130_fd_sc_hd__buf_4 _12881_ (.A(_03142_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_4 _12882_ (.A(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__or2_4 _12883_ (.A(_04005_),
    .B(_03988_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_4 clone66 (.A(net605),
    .X(net66));
 sky130_fd_sc_hd__nor2_2 _12885_ (.A(_03177_),
    .B(_04031_),
    .Y(_04033_));
 sky130_fd_sc_hd__a21oi_1 _12886_ (.A1(\samples_imag[0][11] ),
    .A2(_03207_),
    .B1(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__xnor2_2 _12887_ (.A(_03898_),
    .B(net543),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_8 _12888_ (.A(_04035_),
    .B(_04010_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_1 _12889_ (.A(_03314_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__a21oi_1 _12890_ (.A1(_04034_),
    .A2(_03310_),
    .B1(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__nor2b_1 _12891_ (.A(_04023_),
    .B_N(net47),
    .Y(_04039_));
 sky130_fd_sc_hd__buf_4 _12892_ (.A(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__a21oi_1 _12893_ (.A1(_04030_),
    .A2(_04038_),
    .B1(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_1 _12894_ (.A(\samples_imag[0][11] ),
    .B(_04027_),
    .Y(_04042_));
 sky130_fd_sc_hd__o21ai_1 _12895_ (.A1(_04003_),
    .A2(_04041_),
    .B1(_04042_),
    .Y(_00294_));
 sky130_fd_sc_hd__buf_2 _12896_ (.A(_03892_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_4 _12897_ (.A(_03176_),
    .X(_04044_));
 sky130_fd_sc_hd__or2_4 _12898_ (.A(net77),
    .B(_03974_),
    .X(_04045_));
 sky130_fd_sc_hd__buf_6 clone55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__nor2_1 _12900_ (.A(_04044_),
    .B(_04045_),
    .Y(_04047_));
 sky130_fd_sc_hd__a21oi_1 _12901_ (.A1(\samples_imag[0][12] ),
    .A2(_03207_),
    .B1(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__o21bai_1 _12902_ (.A1(_03899_),
    .A2(_04018_),
    .B1_N(_07865_),
    .Y(_04049_));
 sky130_fd_sc_hd__a21oi_2 _12903_ (.A1(_03898_),
    .A2(_04049_),
    .B1(_07860_),
    .Y(_04050_));
 sky130_fd_sc_hd__xnor2_2 _12904_ (.A(_03897_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__nor2_8 _12905_ (.A(_04051_),
    .B(_04010_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor2_1 _12906_ (.A(_03314_),
    .B(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__a21oi_1 _12907_ (.A1(_04048_),
    .A2(_03310_),
    .B1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__clkbuf_4 _12908_ (.A(\state[1] ),
    .X(_04055_));
 sky130_fd_sc_hd__nor2b_1 _12909_ (.A(_04055_),
    .B_N(net48),
    .Y(_04056_));
 sky130_fd_sc_hd__buf_6 _12910_ (.A(_04056_),
    .X(_04057_));
 sky130_fd_sc_hd__a21oi_1 _12911_ (.A1(_04054_),
    .A2(_04030_),
    .B1(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand2_1 _12912_ (.A(\samples_imag[0][12] ),
    .B(_04027_),
    .Y(_04059_));
 sky130_fd_sc_hd__o21ai_1 _12913_ (.A1(_04043_),
    .A2(_04058_),
    .B1(_04059_),
    .Y(_00295_));
 sky130_fd_sc_hd__clkbuf_4 _12914_ (.A(_03176_),
    .X(_04060_));
 sky130_fd_sc_hd__or2_4 _12915_ (.A(net77),
    .B(_03973_),
    .X(_04061_));
 sky130_fd_sc_hd__buf_8 clone65 (.A(net526),
    .X(net65));
 sky130_fd_sc_hd__nor2_1 _12917_ (.A(_04044_),
    .B(_04061_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21oi_1 _12918_ (.A1(\samples_imag[0][13] ),
    .A2(_04060_),
    .B1(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__xnor2_2 _12919_ (.A(_03896_),
    .B(_03919_),
    .Y(_04065_));
 sky130_fd_sc_hd__nor2_8 _12920_ (.A(_04065_),
    .B(_04010_),
    .Y(_04066_));
 sky130_fd_sc_hd__nor2_1 _12921_ (.A(_03314_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a21oi_1 _12922_ (.A1(_04064_),
    .A2(_03310_),
    .B1(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2b_1 _12923_ (.A(_04023_),
    .B_N(net57),
    .Y(_04069_));
 sky130_fd_sc_hd__buf_6 _12924_ (.A(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__a21oi_1 _12925_ (.A1(_04030_),
    .A2(_04068_),
    .B1(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _12926_ (.A(\samples_imag[0][13] ),
    .B(_04027_),
    .Y(_04072_));
 sky130_fd_sc_hd__o21ai_1 _12927_ (.A1(_04043_),
    .A2(_04071_),
    .B1(_04072_),
    .Y(_00296_));
 sky130_fd_sc_hd__or2_4 _12928_ (.A(net77),
    .B(_03972_),
    .X(_04073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__nor2_2 _12930_ (.A(_04073_),
    .B(_04044_),
    .Y(_04075_));
 sky130_fd_sc_hd__a21oi_1 _12931_ (.A1(\samples_imag[0][14] ),
    .A2(_04060_),
    .B1(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__o21bai_1 _12932_ (.A1(_03897_),
    .A2(_04050_),
    .B1_N(_07855_),
    .Y(_04077_));
 sky130_fd_sc_hd__a21oi_2 _12933_ (.A1(_03896_),
    .A2(_04077_),
    .B1(_07841_),
    .Y(_04078_));
 sky130_fd_sc_hd__xor2_2 _12934_ (.A(_04078_),
    .B(_07837_),
    .X(_04079_));
 sky130_fd_sc_hd__nor2_8 _12935_ (.A(net62),
    .B(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__nor2_1 _12936_ (.A(_03314_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21oi_1 _12937_ (.A1(_04076_),
    .A2(_03310_),
    .B1(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__nor2b_1 _12938_ (.A(_04023_),
    .B_N(net58),
    .Y(_04083_));
 sky130_fd_sc_hd__buf_4 _12939_ (.A(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__a21oi_1 _12940_ (.A1(_04082_),
    .A2(_04030_),
    .B1(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _12941_ (.A(\samples_imag[0][14] ),
    .B(_04027_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21ai_1 _12942_ (.A1(_04085_),
    .A2(_04043_),
    .B1(_04086_),
    .Y(_00297_));
 sky130_fd_sc_hd__clkbuf_4 _12943_ (.A(_03893_),
    .X(_04087_));
 sky130_fd_sc_hd__buf_4 _12944_ (.A(_03142_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_4 _12945_ (.A(_03176_),
    .X(_04089_));
 sky130_fd_sc_hd__a31oi_4 _12946_ (.A1(\temp_imag[0] ),
    .A2(_07852_),
    .A3(net542),
    .B1(net545),
    .Y(_04090_));
 sky130_fd_sc_hd__clkbuf_4 _12947_ (.A(_03176_),
    .X(_04091_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(\samples_imag[0][15] ),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__o211ai_1 _12949_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_04092_),
    .C1(_03309_),
    .Y(_04093_));
 sky130_fd_sc_hd__o21ai_0 _12950_ (.A1(_03894_),
    .A2(net524),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__nor2_4 _12951_ (.A(_03142_),
    .B(net59),
    .Y(_04095_));
 sky130_fd_sc_hd__a211oi_1 _12952_ (.A1(_04088_),
    .A2(_04094_),
    .B1(_04095_),
    .C1(_04087_),
    .Y(_04096_));
 sky130_fd_sc_hd__a21o_1 _12953_ (.A1(\samples_imag[0][15] ),
    .A2(_04087_),
    .B1(_04096_),
    .X(_00298_));
 sky130_fd_sc_hd__or2_4 _12954_ (.A(net77),
    .B(_05901_),
    .X(_04097_));
 sky130_fd_sc_hd__buf_12 clone62 (.A(_03923_),
    .X(net62));
 sky130_fd_sc_hd__nor2_2 _12956_ (.A(_04044_),
    .B(net647),
    .Y(_04099_));
 sky130_fd_sc_hd__a21oi_1 _12957_ (.A1(\samples_imag[0][1] ),
    .A2(_04060_),
    .B1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__nor2_8 _12958_ (.A(_04010_),
    .B(_05905_),
    .Y(_04101_));
 sky130_fd_sc_hd__nor2_1 _12959_ (.A(_03314_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__a21oi_1 _12960_ (.A1(_04100_),
    .A2(_03310_),
    .B1(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nor2b_1 _12961_ (.A(_04055_),
    .B_N(net60),
    .Y(_04104_));
 sky130_fd_sc_hd__clkbuf_8 _12962_ (.A(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__a21oi_1 _12963_ (.A1(_04030_),
    .A2(_04103_),
    .B1(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_1 _12964_ (.A(\samples_imag[0][1] ),
    .B(_04027_),
    .Y(_04107_));
 sky130_fd_sc_hd__o21ai_1 _12965_ (.A1(_04043_),
    .A2(_04106_),
    .B1(_04107_),
    .Y(_00299_));
 sky130_fd_sc_hd__clkbuf_4 _12966_ (.A(_03309_),
    .X(_04108_));
 sky130_fd_sc_hd__or2_4 _12967_ (.A(_03978_),
    .B(_04005_),
    .X(_04109_));
 sky130_fd_sc_hd__buf_6 clone77 (.A(_03992_),
    .X(net77));
 sky130_fd_sc_hd__nor2_1 _12969_ (.A(_04044_),
    .B(_04109_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21oi_1 _12970_ (.A1(\samples_imag[0][2] ),
    .A2(_04060_),
    .B1(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_2 _12971_ (.A(_03907_),
    .B(_05904_),
    .Y(_04113_));
 sky130_fd_sc_hd__nor2_8 _12972_ (.A(_04113_),
    .B(net62),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _12973_ (.A(_03314_),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__a21oi_1 _12974_ (.A1(_04112_),
    .A2(_04108_),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nor2b_1 _12975_ (.A(_04023_),
    .B_N(net61),
    .Y(_04117_));
 sky130_fd_sc_hd__buf_6 _12976_ (.A(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_1 _12977_ (.A1(_04116_),
    .A2(_04030_),
    .B1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _12978_ (.A(\samples_imag[0][2] ),
    .B(_04027_),
    .Y(_04120_));
 sky130_fd_sc_hd__o21ai_1 _12979_ (.A1(_04043_),
    .A2(_04119_),
    .B1(_04120_),
    .Y(_00300_));
 sky130_fd_sc_hd__or2_4 _12980_ (.A(net77),
    .B(_03977_),
    .X(_04121_));
 sky130_fd_sc_hd__dlymetal6s2s_1 split67 (.A(net528),
    .X(net67));
 sky130_fd_sc_hd__nor2_1 _12982_ (.A(_04044_),
    .B(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__a21oi_1 _12983_ (.A1(\samples_imag[0][3] ),
    .A2(_04060_),
    .B1(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_2 _12984_ (.A(_07901_),
    .B(net544),
    .Y(_04125_));
 sky130_fd_sc_hd__nor2_8 _12985_ (.A(_04125_),
    .B(_04010_),
    .Y(_04126_));
 sky130_fd_sc_hd__nor2_1 _12986_ (.A(_03314_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__a21oi_1 _12987_ (.A1(_04124_),
    .A2(_04108_),
    .B1(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__nor2b_1 _12988_ (.A(_04055_),
    .B_N(net63),
    .Y(_04129_));
 sky130_fd_sc_hd__buf_6 _12989_ (.A(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__a21oi_1 _12990_ (.A1(_04030_),
    .A2(_04128_),
    .B1(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _12991_ (.A(\samples_imag[0][3] ),
    .B(_04027_),
    .Y(_04132_));
 sky130_fd_sc_hd__o21ai_1 _12992_ (.A1(_04043_),
    .A2(_04131_),
    .B1(_04132_),
    .Y(_00301_));
 sky130_fd_sc_hd__or2_4 _12993_ (.A(_04005_),
    .B(_03979_),
    .X(_04133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__nor2_1 _12995_ (.A(_04044_),
    .B(_04133_),
    .Y(_04135_));
 sky130_fd_sc_hd__a21oi_1 _12996_ (.A1(\samples_imag[0][4] ),
    .A2(_04060_),
    .B1(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__xnor2_2 _12997_ (.A(_03905_),
    .B(_04012_),
    .Y(_04137_));
 sky130_fd_sc_hd__nor2_8 _12998_ (.A(net62),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__nor2_1 _12999_ (.A(_03314_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__a21oi_1 _13000_ (.A1(_04136_),
    .A2(_04108_),
    .B1(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__nor2b_1 _13001_ (.A(_04023_),
    .B_N(net68),
    .Y(_04141_));
 sky130_fd_sc_hd__buf_4 _13002_ (.A(_04141_),
    .X(_04142_));
 sky130_fd_sc_hd__a21oi_1 _13003_ (.A1(_04030_),
    .A2(_04140_),
    .B1(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand2_1 _13004_ (.A(\samples_imag[0][4] ),
    .B(_04027_),
    .Y(_04144_));
 sky130_fd_sc_hd__o21ai_1 _13005_ (.A1(_04043_),
    .A2(_04143_),
    .B1(_04144_),
    .Y(_00302_));
 sky130_fd_sc_hd__or2_4 _13006_ (.A(_04005_),
    .B(_03976_),
    .X(_04145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__nor2_1 _13008_ (.A(_04145_),
    .B(_04044_),
    .Y(_04147_));
 sky130_fd_sc_hd__a21oi_1 _13009_ (.A1(\samples_imag[0][5] ),
    .A2(_04060_),
    .B1(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__xnor2_2 _13010_ (.A(_03904_),
    .B(_03911_),
    .Y(_04149_));
 sky130_fd_sc_hd__nor2_8 _13011_ (.A(net62),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__nor2_1 _13012_ (.A(_03894_),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__a21oi_1 _13013_ (.A1(_04108_),
    .A2(_04148_),
    .B1(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nor2b_1 _13014_ (.A(_04023_),
    .B_N(net69),
    .Y(_04153_));
 sky130_fd_sc_hd__clkbuf_8 _13015_ (.A(_04153_),
    .X(_04154_));
 sky130_fd_sc_hd__a21oi_2 _13016_ (.A1(_04152_),
    .A2(_04030_),
    .B1(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _13017_ (.A(\samples_imag[0][5] ),
    .B(_04027_),
    .Y(_04156_));
 sky130_fd_sc_hd__o21ai_1 _13018_ (.A1(_04043_),
    .A2(_04155_),
    .B1(_04156_),
    .Y(_00303_));
 sky130_fd_sc_hd__or2_1 _13019_ (.A(_03975_),
    .B(_03992_),
    .X(_04157_));
 sky130_fd_sc_hd__buf_6 _13020_ (.A(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__nor2_1 _13021_ (.A(_04044_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__a21oi_1 _13022_ (.A1(\samples_imag[0][6] ),
    .A2(_04060_),
    .B1(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__xnor2_2 _13023_ (.A(_03903_),
    .B(_04014_),
    .Y(_04161_));
 sky130_fd_sc_hd__nor2_8 _13024_ (.A(net518),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__nor2_1 _13025_ (.A(_03894_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_1 _13026_ (.A1(_04108_),
    .A2(_04160_),
    .B1(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__nor2b_1 _13027_ (.A(_04023_),
    .B_N(net70),
    .Y(_04165_));
 sky130_fd_sc_hd__clkbuf_8 _13028_ (.A(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__a21oi_1 _13029_ (.A1(_04030_),
    .A2(_04164_),
    .B1(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__buf_4 _13030_ (.A(_03893_),
    .X(_04168_));
 sky130_fd_sc_hd__nand2_1 _13031_ (.A(\samples_imag[0][6] ),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__o21ai_1 _13032_ (.A1(_04043_),
    .A2(_04167_),
    .B1(_04169_),
    .Y(_00304_));
 sky130_fd_sc_hd__buf_4 _13033_ (.A(_03142_),
    .X(_04170_));
 sky130_fd_sc_hd__buf_4 _13034_ (.A(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__or2_1 _13035_ (.A(_03983_),
    .B(_03992_),
    .X(_04172_));
 sky130_fd_sc_hd__buf_6 _13036_ (.A(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__nor2_2 _13037_ (.A(_04044_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__a21oi_1 _13038_ (.A1(\samples_imag[0][7] ),
    .A2(_04060_),
    .B1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__xnor2_2 _13039_ (.A(_03902_),
    .B(net541),
    .Y(_04176_));
 sky130_fd_sc_hd__nor2_8 _13040_ (.A(net518),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__nor2_2 _13041_ (.A(_03894_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a21oi_1 _13042_ (.A1(_04108_),
    .A2(_04175_),
    .B1(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nor2b_1 _13043_ (.A(_04055_),
    .B_N(net71),
    .Y(_04180_));
 sky130_fd_sc_hd__buf_4 _13044_ (.A(_04180_),
    .X(_04181_));
 sky130_fd_sc_hd__a21oi_1 _13045_ (.A1(_04171_),
    .A2(_04179_),
    .B1(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(\samples_imag[0][7] ),
    .B(_04168_),
    .Y(_04183_));
 sky130_fd_sc_hd__o21ai_1 _13047_ (.A1(_04043_),
    .A2(_04182_),
    .B1(_04183_),
    .Y(_00305_));
 sky130_fd_sc_hd__buf_4 _13048_ (.A(_03892_),
    .X(_04184_));
 sky130_fd_sc_hd__or2_1 _13049_ (.A(_03982_),
    .B(_03992_),
    .X(_04185_));
 sky130_fd_sc_hd__buf_6 _13050_ (.A(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__nor2_1 _13051_ (.A(_04089_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__a21oi_1 _13052_ (.A1(\samples_imag[0][8] ),
    .A2(_04060_),
    .B1(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__xnor2_2 _13053_ (.A(_03901_),
    .B(net639),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_8 _13054_ (.A(net518),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__nor2_1 _13055_ (.A(_03894_),
    .B(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21oi_1 _13056_ (.A1(_04108_),
    .A2(_04188_),
    .B1(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2b_1 _13057_ (.A(_04055_),
    .B_N(net72),
    .Y(_04193_));
 sky130_fd_sc_hd__buf_6 _13058_ (.A(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__a21oi_1 _13059_ (.A1(_04171_),
    .A2(_04192_),
    .B1(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _13060_ (.A(\samples_imag[0][8] ),
    .B(_04168_),
    .Y(_04196_));
 sky130_fd_sc_hd__o21ai_1 _13061_ (.A1(_04184_),
    .A2(_04195_),
    .B1(_04196_),
    .Y(_00306_));
 sky130_fd_sc_hd__or2_1 _13062_ (.A(_03986_),
    .B(_03992_),
    .X(_04197_));
 sky130_fd_sc_hd__buf_6 _13063_ (.A(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__nor2_1 _13064_ (.A(_04089_),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__a21oi_1 _13065_ (.A1(\samples_imag[0][9] ),
    .A2(_03715_),
    .B1(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__xnor2_2 _13066_ (.A(_03900_),
    .B(_03915_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_8 _13067_ (.A(net518),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__nor2_1 _13068_ (.A(_03894_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21oi_1 _13069_ (.A1(_04108_),
    .A2(_04200_),
    .B1(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__nor2b_1 _13070_ (.A(_04023_),
    .B_N(net73),
    .Y(_04205_));
 sky130_fd_sc_hd__buf_6 _13071_ (.A(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__a21oi_1 _13072_ (.A1(_04171_),
    .A2(_04204_),
    .B1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand2_1 _13073_ (.A(\samples_imag[0][9] ),
    .B(_04168_),
    .Y(_04208_));
 sky130_fd_sc_hd__o21ai_0 _13074_ (.A1(_04184_),
    .A2(_04207_),
    .B1(_04208_),
    .Y(_00307_));
 sky130_fd_sc_hd__nor3b_1 _13075_ (.A(_03837_),
    .B(_03839_),
    .C_N(_03835_),
    .Y(_04209_));
 sky130_fd_sc_hd__a21boi_4 _13076_ (.A1(_03137_),
    .A2(_03887_),
    .B1_N(_03891_),
    .Y(_04210_));
 sky130_fd_sc_hd__o21ai_4 _13077_ (.A1(_03888_),
    .A2(_04209_),
    .B1(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__buf_4 _13078_ (.A(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__buf_4 _13079_ (.A(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_4 _13080_ (.A(_03469_),
    .X(_04214_));
 sky130_fd_sc_hd__or3_1 _13081_ (.A(_03146_),
    .B(net516),
    .C(_03151_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_4 _13082_ (.A(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__buf_4 _13083_ (.A(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__buf_4 _13084_ (.A(_04216_),
    .X(_04218_));
 sky130_fd_sc_hd__nor2_1 _13085_ (.A(_04218_),
    .B(_04211_),
    .Y(_04219_));
 sky130_fd_sc_hd__a22oi_1 _13086_ (.A1(\samples_imag[1][0] ),
    .A2(_04217_),
    .B1(_03994_),
    .B2(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _13087_ (.A(_04214_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_4 _13088_ (.A(net44),
    .B(_03276_),
    .Y(_04222_));
 sky130_fd_sc_hd__nor3_2 _13089_ (.A(_04222_),
    .B(_04212_),
    .C(_03925_),
    .Y(_04223_));
 sky130_fd_sc_hd__o21ai_1 _13090_ (.A1(_04223_),
    .A2(_04221_),
    .B1(_04004_),
    .Y(_04224_));
 sky130_fd_sc_hd__clkbuf_4 _13091_ (.A(_04212_),
    .X(_04225_));
 sky130_fd_sc_hd__nand2_1 _13092_ (.A(\samples_imag[1][0] ),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__o211ai_2 _13093_ (.A1(_04001_),
    .A2(_04213_),
    .B1(_04226_),
    .C1(_04224_),
    .Y(_00308_));
 sky130_fd_sc_hd__buf_4 _13094_ (.A(_04211_),
    .X(_04227_));
 sky130_fd_sc_hd__buf_4 _13095_ (.A(_03469_),
    .X(_04228_));
 sky130_fd_sc_hd__nor2_1 _13096_ (.A(_04006_),
    .B(_04218_),
    .Y(_04229_));
 sky130_fd_sc_hd__a21oi_1 _13097_ (.A1(\samples_imag[1][10] ),
    .A2(_04217_),
    .B1(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__clkbuf_4 _13098_ (.A(_03279_),
    .X(_04231_));
 sky130_fd_sc_hd__nand2_1 _13099_ (.A(_04231_),
    .B(_04020_),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ai_1 _13100_ (.A1(_04228_),
    .A2(_04230_),
    .B1(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__a21oi_1 _13101_ (.A1(_04171_),
    .A2(_04233_),
    .B1(_04025_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _13102_ (.A(\samples_imag[1][10] ),
    .B(_04213_),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ai_1 _13103_ (.A1(_04227_),
    .A2(_04234_),
    .B1(_04235_),
    .Y(_00309_));
 sky130_fd_sc_hd__buf_4 _13104_ (.A(_03142_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_8 _13105_ (.A(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_4 _13106_ (.A(_03279_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_4 _13107_ (.A(_04216_),
    .X(_04239_));
 sky130_fd_sc_hd__buf_4 _13108_ (.A(_04216_),
    .X(_04240_));
 sky130_fd_sc_hd__nor2_1 _13109_ (.A(_04031_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__a21oi_1 _13110_ (.A1(\samples_imag[1][11] ),
    .A2(_04239_),
    .B1(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__clkbuf_4 _13111_ (.A(_03279_),
    .X(_04243_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_04243_),
    .B(_04036_),
    .Y(_04244_));
 sky130_fd_sc_hd__o21ai_1 _13113_ (.A1(_04238_),
    .A2(_04242_),
    .B1(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__buf_4 _13114_ (.A(_04212_),
    .X(_04246_));
 sky130_fd_sc_hd__a211oi_1 _13115_ (.A1(_04245_),
    .A2(_04237_),
    .B1(_04246_),
    .C1(_04040_),
    .Y(_04247_));
 sky130_fd_sc_hd__a21oi_1 _13116_ (.A1(_03305_),
    .A2(_04213_),
    .B1(_04247_),
    .Y(_00310_));
 sky130_fd_sc_hd__nor2_1 _13117_ (.A(_04045_),
    .B(_04218_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21oi_1 _13118_ (.A1(\samples_imag[1][12] ),
    .A2(_04217_),
    .B1(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _13119_ (.A(_04231_),
    .B(_04052_),
    .Y(_04250_));
 sky130_fd_sc_hd__o21ai_1 _13120_ (.A1(_04228_),
    .A2(_04249_),
    .B1(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21oi_1 _13121_ (.A1(_04171_),
    .A2(_04251_),
    .B1(_04057_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _13122_ (.A(\samples_imag[1][12] ),
    .B(_04213_),
    .Y(_04253_));
 sky130_fd_sc_hd__o21ai_1 _13123_ (.A1(_04227_),
    .A2(_04252_),
    .B1(_04253_),
    .Y(_00311_));
 sky130_fd_sc_hd__nor2_1 _13124_ (.A(_04061_),
    .B(_04240_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21oi_1 _13125_ (.A1(\samples_imag[1][13] ),
    .A2(_04239_),
    .B1(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_1 _13126_ (.A(_04243_),
    .B(_04066_),
    .Y(_04256_));
 sky130_fd_sc_hd__o21ai_1 _13127_ (.A1(_04238_),
    .A2(_04255_),
    .B1(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__a211oi_1 _13128_ (.A1(_04257_),
    .A2(_04237_),
    .B1(_04246_),
    .C1(_04070_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21oi_1 _13129_ (.A1(_03761_),
    .A2(_04213_),
    .B1(_04258_),
    .Y(_00312_));
 sky130_fd_sc_hd__nor2_1 _13130_ (.A(_04218_),
    .B(_04073_),
    .Y(_04259_));
 sky130_fd_sc_hd__a21oi_1 _13131_ (.A1(\samples_imag[1][14] ),
    .A2(_04217_),
    .B1(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__nand2_1 _13132_ (.A(_04231_),
    .B(_04080_),
    .Y(_04261_));
 sky130_fd_sc_hd__o21ai_1 _13133_ (.A1(_04228_),
    .A2(_04260_),
    .B1(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21oi_1 _13134_ (.A1(_04171_),
    .A2(_04262_),
    .B1(_04084_),
    .Y(_04263_));
 sky130_fd_sc_hd__nand2_1 _13135_ (.A(\samples_imag[1][14] ),
    .B(_04213_),
    .Y(_04264_));
 sky130_fd_sc_hd__o21ai_1 _13136_ (.A1(_04227_),
    .A2(_04263_),
    .B1(_04264_),
    .Y(_00313_));
 sky130_fd_sc_hd__clkbuf_4 _13137_ (.A(_04216_),
    .X(_04265_));
 sky130_fd_sc_hd__nand2_1 _13138_ (.A(\samples_imag[1][15] ),
    .B(_04216_),
    .Y(_04266_));
 sky130_fd_sc_hd__o211ai_1 _13139_ (.A1(_04265_),
    .A2(_04090_),
    .B1(_04266_),
    .C1(_04222_),
    .Y(_04267_));
 sky130_fd_sc_hd__o21ai_0 _13140_ (.A1(_04222_),
    .A2(net524),
    .B1(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__a211oi_1 _13141_ (.A1(_04088_),
    .A2(_04268_),
    .B1(_04212_),
    .C1(_04095_),
    .Y(_04269_));
 sky130_fd_sc_hd__a21o_1 _13142_ (.A1(\samples_imag[1][15] ),
    .A2(_04246_),
    .B1(_04269_),
    .X(_00314_));
 sky130_fd_sc_hd__nor2_1 _13143_ (.A(_04240_),
    .B(net647),
    .Y(_04270_));
 sky130_fd_sc_hd__a21oi_1 _13144_ (.A1(\samples_imag[1][1] ),
    .A2(_04239_),
    .B1(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_1 _13145_ (.A(_04101_),
    .B(_04243_),
    .Y(_04272_));
 sky130_fd_sc_hd__o21ai_1 _13146_ (.A1(_04238_),
    .A2(_04271_),
    .B1(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a211oi_1 _13147_ (.A1(_04273_),
    .A2(_04237_),
    .B1(_04246_),
    .C1(_04105_),
    .Y(_04274_));
 sky130_fd_sc_hd__a21oi_1 _13148_ (.A1(_03214_),
    .A2(_04213_),
    .B1(_04274_),
    .Y(_00315_));
 sky130_fd_sc_hd__nor2_1 _13149_ (.A(_04109_),
    .B(_04218_),
    .Y(_04275_));
 sky130_fd_sc_hd__a21oi_1 _13150_ (.A1(\samples_imag[1][2] ),
    .A2(_04217_),
    .B1(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(_04231_),
    .B(_04114_),
    .Y(_04277_));
 sky130_fd_sc_hd__o21ai_1 _13152_ (.A1(_04228_),
    .A2(_04276_),
    .B1(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__a21oi_1 _13153_ (.A1(_04171_),
    .A2(_04278_),
    .B1(_04118_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _13154_ (.A(\samples_imag[1][2] ),
    .B(_04213_),
    .Y(_04280_));
 sky130_fd_sc_hd__o21ai_1 _13155_ (.A1(_04279_),
    .A2(_04227_),
    .B1(_04280_),
    .Y(_00316_));
 sky130_fd_sc_hd__nor2_1 _13156_ (.A(_04218_),
    .B(_04121_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21oi_1 _13157_ (.A1(\samples_imag[1][3] ),
    .A2(_04217_),
    .B1(_04281_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_1 _13158_ (.A(_04238_),
    .B(_04126_),
    .Y(_04283_));
 sky130_fd_sc_hd__o21ai_1 _13159_ (.A1(_04228_),
    .A2(_04282_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__a21oi_1 _13160_ (.A1(_04284_),
    .A2(_04171_),
    .B1(_04130_),
    .Y(_04285_));
 sky130_fd_sc_hd__buf_4 _13161_ (.A(_04212_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_1 _13162_ (.A(\samples_imag[1][3] ),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__o21ai_1 _13163_ (.A1(_04227_),
    .A2(_04285_),
    .B1(_04287_),
    .Y(_00317_));
 sky130_fd_sc_hd__nor2_1 _13164_ (.A(_04133_),
    .B(_04218_),
    .Y(_04288_));
 sky130_fd_sc_hd__a21oi_1 _13165_ (.A1(\samples_imag[1][4] ),
    .A2(_04217_),
    .B1(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _13166_ (.A(_04238_),
    .B(_04138_),
    .Y(_04290_));
 sky130_fd_sc_hd__o21ai_1 _13167_ (.A1(_04231_),
    .A2(_04289_),
    .B1(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a21oi_1 _13168_ (.A1(_04171_),
    .A2(_04291_),
    .B1(_04142_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand2_1 _13169_ (.A(\samples_imag[1][4] ),
    .B(_04286_),
    .Y(_04293_));
 sky130_fd_sc_hd__o21ai_1 _13170_ (.A1(_04227_),
    .A2(_04292_),
    .B1(_04293_),
    .Y(_00318_));
 sky130_fd_sc_hd__nor2_1 _13171_ (.A(_04145_),
    .B(_04218_),
    .Y(_04294_));
 sky130_fd_sc_hd__a21oi_1 _13172_ (.A1(\samples_imag[1][5] ),
    .A2(_04239_),
    .B1(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _13173_ (.A(_04238_),
    .B(_04150_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_1 _13174_ (.A1(_04231_),
    .A2(_04295_),
    .B1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a21oi_1 _13175_ (.A1(_04171_),
    .A2(_04297_),
    .B1(_04154_),
    .Y(_04298_));
 sky130_fd_sc_hd__nand2_1 _13176_ (.A(\samples_imag[1][5] ),
    .B(_04286_),
    .Y(_04299_));
 sky130_fd_sc_hd__o21ai_1 _13177_ (.A1(_04227_),
    .A2(_04298_),
    .B1(_04299_),
    .Y(_00319_));
 sky130_fd_sc_hd__clkbuf_4 _13178_ (.A(_04170_),
    .X(_04300_));
 sky130_fd_sc_hd__nor2_2 _13179_ (.A(_04218_),
    .B(_04158_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _13180_ (.A1(\samples_imag[1][6] ),
    .A2(_04239_),
    .B1(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _13181_ (.A(_04238_),
    .B(_04162_),
    .Y(_04303_));
 sky130_fd_sc_hd__o21ai_1 _13182_ (.A1(_04231_),
    .A2(_04302_),
    .B1(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__a21oi_1 _13183_ (.A1(_04300_),
    .A2(_04304_),
    .B1(_04166_),
    .Y(_04305_));
 sky130_fd_sc_hd__nand2_1 _13184_ (.A(\samples_imag[1][6] ),
    .B(_04286_),
    .Y(_04306_));
 sky130_fd_sc_hd__o21ai_1 _13185_ (.A1(_04227_),
    .A2(_04305_),
    .B1(_04306_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_1 _13186_ (.A(_04216_),
    .B(_04173_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_1 _13187_ (.A1(\samples_imag[1][7] ),
    .A2(_04239_),
    .B1(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_04243_),
    .B(_04177_),
    .Y(_04309_));
 sky130_fd_sc_hd__o21ai_1 _13189_ (.A1(_04243_),
    .A2(_04308_),
    .B1(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__a211oi_2 _13190_ (.A1(_04237_),
    .A2(_04310_),
    .B1(_04212_),
    .C1(_04181_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21oi_1 _13191_ (.A1(_03359_),
    .A2(_04213_),
    .B1(_04311_),
    .Y(_00321_));
 sky130_fd_sc_hd__nor2_2 _13192_ (.A(_04265_),
    .B(_04186_),
    .Y(_04312_));
 sky130_fd_sc_hd__a21oi_1 _13193_ (.A1(\samples_imag[1][8] ),
    .A2(_04239_),
    .B1(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _13194_ (.A(_04238_),
    .B(_04190_),
    .Y(_04314_));
 sky130_fd_sc_hd__o21ai_1 _13195_ (.A1(_04231_),
    .A2(_04313_),
    .B1(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__a21oi_1 _13196_ (.A1(_04300_),
    .A2(_04315_),
    .B1(_04194_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(\samples_imag[1][8] ),
    .B(_04286_),
    .Y(_04317_));
 sky130_fd_sc_hd__o21ai_1 _13198_ (.A1(_04227_),
    .A2(_04316_),
    .B1(_04317_),
    .Y(_00322_));
 sky130_fd_sc_hd__buf_4 _13199_ (.A(_04211_),
    .X(_04318_));
 sky130_fd_sc_hd__nor2_1 _13200_ (.A(_04265_),
    .B(_04198_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _13201_ (.A1(\samples_imag[1][9] ),
    .A2(_04239_),
    .B1(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_1 _13202_ (.A(_04238_),
    .B(_04202_),
    .Y(_04321_));
 sky130_fd_sc_hd__o21ai_1 _13203_ (.A1(_04231_),
    .A2(_04320_),
    .B1(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21oi_1 _13204_ (.A1(_04300_),
    .A2(_04322_),
    .B1(_04206_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(\samples_imag[1][9] ),
    .B(_04286_),
    .Y(_04324_));
 sky130_fd_sc_hd__o21ai_1 _13206_ (.A1(_04318_),
    .A2(_04323_),
    .B1(_04324_),
    .Y(_00323_));
 sky130_fd_sc_hd__nor3b_1 _13207_ (.A(_03835_),
    .B(_03839_),
    .C_N(_03837_),
    .Y(_04325_));
 sky130_fd_sc_hd__o21ai_4 _13208_ (.A1(_03888_),
    .A2(_04325_),
    .B1(_04210_),
    .Y(_04326_));
 sky130_fd_sc_hd__clkbuf_4 _13209_ (.A(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__buf_4 _13210_ (.A(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_4 _13211_ (.A(_03437_),
    .X(_04329_));
 sky130_fd_sc_hd__nand2b_1 _13212_ (.A_N(net539),
    .B(_03151_),
    .Y(_04330_));
 sky130_fd_sc_hd__clkbuf_4 _13213_ (.A(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_4 _13214_ (.A(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__buf_4 _13215_ (.A(_04331_),
    .X(_04333_));
 sky130_fd_sc_hd__nor2_1 _13216_ (.A(_04333_),
    .B(_04326_),
    .Y(_04334_));
 sky130_fd_sc_hd__a22oi_1 _13217_ (.A1(\samples_imag[2][0] ),
    .A2(_04332_),
    .B1(_03994_),
    .B2(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__nor2_1 _13218_ (.A(_04329_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_4 _13219_ (.A(_03296_),
    .B(_03292_),
    .Y(_04337_));
 sky130_fd_sc_hd__nor3_2 _13220_ (.A(_04337_),
    .B(_04327_),
    .C(_03925_),
    .Y(_04338_));
 sky130_fd_sc_hd__o21ai_1 _13221_ (.A1(_04336_),
    .A2(_04338_),
    .B1(_04004_),
    .Y(_04339_));
 sky130_fd_sc_hd__clkbuf_4 _13222_ (.A(_04327_),
    .X(_04340_));
 sky130_fd_sc_hd__nand2_1 _13223_ (.A(\samples_imag[2][0] ),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__o211ai_1 _13224_ (.A1(_04001_),
    .A2(_04328_),
    .B1(_04341_),
    .C1(_04339_),
    .Y(_00324_));
 sky130_fd_sc_hd__clkbuf_4 _13225_ (.A(_04326_),
    .X(_04342_));
 sky130_fd_sc_hd__buf_4 _13226_ (.A(_03437_),
    .X(_04343_));
 sky130_fd_sc_hd__nor2_1 _13227_ (.A(_04333_),
    .B(_04006_),
    .Y(_04344_));
 sky130_fd_sc_hd__a21oi_1 _13228_ (.A1(\samples_imag[2][10] ),
    .A2(_04332_),
    .B1(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__clkbuf_4 _13229_ (.A(_03275_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _13230_ (.A(_04346_),
    .B(_04020_),
    .Y(_04347_));
 sky130_fd_sc_hd__o21ai_1 _13231_ (.A1(_04343_),
    .A2(_04345_),
    .B1(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(_04300_),
    .A2(_04348_),
    .B1(_04025_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _13233_ (.A(\samples_imag[2][10] ),
    .B(_04328_),
    .Y(_04350_));
 sky130_fd_sc_hd__o21ai_1 _13234_ (.A1(_04342_),
    .A2(_04349_),
    .B1(_04350_),
    .Y(_00325_));
 sky130_fd_sc_hd__nor2_1 _13235_ (.A(_04031_),
    .B(_04333_),
    .Y(_04351_));
 sky130_fd_sc_hd__a21oi_1 _13236_ (.A1(\samples_imag[2][11] ),
    .A2(_04332_),
    .B1(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__clkbuf_4 _13237_ (.A(_03437_),
    .X(_04353_));
 sky130_fd_sc_hd__nand2_1 _13238_ (.A(_04353_),
    .B(_04036_),
    .Y(_04354_));
 sky130_fd_sc_hd__o21ai_1 _13239_ (.A1(_04343_),
    .A2(_04352_),
    .B1(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__a21oi_1 _13240_ (.A1(_04300_),
    .A2(_04355_),
    .B1(_04040_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2_1 _13241_ (.A(\samples_imag[2][11] ),
    .B(_04328_),
    .Y(_04357_));
 sky130_fd_sc_hd__o21ai_1 _13242_ (.A1(_04342_),
    .A2(_04356_),
    .B1(_04357_),
    .Y(_00326_));
 sky130_fd_sc_hd__clkbuf_4 _13243_ (.A(_04331_),
    .X(_04358_));
 sky130_fd_sc_hd__nor2_2 _13244_ (.A(_04333_),
    .B(_04045_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21oi_1 _13245_ (.A1(\samples_imag[2][12] ),
    .A2(_04358_),
    .B1(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_1 _13246_ (.A(_04353_),
    .B(_04052_),
    .Y(_04361_));
 sky130_fd_sc_hd__o21ai_1 _13247_ (.A1(_04343_),
    .A2(_04360_),
    .B1(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__a21oi_1 _13248_ (.A1(_04300_),
    .A2(_04362_),
    .B1(_04057_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _13249_ (.A(\samples_imag[2][12] ),
    .B(_04328_),
    .Y(_04364_));
 sky130_fd_sc_hd__o21ai_1 _13250_ (.A1(_04342_),
    .A2(_04363_),
    .B1(_04364_),
    .Y(_00327_));
 sky130_fd_sc_hd__nor2_1 _13251_ (.A(_04061_),
    .B(_04333_),
    .Y(_04365_));
 sky130_fd_sc_hd__a21oi_1 _13252_ (.A1(\samples_imag[2][13] ),
    .A2(_04358_),
    .B1(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _13253_ (.A(_04353_),
    .B(_04066_),
    .Y(_04367_));
 sky130_fd_sc_hd__o21ai_1 _13254_ (.A1(_04343_),
    .A2(_04366_),
    .B1(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__a21oi_1 _13255_ (.A1(_04300_),
    .A2(_04368_),
    .B1(_04070_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _13256_ (.A(\samples_imag[2][13] ),
    .B(_04328_),
    .Y(_04370_));
 sky130_fd_sc_hd__o21ai_1 _13257_ (.A1(_04342_),
    .A2(_04369_),
    .B1(_04370_),
    .Y(_00328_));
 sky130_fd_sc_hd__nor2_1 _13258_ (.A(_04333_),
    .B(_04073_),
    .Y(_04371_));
 sky130_fd_sc_hd__a21oi_1 _13259_ (.A1(\samples_imag[2][14] ),
    .A2(_04358_),
    .B1(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _13260_ (.A(_04353_),
    .B(_04080_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21ai_1 _13261_ (.A1(_04343_),
    .A2(_04372_),
    .B1(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__a21oi_1 _13262_ (.A1(_04300_),
    .A2(_04374_),
    .B1(_04084_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand2_1 _13263_ (.A(\samples_imag[2][14] ),
    .B(_04328_),
    .Y(_04376_));
 sky130_fd_sc_hd__o21ai_1 _13264_ (.A1(_04375_),
    .A2(_04342_),
    .B1(_04376_),
    .Y(_00329_));
 sky130_fd_sc_hd__buf_4 _13265_ (.A(_04327_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_4 _13266_ (.A(_04331_),
    .X(_04378_));
 sky130_fd_sc_hd__nand2_1 _13267_ (.A(\samples_imag[2][15] ),
    .B(_04331_),
    .Y(_04379_));
 sky130_fd_sc_hd__o211ai_1 _13268_ (.A1(_04378_),
    .A2(_04090_),
    .B1(_04379_),
    .C1(_04337_),
    .Y(_04380_));
 sky130_fd_sc_hd__o21ai_1 _13269_ (.A1(_04337_),
    .A2(net54),
    .B1(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__a211oi_2 _13270_ (.A1(_04088_),
    .A2(_04381_),
    .B1(_04327_),
    .C1(_04095_),
    .Y(_04382_));
 sky130_fd_sc_hd__a21o_1 _13271_ (.A1(\samples_imag[2][15] ),
    .A2(_04377_),
    .B1(_04382_),
    .X(_00330_));
 sky130_fd_sc_hd__nor2_2 _13272_ (.A(_04333_),
    .B(_04097_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21oi_1 _13273_ (.A1(\samples_imag[2][1] ),
    .A2(_04358_),
    .B1(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__nand2_1 _13274_ (.A(_04353_),
    .B(_04101_),
    .Y(_04385_));
 sky130_fd_sc_hd__o21ai_1 _13275_ (.A1(_04346_),
    .A2(_04384_),
    .B1(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__a21oi_1 _13276_ (.A1(_04300_),
    .A2(_04386_),
    .B1(_04105_),
    .Y(_04387_));
 sky130_fd_sc_hd__buf_4 _13277_ (.A(_04327_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _13278_ (.A(\samples_imag[2][1] ),
    .B(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__o21ai_1 _13279_ (.A1(_04387_),
    .A2(_04342_),
    .B1(_04389_),
    .Y(_00331_));
 sky130_fd_sc_hd__nor2_1 _13280_ (.A(_04109_),
    .B(_04378_),
    .Y(_04390_));
 sky130_fd_sc_hd__a21oi_1 _13281_ (.A1(\samples_imag[2][2] ),
    .A2(_04358_),
    .B1(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2_1 _13282_ (.A(_04353_),
    .B(_04114_),
    .Y(_04392_));
 sky130_fd_sc_hd__o21ai_1 _13283_ (.A1(_04346_),
    .A2(_04391_),
    .B1(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a21oi_1 _13284_ (.A1(_04300_),
    .A2(_04393_),
    .B1(_04118_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(\samples_imag[2][2] ),
    .B(_04388_),
    .Y(_04395_));
 sky130_fd_sc_hd__o21ai_1 _13286_ (.A1(_04342_),
    .A2(_04394_),
    .B1(_04395_),
    .Y(_00332_));
 sky130_fd_sc_hd__buf_2 _13287_ (.A(_04170_),
    .X(_04396_));
 sky130_fd_sc_hd__nor2_2 _13288_ (.A(_04378_),
    .B(_04121_),
    .Y(_04397_));
 sky130_fd_sc_hd__a21oi_1 _13289_ (.A1(\samples_imag[2][3] ),
    .A2(_04358_),
    .B1(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _13290_ (.A(_04353_),
    .B(_04126_),
    .Y(_04399_));
 sky130_fd_sc_hd__o21ai_1 _13291_ (.A1(_04346_),
    .A2(_04398_),
    .B1(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__a21oi_1 _13292_ (.A1(_04396_),
    .A2(_04400_),
    .B1(_04130_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _13293_ (.A(\samples_imag[2][3] ),
    .B(_04388_),
    .Y(_04402_));
 sky130_fd_sc_hd__o21ai_1 _13294_ (.A1(_04342_),
    .A2(_04401_),
    .B1(_04402_),
    .Y(_00333_));
 sky130_fd_sc_hd__nor2_1 _13295_ (.A(_04133_),
    .B(_04378_),
    .Y(_04403_));
 sky130_fd_sc_hd__a21oi_1 _13296_ (.A1(\samples_imag[2][4] ),
    .A2(_04358_),
    .B1(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(_04353_),
    .B(_04138_),
    .Y(_04405_));
 sky130_fd_sc_hd__o21ai_1 _13298_ (.A1(_04346_),
    .A2(_04404_),
    .B1(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__a21oi_1 _13299_ (.A1(_04396_),
    .A2(_04406_),
    .B1(_04142_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_1 _13300_ (.A(\samples_imag[2][4] ),
    .B(_04388_),
    .Y(_04408_));
 sky130_fd_sc_hd__o21ai_1 _13301_ (.A1(_04342_),
    .A2(_04407_),
    .B1(_04408_),
    .Y(_00334_));
 sky130_fd_sc_hd__buf_4 _13302_ (.A(_04326_),
    .X(_04409_));
 sky130_fd_sc_hd__nor2_2 _13303_ (.A(_04378_),
    .B(_04145_),
    .Y(_04410_));
 sky130_fd_sc_hd__a21oi_1 _13304_ (.A1(\samples_imag[2][5] ),
    .A2(_04358_),
    .B1(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand2_1 _13305_ (.A(_04353_),
    .B(_04150_),
    .Y(_04412_));
 sky130_fd_sc_hd__o21ai_1 _13306_ (.A1(_04346_),
    .A2(_04411_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a21oi_1 _13307_ (.A1(_04396_),
    .A2(_04413_),
    .B1(_04154_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand2_1 _13308_ (.A(\samples_imag[2][5] ),
    .B(_04388_),
    .Y(_04415_));
 sky130_fd_sc_hd__o21ai_1 _13309_ (.A1(_04409_),
    .A2(_04414_),
    .B1(_04415_),
    .Y(_00335_));
 sky130_fd_sc_hd__nor2_1 _13310_ (.A(_04378_),
    .B(_04158_),
    .Y(_04416_));
 sky130_fd_sc_hd__a21oi_1 _13311_ (.A1(\samples_imag[2][6] ),
    .A2(_04358_),
    .B1(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(_04353_),
    .B(_04162_),
    .Y(_04418_));
 sky130_fd_sc_hd__o21ai_1 _13313_ (.A1(_04346_),
    .A2(_04417_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a21oi_1 _13314_ (.A1(_04396_),
    .A2(_04419_),
    .B1(_04166_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand2_1 _13315_ (.A(\samples_imag[2][6] ),
    .B(_04388_),
    .Y(_04421_));
 sky130_fd_sc_hd__o21ai_1 _13316_ (.A1(_04409_),
    .A2(_04420_),
    .B1(_04421_),
    .Y(_00336_));
 sky130_fd_sc_hd__nor2_1 _13317_ (.A(_04378_),
    .B(_04173_),
    .Y(_04422_));
 sky130_fd_sc_hd__a21oi_1 _13318_ (.A1(\samples_imag[2][7] ),
    .A2(_04358_),
    .B1(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__clkbuf_4 _13319_ (.A(_03275_),
    .X(_04424_));
 sky130_fd_sc_hd__nand2_1 _13320_ (.A(_04424_),
    .B(_04177_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_1 _13321_ (.A1(_04346_),
    .A2(_04423_),
    .B1(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a21oi_1 _13322_ (.A1(_04396_),
    .A2(_04426_),
    .B1(_04181_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _13323_ (.A(\samples_imag[2][7] ),
    .B(_04388_),
    .Y(_04428_));
 sky130_fd_sc_hd__o21ai_1 _13324_ (.A1(_04409_),
    .A2(_04427_),
    .B1(_04428_),
    .Y(_00337_));
 sky130_fd_sc_hd__buf_4 _13325_ (.A(_04331_),
    .X(_04429_));
 sky130_fd_sc_hd__nor2_1 _13326_ (.A(_04331_),
    .B(_04186_),
    .Y(_04430_));
 sky130_fd_sc_hd__a21oi_1 _13327_ (.A1(\samples_imag[2][8] ),
    .A2(_04429_),
    .B1(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_04424_),
    .B(_04190_),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_1 _13329_ (.A1(_04424_),
    .A2(_04431_),
    .B1(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__a211oi_2 _13330_ (.A1(_04237_),
    .A2(_04433_),
    .B1(_04377_),
    .C1(_04194_),
    .Y(_04434_));
 sky130_fd_sc_hd__a21oi_1 _13331_ (.A1(_03347_),
    .A2(_04328_),
    .B1(_04434_),
    .Y(_00338_));
 sky130_fd_sc_hd__nor2_1 _13332_ (.A(_04378_),
    .B(_04198_),
    .Y(_04435_));
 sky130_fd_sc_hd__a21oi_1 _13333_ (.A1(\samples_imag[2][9] ),
    .A2(_04429_),
    .B1(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand2_1 _13334_ (.A(_04424_),
    .B(_04202_),
    .Y(_04437_));
 sky130_fd_sc_hd__o21ai_1 _13335_ (.A1(_04346_),
    .A2(_04436_),
    .B1(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__a21oi_1 _13336_ (.A1(_04396_),
    .A2(_04438_),
    .B1(_04206_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _13337_ (.A(\samples_imag[2][9] ),
    .B(_04388_),
    .Y(_04440_));
 sky130_fd_sc_hd__o21ai_1 _13338_ (.A1(_04409_),
    .A2(_04439_),
    .B1(_04440_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _13339_ (.A(_03837_),
    .B(_03835_),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_1 _13340_ (.A(_03839_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__o21ai_4 _13341_ (.A1(_03888_),
    .A2(_04442_),
    .B1(_04210_),
    .Y(_04443_));
 sky130_fd_sc_hd__buf_4 _13342_ (.A(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__or2_0 _13343_ (.A(_03158_),
    .B(net539),
    .X(_04445_));
 sky130_fd_sc_hd__buf_4 _13344_ (.A(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__buf_4 _13345_ (.A(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__nor2_1 _13346_ (.A(_04446_),
    .B(_04444_),
    .Y(_04448_));
 sky130_fd_sc_hd__a22oi_1 _13347_ (.A1(\samples_imag[3][0] ),
    .A2(_04447_),
    .B1(_03994_),
    .B2(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__nand2_4 _13348_ (.A(_03296_),
    .B(_03287_),
    .Y(_04450_));
 sky130_fd_sc_hd__or2_1 _13349_ (.A(_04450_),
    .B(_04444_),
    .X(_04451_));
 sky130_fd_sc_hd__o22ai_2 _13350_ (.A1(_03439_),
    .A2(_04449_),
    .B1(_04451_),
    .B2(_03925_),
    .Y(_04452_));
 sky130_fd_sc_hd__nor2_1 _13351_ (.A(_04001_),
    .B(_04444_),
    .Y(_04453_));
 sky130_fd_sc_hd__a221o_1 _13352_ (.A1(\samples_imag[3][0] ),
    .A2(_04444_),
    .B1(_04452_),
    .B2(_03999_),
    .C1(_04453_),
    .X(_00340_));
 sky130_fd_sc_hd__buf_4 _13353_ (.A(_04444_),
    .X(_04454_));
 sky130_fd_sc_hd__buf_4 _13354_ (.A(_03439_),
    .X(_04455_));
 sky130_fd_sc_hd__buf_4 _13355_ (.A(_04446_),
    .X(_04456_));
 sky130_fd_sc_hd__nor2_2 _13356_ (.A(_04447_),
    .B(_04006_),
    .Y(_04457_));
 sky130_fd_sc_hd__a21oi_1 _13357_ (.A1(\samples_imag[3][10] ),
    .A2(_04456_),
    .B1(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__clkbuf_4 _13358_ (.A(_03439_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _13359_ (.A(_04459_),
    .B(_04020_),
    .Y(_04460_));
 sky130_fd_sc_hd__o21ai_1 _13360_ (.A1(_04455_),
    .A2(_04458_),
    .B1(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__a21oi_1 _13361_ (.A1(_04396_),
    .A2(_04461_),
    .B1(_04025_),
    .Y(_04462_));
 sky130_fd_sc_hd__buf_2 _13362_ (.A(_04444_),
    .X(_04463_));
 sky130_fd_sc_hd__nand2_1 _13363_ (.A(\samples_imag[3][10] ),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__o21ai_1 _13364_ (.A1(_04462_),
    .A2(_04454_),
    .B1(_04464_),
    .Y(_00341_));
 sky130_fd_sc_hd__nor2_2 _13365_ (.A(_04031_),
    .B(_04447_),
    .Y(_04465_));
 sky130_fd_sc_hd__a21oi_1 _13366_ (.A1(\samples_imag[3][11] ),
    .A2(_04456_),
    .B1(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__buf_2 _13367_ (.A(_03439_),
    .X(_04467_));
 sky130_fd_sc_hd__nand2_1 _13368_ (.A(_04467_),
    .B(_04036_),
    .Y(_04468_));
 sky130_fd_sc_hd__o21ai_1 _13369_ (.A1(_04455_),
    .A2(_04466_),
    .B1(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__a21oi_1 _13370_ (.A1(_04396_),
    .A2(_04469_),
    .B1(_04040_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _13371_ (.A(\samples_imag[3][11] ),
    .B(_04463_),
    .Y(_04471_));
 sky130_fd_sc_hd__o21ai_1 _13372_ (.A1(_04470_),
    .A2(_04454_),
    .B1(_04471_),
    .Y(_00342_));
 sky130_fd_sc_hd__clkbuf_2 _13373_ (.A(_04443_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_2 _13374_ (.A(_04447_),
    .B(_04045_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21oi_1 _13375_ (.A1(\samples_imag[3][12] ),
    .A2(_04456_),
    .B1(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__nand2_1 _13376_ (.A(_04052_),
    .B(_04467_),
    .Y(_04475_));
 sky130_fd_sc_hd__o21ai_1 _13377_ (.A1(_04455_),
    .A2(_04474_),
    .B1(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21oi_1 _13378_ (.A1(_04476_),
    .A2(_04396_),
    .B1(_04057_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_1 _13379_ (.A(\samples_imag[3][12] ),
    .B(_04463_),
    .Y(_04478_));
 sky130_fd_sc_hd__o21ai_1 _13380_ (.A1(_04472_),
    .A2(_04477_),
    .B1(_04478_),
    .Y(_00343_));
 sky130_fd_sc_hd__nor2_2 _13381_ (.A(_04061_),
    .B(_04447_),
    .Y(_04479_));
 sky130_fd_sc_hd__a21oi_1 _13382_ (.A1(\samples_imag[3][13] ),
    .A2(_04456_),
    .B1(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2_1 _13383_ (.A(_04467_),
    .B(_04066_),
    .Y(_04481_));
 sky130_fd_sc_hd__o21ai_1 _13384_ (.A1(_04455_),
    .A2(_04480_),
    .B1(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__a21oi_1 _13385_ (.A1(_04396_),
    .A2(_04482_),
    .B1(_04070_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _13386_ (.A(\samples_imag[3][13] ),
    .B(_04463_),
    .Y(_04484_));
 sky130_fd_sc_hd__o21ai_1 _13387_ (.A1(_04472_),
    .A2(_04483_),
    .B1(_04484_),
    .Y(_00344_));
 sky130_fd_sc_hd__buf_2 _13388_ (.A(_04170_),
    .X(_04485_));
 sky130_fd_sc_hd__buf_2 _13389_ (.A(_04446_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _13390_ (.A(_04073_),
    .B(_04447_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_1 _13391_ (.A1(\samples_imag[3][14] ),
    .A2(_04486_),
    .B1(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_1 _13392_ (.A(_04467_),
    .B(_04080_),
    .Y(_04489_));
 sky130_fd_sc_hd__o21ai_1 _13393_ (.A1(_04455_),
    .A2(_04488_),
    .B1(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__a21oi_1 _13394_ (.A1(_04485_),
    .A2(_04490_),
    .B1(_04084_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2_1 _13395_ (.A(\samples_imag[3][14] ),
    .B(_04463_),
    .Y(_04492_));
 sky130_fd_sc_hd__o21ai_1 _13396_ (.A1(_04472_),
    .A2(_04491_),
    .B1(_04492_),
    .Y(_00345_));
 sky130_fd_sc_hd__buf_2 _13397_ (.A(_04444_),
    .X(_04493_));
 sky130_fd_sc_hd__buf_4 _13398_ (.A(_04446_),
    .X(_04494_));
 sky130_fd_sc_hd__nand2_1 _13399_ (.A(\samples_imag[3][15] ),
    .B(_04446_),
    .Y(_04495_));
 sky130_fd_sc_hd__o211ai_1 _13400_ (.A1(_04494_),
    .A2(_04090_),
    .B1(_04495_),
    .C1(_04450_),
    .Y(_04496_));
 sky130_fd_sc_hd__o21ai_0 _13401_ (.A1(_04450_),
    .A2(net54),
    .B1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__a211oi_1 _13402_ (.A1(_04088_),
    .A2(_04497_),
    .B1(_04493_),
    .C1(_04095_),
    .Y(_04498_));
 sky130_fd_sc_hd__a21o_1 _13403_ (.A1(\samples_imag[3][15] ),
    .A2(_04493_),
    .B1(_04498_),
    .X(_00346_));
 sky130_fd_sc_hd__nor2_1 _13404_ (.A(_04447_),
    .B(_04097_),
    .Y(_04499_));
 sky130_fd_sc_hd__a21oi_1 _13405_ (.A1(\samples_imag[3][1] ),
    .A2(_04486_),
    .B1(_04499_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(_04467_),
    .B(_04101_),
    .Y(_04501_));
 sky130_fd_sc_hd__o21ai_1 _13407_ (.A1(_04455_),
    .A2(_04500_),
    .B1(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__a21oi_1 _13408_ (.A1(_04485_),
    .A2(_04502_),
    .B1(_04105_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(\samples_imag[3][1] ),
    .B(_04463_),
    .Y(_04504_));
 sky130_fd_sc_hd__o21ai_1 _13410_ (.A1(_04472_),
    .A2(_04503_),
    .B1(_04504_),
    .Y(_00347_));
 sky130_fd_sc_hd__nor2_2 _13411_ (.A(_04447_),
    .B(_04109_),
    .Y(_04505_));
 sky130_fd_sc_hd__a21oi_1 _13412_ (.A1(\samples_imag[3][2] ),
    .A2(_04486_),
    .B1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2_1 _13413_ (.A(_04467_),
    .B(_04114_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21ai_1 _13414_ (.A1(_04459_),
    .A2(_04506_),
    .B1(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21oi_1 _13415_ (.A1(_04485_),
    .A2(_04508_),
    .B1(_04118_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _13416_ (.A(\samples_imag[3][2] ),
    .B(_04463_),
    .Y(_04510_));
 sky130_fd_sc_hd__o21ai_1 _13417_ (.A1(_04472_),
    .A2(_04509_),
    .B1(_04510_),
    .Y(_00348_));
 sky130_fd_sc_hd__nor2_2 _13418_ (.A(_04494_),
    .B(_04121_),
    .Y(_04511_));
 sky130_fd_sc_hd__a21oi_1 _13419_ (.A1(\samples_imag[3][3] ),
    .A2(_04486_),
    .B1(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand2_1 _13420_ (.A(_04467_),
    .B(_04126_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_1 _13421_ (.A1(_04459_),
    .A2(_04512_),
    .B1(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__a21oi_1 _13422_ (.A1(_04485_),
    .A2(_04514_),
    .B1(_04130_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _13423_ (.A(\samples_imag[3][3] ),
    .B(_04463_),
    .Y(_04516_));
 sky130_fd_sc_hd__o21ai_1 _13424_ (.A1(_04472_),
    .A2(_04515_),
    .B1(_04516_),
    .Y(_00349_));
 sky130_fd_sc_hd__nor2_1 _13425_ (.A(_04133_),
    .B(_04494_),
    .Y(_04517_));
 sky130_fd_sc_hd__a21oi_1 _13426_ (.A1(\samples_imag[3][4] ),
    .A2(_04486_),
    .B1(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_1 _13427_ (.A(_04467_),
    .B(_04138_),
    .Y(_04519_));
 sky130_fd_sc_hd__o21ai_1 _13428_ (.A1(_04459_),
    .A2(_04518_),
    .B1(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__a21oi_1 _13429_ (.A1(_04485_),
    .A2(_04520_),
    .B1(_04142_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _13430_ (.A(\samples_imag[3][4] ),
    .B(_04463_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21ai_1 _13431_ (.A1(_04472_),
    .A2(_04521_),
    .B1(_04522_),
    .Y(_00350_));
 sky130_fd_sc_hd__nor2_1 _13432_ (.A(_04145_),
    .B(_04494_),
    .Y(_04523_));
 sky130_fd_sc_hd__a21oi_1 _13433_ (.A1(\samples_imag[3][5] ),
    .A2(_04486_),
    .B1(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand2_1 _13434_ (.A(_04467_),
    .B(_04150_),
    .Y(_04525_));
 sky130_fd_sc_hd__o21ai_1 _13435_ (.A1(_04459_),
    .A2(_04524_),
    .B1(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21oi_1 _13436_ (.A1(_04485_),
    .A2(_04526_),
    .B1(_04154_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_1 _13437_ (.A(\samples_imag[3][5] ),
    .B(_04463_),
    .Y(_04528_));
 sky130_fd_sc_hd__o21ai_1 _13438_ (.A1(_04472_),
    .A2(_04527_),
    .B1(_04528_),
    .Y(_00351_));
 sky130_fd_sc_hd__nor2_1 _13439_ (.A(_04494_),
    .B(_04158_),
    .Y(_04529_));
 sky130_fd_sc_hd__a21oi_1 _13440_ (.A1(\samples_imag[3][6] ),
    .A2(_04486_),
    .B1(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__nand2_1 _13441_ (.A(_04467_),
    .B(_04162_),
    .Y(_04531_));
 sky130_fd_sc_hd__o21ai_1 _13442_ (.A1(_04459_),
    .A2(_04530_),
    .B1(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__a21oi_1 _13443_ (.A1(_04485_),
    .A2(_04532_),
    .B1(_04166_),
    .Y(_04533_));
 sky130_fd_sc_hd__buf_4 _13444_ (.A(_04444_),
    .X(_04534_));
 sky130_fd_sc_hd__nand2_1 _13445_ (.A(\samples_imag[3][6] ),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__o21ai_1 _13446_ (.A1(_04472_),
    .A2(_04533_),
    .B1(_04535_),
    .Y(_00352_));
 sky130_fd_sc_hd__nor2_1 _13447_ (.A(_04494_),
    .B(_04173_),
    .Y(_04536_));
 sky130_fd_sc_hd__a21oi_1 _13448_ (.A1(\samples_imag[3][7] ),
    .A2(_04486_),
    .B1(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _13449_ (.A(_03439_),
    .B(_04177_),
    .Y(_04538_));
 sky130_fd_sc_hd__o21ai_1 _13450_ (.A1(_04459_),
    .A2(_04537_),
    .B1(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__a21oi_1 _13451_ (.A1(_04485_),
    .A2(_04539_),
    .B1(_04181_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _13452_ (.A(\samples_imag[3][7] ),
    .B(_04534_),
    .Y(_04541_));
 sky130_fd_sc_hd__o21ai_1 _13453_ (.A1(_04472_),
    .A2(_04540_),
    .B1(_04541_),
    .Y(_00353_));
 sky130_fd_sc_hd__buf_4 _13454_ (.A(_04443_),
    .X(_04542_));
 sky130_fd_sc_hd__nor2_1 _13455_ (.A(_04494_),
    .B(_04186_),
    .Y(_04543_));
 sky130_fd_sc_hd__a21oi_1 _13456_ (.A1(\samples_imag[3][8] ),
    .A2(_04486_),
    .B1(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _13457_ (.A(_03439_),
    .B(_04190_),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ai_1 _13458_ (.A1(_04459_),
    .A2(_04544_),
    .B1(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__a21oi_1 _13459_ (.A1(_04485_),
    .A2(_04546_),
    .B1(_04194_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(\samples_imag[3][8] ),
    .B(_04534_),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ai_1 _13461_ (.A1(_04542_),
    .A2(_04547_),
    .B1(_04548_),
    .Y(_00354_));
 sky130_fd_sc_hd__nor2_2 _13462_ (.A(_04494_),
    .B(_04198_),
    .Y(_04549_));
 sky130_fd_sc_hd__a21oi_1 _13463_ (.A1(\samples_imag[3][9] ),
    .A2(_04486_),
    .B1(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_2 _13464_ (.A(_03439_),
    .B(_04202_),
    .Y(_04551_));
 sky130_fd_sc_hd__o21ai_1 _13465_ (.A1(_04459_),
    .A2(_04550_),
    .B1(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21oi_1 _13466_ (.A1(_04485_),
    .A2(_04552_),
    .B1(_04206_),
    .Y(_04553_));
 sky130_fd_sc_hd__nand2_1 _13467_ (.A(\samples_imag[3][9] ),
    .B(_04534_),
    .Y(_04554_));
 sky130_fd_sc_hd__o21ai_1 _13468_ (.A1(_04542_),
    .A2(_04553_),
    .B1(_04554_),
    .Y(_00355_));
 sky130_fd_sc_hd__nor3b_1 _13469_ (.A(_03837_),
    .B(_03835_),
    .C_N(_03839_),
    .Y(_04555_));
 sky130_fd_sc_hd__o21ai_4 _13470_ (.A1(_03888_),
    .A2(_04555_),
    .B1(_04210_),
    .Y(_04556_));
 sky130_fd_sc_hd__buf_2 _13471_ (.A(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__buf_2 _13472_ (.A(_03467_),
    .X(_04558_));
 sky130_fd_sc_hd__nand2_2 _13473_ (.A(_03146_),
    .B(_03160_),
    .Y(_04559_));
 sky130_fd_sc_hd__clkbuf_4 _13474_ (.A(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_4 _13475_ (.A(_04559_),
    .X(_04561_));
 sky130_fd_sc_hd__nor2_1 _13476_ (.A(_04561_),
    .B(_04556_),
    .Y(_04562_));
 sky130_fd_sc_hd__a22oi_1 _13477_ (.A1(\samples_imag[4][0] ),
    .A2(_04560_),
    .B1(_03994_),
    .B2(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__clkbuf_4 _13478_ (.A(_03272_),
    .X(_04564_));
 sky130_fd_sc_hd__nor2_1 _13479_ (.A(_04557_),
    .B(_03925_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _13480_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__o21ai_1 _13481_ (.A1(_04558_),
    .A2(_04563_),
    .B1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__nor2_1 _13482_ (.A(_04001_),
    .B(_04557_),
    .Y(_04568_));
 sky130_fd_sc_hd__a221o_1 _13483_ (.A1(\samples_imag[4][0] ),
    .A2(_04557_),
    .B1(_03999_),
    .B2(_04567_),
    .C1(_04568_),
    .X(_00356_));
 sky130_fd_sc_hd__clkbuf_4 _13484_ (.A(_04557_),
    .X(_04569_));
 sky130_fd_sc_hd__buf_2 _13485_ (.A(_04170_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_4 _13486_ (.A(_03467_),
    .X(_04571_));
 sky130_fd_sc_hd__buf_2 _13487_ (.A(_04561_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_4 _13488_ (.A(_04559_),
    .X(_04573_));
 sky130_fd_sc_hd__nor2_2 _13489_ (.A(_04573_),
    .B(_04006_),
    .Y(_04574_));
 sky130_fd_sc_hd__a21oi_1 _13490_ (.A1(\samples_imag[4][10] ),
    .A2(_04572_),
    .B1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__buf_2 _13491_ (.A(_03467_),
    .X(_04576_));
 sky130_fd_sc_hd__nand2_1 _13492_ (.A(_04576_),
    .B(_04020_),
    .Y(_04577_));
 sky130_fd_sc_hd__o21ai_1 _13493_ (.A1(_04575_),
    .A2(_04571_),
    .B1(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__a21oi_1 _13494_ (.A1(_04570_),
    .A2(_04578_),
    .B1(_04025_),
    .Y(_04579_));
 sky130_fd_sc_hd__clkbuf_4 _13495_ (.A(_04557_),
    .X(_04580_));
 sky130_fd_sc_hd__nand2_1 _13496_ (.A(\samples_imag[4][10] ),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o21ai_1 _13497_ (.A1(_04569_),
    .A2(_04579_),
    .B1(_04581_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_2 _13498_ (.A(_04031_),
    .B(_04573_),
    .Y(_04582_));
 sky130_fd_sc_hd__a21oi_1 _13499_ (.A1(\samples_imag[4][11] ),
    .A2(_04572_),
    .B1(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _13500_ (.A(_04576_),
    .B(_04036_),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_1 _13501_ (.A1(_04571_),
    .A2(_04583_),
    .B1(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21oi_1 _13502_ (.A1(_04570_),
    .A2(_04585_),
    .B1(_04040_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand2_1 _13503_ (.A(\samples_imag[4][11] ),
    .B(_04580_),
    .Y(_04587_));
 sky130_fd_sc_hd__o21ai_1 _13504_ (.A1(_04569_),
    .A2(_04586_),
    .B1(_04587_),
    .Y(_00358_));
 sky130_fd_sc_hd__clkbuf_4 _13505_ (.A(_04559_),
    .X(_04588_));
 sky130_fd_sc_hd__nor2_2 _13506_ (.A(_04561_),
    .B(net646),
    .Y(_04589_));
 sky130_fd_sc_hd__a21oi_1 _13507_ (.A1(\samples_imag[4][12] ),
    .A2(_04588_),
    .B1(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _13508_ (.A(_04564_),
    .B(_04052_),
    .Y(_04591_));
 sky130_fd_sc_hd__o21ai_1 _13509_ (.A1(_04564_),
    .A2(_04590_),
    .B1(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__clkbuf_4 _13510_ (.A(_04557_),
    .X(_04593_));
 sky130_fd_sc_hd__a211oi_1 _13511_ (.A1(_04592_),
    .A2(_04237_),
    .B1(_04593_),
    .C1(_04057_),
    .Y(_04594_));
 sky130_fd_sc_hd__a21oi_1 _13512_ (.A1(_03253_),
    .A2(_04580_),
    .B1(_04594_),
    .Y(_00359_));
 sky130_fd_sc_hd__clkbuf_2 _13513_ (.A(_04556_),
    .X(_04595_));
 sky130_fd_sc_hd__nor2_1 _13514_ (.A(_04061_),
    .B(_04573_),
    .Y(_04596_));
 sky130_fd_sc_hd__a21oi_1 _13515_ (.A1(\samples_imag[4][13] ),
    .A2(_04572_),
    .B1(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _13516_ (.A(_04576_),
    .B(_04066_),
    .Y(_04598_));
 sky130_fd_sc_hd__o21ai_1 _13517_ (.A1(_04597_),
    .A2(_04571_),
    .B1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__a21oi_1 _13518_ (.A1(_04599_),
    .A2(_04570_),
    .B1(_04070_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2_1 _13519_ (.A(\samples_imag[4][13] ),
    .B(_04580_),
    .Y(_04601_));
 sky130_fd_sc_hd__o21ai_1 _13520_ (.A1(_04595_),
    .A2(_04600_),
    .B1(_04601_),
    .Y(_00360_));
 sky130_fd_sc_hd__nor2_2 _13521_ (.A(_04573_),
    .B(_04073_),
    .Y(_04602_));
 sky130_fd_sc_hd__a21oi_1 _13522_ (.A1(\samples_imag[4][14] ),
    .A2(_04572_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2_1 _13523_ (.A(_04576_),
    .B(_04080_),
    .Y(_04604_));
 sky130_fd_sc_hd__o21ai_1 _13524_ (.A1(_04571_),
    .A2(_04603_),
    .B1(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__a21oi_1 _13525_ (.A1(_04570_),
    .A2(_04605_),
    .B1(_04084_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_1 _13526_ (.A(\samples_imag[4][14] ),
    .B(_04580_),
    .Y(_04607_));
 sky130_fd_sc_hd__o21ai_1 _13527_ (.A1(_04595_),
    .A2(_04606_),
    .B1(_04607_),
    .Y(_00361_));
 sky130_fd_sc_hd__nor2_1 _13528_ (.A(\samples_imag[4][15] ),
    .B(net549),
    .Y(_04608_));
 sky130_fd_sc_hd__a211oi_1 _13529_ (.A1(net550),
    .A2(_04090_),
    .B1(_04608_),
    .C1(_03467_),
    .Y(_04609_));
 sky130_fd_sc_hd__a21oi_1 _13530_ (.A1(_04564_),
    .A2(net54),
    .B1(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__a211oi_1 _13531_ (.A1(_04088_),
    .A2(_04610_),
    .B1(_04593_),
    .C1(_04095_),
    .Y(_04611_));
 sky130_fd_sc_hd__a21o_1 _13532_ (.A1(\samples_imag[4][15] ),
    .A2(_04593_),
    .B1(_04611_),
    .X(_00362_));
 sky130_fd_sc_hd__nor2_1 _13533_ (.A(_04573_),
    .B(_04097_),
    .Y(_04612_));
 sky130_fd_sc_hd__a21oi_1 _13534_ (.A1(\samples_imag[4][1] ),
    .A2(_04572_),
    .B1(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(_04558_),
    .B(_04101_),
    .Y(_04614_));
 sky130_fd_sc_hd__o21ai_1 _13536_ (.A1(_04613_),
    .A2(_04571_),
    .B1(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__a21oi_1 _13537_ (.A1(_04570_),
    .A2(_04615_),
    .B1(_04105_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _13538_ (.A(\samples_imag[4][1] ),
    .B(_04580_),
    .Y(_04617_));
 sky130_fd_sc_hd__o21ai_1 _13539_ (.A1(_04595_),
    .A2(_04616_),
    .B1(_04617_),
    .Y(_00363_));
 sky130_fd_sc_hd__nor2_2 _13540_ (.A(_04109_),
    .B(_04573_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21oi_1 _13541_ (.A1(\samples_imag[4][2] ),
    .A2(_04572_),
    .B1(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _13542_ (.A(_04558_),
    .B(_04114_),
    .Y(_04620_));
 sky130_fd_sc_hd__o21ai_1 _13543_ (.A1(_04619_),
    .A2(_04571_),
    .B1(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21oi_1 _13544_ (.A1(_04621_),
    .A2(_04570_),
    .B1(_04118_),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _13545_ (.A(\samples_imag[4][2] ),
    .B(_04580_),
    .Y(_04623_));
 sky130_fd_sc_hd__o21ai_1 _13546_ (.A1(_04595_),
    .A2(_04622_),
    .B1(_04623_),
    .Y(_00364_));
 sky130_fd_sc_hd__nor2_1 _13547_ (.A(_04121_),
    .B(_04561_),
    .Y(_04624_));
 sky130_fd_sc_hd__a21oi_1 _13548_ (.A1(\samples_imag[4][3] ),
    .A2(_04588_),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _13549_ (.A(_04564_),
    .B(_04126_),
    .Y(_04626_));
 sky130_fd_sc_hd__o21ai_1 _13550_ (.A1(_04625_),
    .A2(_04564_),
    .B1(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__a211oi_1 _13551_ (.A1(_04627_),
    .A2(_04237_),
    .B1(_04593_),
    .C1(_04130_),
    .Y(_04628_));
 sky130_fd_sc_hd__a21oi_1 _13552_ (.A1(_03398_),
    .A2(_04580_),
    .B1(_04628_),
    .Y(_00365_));
 sky130_fd_sc_hd__nor2_1 _13553_ (.A(_04133_),
    .B(_04573_),
    .Y(_04629_));
 sky130_fd_sc_hd__a21oi_1 _13554_ (.A1(\samples_imag[4][4] ),
    .A2(_04572_),
    .B1(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _13555_ (.A(_04558_),
    .B(_04138_),
    .Y(_04631_));
 sky130_fd_sc_hd__o21ai_1 _13556_ (.A1(_04630_),
    .A2(_04571_),
    .B1(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__a21oi_1 _13557_ (.A1(_04632_),
    .A2(_04570_),
    .B1(_04142_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand2_1 _13558_ (.A(\samples_imag[4][4] ),
    .B(_04580_),
    .Y(_04634_));
 sky130_fd_sc_hd__o21ai_1 _13559_ (.A1(_04595_),
    .A2(_04633_),
    .B1(_04634_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_2 _13560_ (.A(_04573_),
    .B(_04145_),
    .Y(_04635_));
 sky130_fd_sc_hd__a21oi_1 _13561_ (.A1(\samples_imag[4][5] ),
    .A2(_04572_),
    .B1(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_1 _13562_ (.A(_04558_),
    .B(_04150_),
    .Y(_04637_));
 sky130_fd_sc_hd__o21ai_1 _13563_ (.A1(_04576_),
    .A2(_04636_),
    .B1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__a21oi_1 _13564_ (.A1(_04570_),
    .A2(_04638_),
    .B1(_04154_),
    .Y(_04639_));
 sky130_fd_sc_hd__nand2_1 _13565_ (.A(\samples_imag[4][5] ),
    .B(_04580_),
    .Y(_04640_));
 sky130_fd_sc_hd__o21ai_1 _13566_ (.A1(_04639_),
    .A2(_04595_),
    .B1(_04640_),
    .Y(_00367_));
 sky130_fd_sc_hd__nor2_1 _13567_ (.A(_04573_),
    .B(_04158_),
    .Y(_04641_));
 sky130_fd_sc_hd__a21oi_1 _13568_ (.A1(\samples_imag[4][6] ),
    .A2(_04572_),
    .B1(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2_1 _13569_ (.A(_04558_),
    .B(_04162_),
    .Y(_04643_));
 sky130_fd_sc_hd__o21ai_1 _13570_ (.A1(_04576_),
    .A2(_04642_),
    .B1(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__a21oi_1 _13571_ (.A1(_04570_),
    .A2(_04644_),
    .B1(_04166_),
    .Y(_04645_));
 sky130_fd_sc_hd__clkbuf_4 _13572_ (.A(_04557_),
    .X(_04646_));
 sky130_fd_sc_hd__nand2_1 _13573_ (.A(\samples_imag[4][6] ),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_1 _13574_ (.A1(_04595_),
    .A2(_04645_),
    .B1(_04647_),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_2 _13575_ (.A(_04573_),
    .B(_04173_),
    .Y(_04648_));
 sky130_fd_sc_hd__a21oi_1 _13576_ (.A1(\samples_imag[4][7] ),
    .A2(_04572_),
    .B1(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _13577_ (.A(_04558_),
    .B(_04177_),
    .Y(_04650_));
 sky130_fd_sc_hd__o21ai_1 _13578_ (.A1(_04576_),
    .A2(_04649_),
    .B1(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__a21oi_1 _13579_ (.A1(_04570_),
    .A2(_04651_),
    .B1(_04181_),
    .Y(_04652_));
 sky130_fd_sc_hd__nand2_1 _13580_ (.A(\samples_imag[4][7] ),
    .B(_04646_),
    .Y(_04653_));
 sky130_fd_sc_hd__o21ai_1 _13581_ (.A1(_04595_),
    .A2(_04652_),
    .B1(_04653_),
    .Y(_00369_));
 sky130_fd_sc_hd__clkbuf_4 _13582_ (.A(_04170_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_4 _13583_ (.A(_04559_),
    .X(_04655_));
 sky130_fd_sc_hd__nor2_1 _13584_ (.A(_04655_),
    .B(_04186_),
    .Y(_04656_));
 sky130_fd_sc_hd__a21oi_1 _13585_ (.A1(\samples_imag[4][8] ),
    .A2(_04588_),
    .B1(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(_04558_),
    .B(_04190_),
    .Y(_04658_));
 sky130_fd_sc_hd__o21ai_1 _13587_ (.A1(_04576_),
    .A2(_04657_),
    .B1(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__a21oi_1 _13588_ (.A1(_04654_),
    .A2(_04659_),
    .B1(_04194_),
    .Y(_04660_));
 sky130_fd_sc_hd__nand2_1 _13589_ (.A(\samples_imag[4][8] ),
    .B(_04646_),
    .Y(_04661_));
 sky130_fd_sc_hd__o21ai_1 _13590_ (.A1(_04595_),
    .A2(_04660_),
    .B1(_04661_),
    .Y(_00370_));
 sky130_fd_sc_hd__nor2_1 _13591_ (.A(_04655_),
    .B(_04198_),
    .Y(_04662_));
 sky130_fd_sc_hd__a21oi_1 _13592_ (.A1(\samples_imag[4][9] ),
    .A2(_04588_),
    .B1(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_1 _13593_ (.A(_04558_),
    .B(_04202_),
    .Y(_04664_));
 sky130_fd_sc_hd__o21ai_1 _13594_ (.A1(_04576_),
    .A2(_04663_),
    .B1(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(_04654_),
    .A2(_04665_),
    .B1(_04206_),
    .Y(_04666_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(\samples_imag[4][9] ),
    .B(_04646_),
    .Y(_04667_));
 sky130_fd_sc_hd__o21ai_1 _13597_ (.A1(_04595_),
    .A2(_04666_),
    .B1(_04667_),
    .Y(_00371_));
 sky130_fd_sc_hd__and3b_1 _13598_ (.A_N(_03837_),
    .B(_03835_),
    .C(_03839_),
    .X(_04668_));
 sky130_fd_sc_hd__o21ai_4 _13599_ (.A1(_03888_),
    .A2(_04668_),
    .B1(_04210_),
    .Y(_04669_));
 sky130_fd_sc_hd__buf_2 _13600_ (.A(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_4 _13601_ (.A(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_4 _13602_ (.A(_03346_),
    .X(_04672_));
 sky130_fd_sc_hd__buf_4 _13603_ (.A(_03773_),
    .X(_04673_));
 sky130_fd_sc_hd__buf_2 _13604_ (.A(_03773_),
    .X(_04674_));
 sky130_fd_sc_hd__nor2_1 _13605_ (.A(_04674_),
    .B(_04669_),
    .Y(_04675_));
 sky130_fd_sc_hd__a22oi_1 _13606_ (.A1(\samples_imag[5][0] ),
    .A2(_04673_),
    .B1(_03994_),
    .B2(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__nor2_1 _13607_ (.A(_04672_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2b_1 _13608_ (.A_N(_03283_),
    .B(_03291_),
    .Y(_04678_));
 sky130_fd_sc_hd__clkbuf_4 _13609_ (.A(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_4 _13610_ (.A(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__nor3_2 _13611_ (.A(_04680_),
    .B(_04670_),
    .C(_03925_),
    .Y(_04681_));
 sky130_fd_sc_hd__o21ai_1 _13612_ (.A1(_04681_),
    .A2(_04677_),
    .B1(_04004_),
    .Y(_04682_));
 sky130_fd_sc_hd__clkbuf_4 _13613_ (.A(_04670_),
    .X(_04683_));
 sky130_fd_sc_hd__nand2_1 _13614_ (.A(\samples_imag[5][0] ),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__o211ai_1 _13615_ (.A1(_04001_),
    .A2(_04671_),
    .B1(_04684_),
    .C1(_04682_),
    .Y(_00372_));
 sky130_fd_sc_hd__clkbuf_4 _13616_ (.A(_04669_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_4 _13617_ (.A(_03346_),
    .X(_04686_));
 sky130_fd_sc_hd__nor2_2 _13618_ (.A(_04674_),
    .B(_04006_),
    .Y(_04687_));
 sky130_fd_sc_hd__a21oi_1 _13619_ (.A1(\samples_imag[5][10] ),
    .A2(_04673_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__buf_2 _13620_ (.A(_03346_),
    .X(_04689_));
 sky130_fd_sc_hd__nand2_1 _13621_ (.A(_04689_),
    .B(_04020_),
    .Y(_04690_));
 sky130_fd_sc_hd__o21ai_1 _13622_ (.A1(_04686_),
    .A2(_04688_),
    .B1(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__a21oi_1 _13623_ (.A1(_04654_),
    .A2(_04691_),
    .B1(_04025_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _13624_ (.A(\samples_imag[5][10] ),
    .B(_04671_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ai_1 _13625_ (.A1(_04685_),
    .A2(_04692_),
    .B1(_04693_),
    .Y(_00373_));
 sky130_fd_sc_hd__nor2_1 _13626_ (.A(_04674_),
    .B(_04031_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21oi_1 _13627_ (.A1(\samples_imag[5][11] ),
    .A2(_04673_),
    .B1(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__buf_2 _13628_ (.A(_03346_),
    .X(_04696_));
 sky130_fd_sc_hd__nand2_1 _13629_ (.A(_04696_),
    .B(_04036_),
    .Y(_04697_));
 sky130_fd_sc_hd__o21ai_1 _13630_ (.A1(_04686_),
    .A2(_04695_),
    .B1(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__a21oi_1 _13631_ (.A1(_04654_),
    .A2(_04698_),
    .B1(_04040_),
    .Y(_04699_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(\samples_imag[5][11] ),
    .B(_04671_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21ai_1 _13633_ (.A1(_04685_),
    .A2(_04699_),
    .B1(_04700_),
    .Y(_00374_));
 sky130_fd_sc_hd__nor2_1 _13634_ (.A(_03773_),
    .B(net646),
    .Y(_04701_));
 sky130_fd_sc_hd__a21oi_1 _13635_ (.A1(\samples_imag[5][12] ),
    .A2(_04674_),
    .B1(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2_1 _13636_ (.A(_03346_),
    .B(_04052_),
    .Y(_04703_));
 sky130_fd_sc_hd__o21ai_1 _13637_ (.A1(_03346_),
    .A2(_04702_),
    .B1(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__a211oi_1 _13638_ (.A1(_04704_),
    .A2(_04237_),
    .B1(_04670_),
    .C1(_04057_),
    .Y(_04705_));
 sky130_fd_sc_hd__a21oi_1 _13639_ (.A1(_03772_),
    .A2(_04671_),
    .B1(_04705_),
    .Y(_00375_));
 sky130_fd_sc_hd__buf_2 _13640_ (.A(_03773_),
    .X(_04706_));
 sky130_fd_sc_hd__nor2_1 _13641_ (.A(_04061_),
    .B(_04674_),
    .Y(_04707_));
 sky130_fd_sc_hd__a21oi_1 _13642_ (.A1(\samples_imag[5][13] ),
    .A2(_04706_),
    .B1(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _13643_ (.A(_04696_),
    .B(_04066_),
    .Y(_04709_));
 sky130_fd_sc_hd__o21ai_1 _13644_ (.A1(_04686_),
    .A2(_04708_),
    .B1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__a21oi_1 _13645_ (.A1(_04654_),
    .A2(_04710_),
    .B1(_04070_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _13646_ (.A(\samples_imag[5][13] ),
    .B(_04671_),
    .Y(_04712_));
 sky130_fd_sc_hd__o21ai_1 _13647_ (.A1(_04685_),
    .A2(_04711_),
    .B1(_04712_),
    .Y(_00376_));
 sky130_fd_sc_hd__nor2_1 _13648_ (.A(_04073_),
    .B(_04674_),
    .Y(_04713_));
 sky130_fd_sc_hd__a21oi_1 _13649_ (.A1(\samples_imag[5][14] ),
    .A2(_04706_),
    .B1(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_1 _13650_ (.A(_04696_),
    .B(_04080_),
    .Y(_04715_));
 sky130_fd_sc_hd__o21ai_1 _13651_ (.A1(_04686_),
    .A2(_04714_),
    .B1(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__a21oi_1 _13652_ (.A1(_04654_),
    .A2(_04716_),
    .B1(_04084_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(\samples_imag[5][14] ),
    .B(_04671_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21ai_1 _13654_ (.A1(_04685_),
    .A2(_04717_),
    .B1(_04718_),
    .Y(_00377_));
 sky130_fd_sc_hd__clkbuf_4 _13655_ (.A(_04670_),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_4 _13656_ (.A(_03773_),
    .X(_04720_));
 sky130_fd_sc_hd__nand2_1 _13657_ (.A(\samples_imag[5][15] ),
    .B(_03773_),
    .Y(_04721_));
 sky130_fd_sc_hd__o211ai_1 _13658_ (.A1(_04720_),
    .A2(_04090_),
    .B1(_04721_),
    .C1(_04679_),
    .Y(_04722_));
 sky130_fd_sc_hd__o21ai_0 _13659_ (.A1(_04679_),
    .A2(net525),
    .B1(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__a211oi_1 _13660_ (.A1(_04088_),
    .A2(_04723_),
    .B1(_04670_),
    .C1(_04095_),
    .Y(_04724_));
 sky130_fd_sc_hd__a21o_1 _13661_ (.A1(\samples_imag[5][15] ),
    .A2(_04719_),
    .B1(_04724_),
    .X(_00378_));
 sky130_fd_sc_hd__nor2_1 _13662_ (.A(_04674_),
    .B(_04097_),
    .Y(_04725_));
 sky130_fd_sc_hd__a21oi_1 _13663_ (.A1(\samples_imag[5][1] ),
    .A2(_04706_),
    .B1(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_1 _13664_ (.A(_04101_),
    .B(_04696_),
    .Y(_04727_));
 sky130_fd_sc_hd__o21ai_1 _13665_ (.A1(_04686_),
    .A2(_04726_),
    .B1(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__a21oi_1 _13666_ (.A1(_04654_),
    .A2(_04728_),
    .B1(_04105_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(\samples_imag[5][1] ),
    .B(_04671_),
    .Y(_04730_));
 sky130_fd_sc_hd__o21ai_1 _13668_ (.A1(_04685_),
    .A2(_04729_),
    .B1(_04730_),
    .Y(_00379_));
 sky130_fd_sc_hd__nor2_1 _13669_ (.A(_04109_),
    .B(_04674_),
    .Y(_04731_));
 sky130_fd_sc_hd__a21oi_1 _13670_ (.A1(\samples_imag[5][2] ),
    .A2(_04706_),
    .B1(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__nand2_1 _13671_ (.A(_04696_),
    .B(_04114_),
    .Y(_04733_));
 sky130_fd_sc_hd__o21ai_1 _13672_ (.A1(_04689_),
    .A2(_04732_),
    .B1(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__a21oi_1 _13673_ (.A1(_04654_),
    .A2(_04734_),
    .B1(_04118_),
    .Y(_04735_));
 sky130_fd_sc_hd__nand2_1 _13674_ (.A(\samples_imag[5][2] ),
    .B(_04671_),
    .Y(_04736_));
 sky130_fd_sc_hd__o21ai_1 _13675_ (.A1(_04685_),
    .A2(_04735_),
    .B1(_04736_),
    .Y(_00380_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(_04121_),
    .B(_04720_),
    .Y(_04737_));
 sky130_fd_sc_hd__a21oi_1 _13677_ (.A1(\samples_imag[5][3] ),
    .A2(_04706_),
    .B1(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand2_1 _13678_ (.A(_04696_),
    .B(_04126_),
    .Y(_04739_));
 sky130_fd_sc_hd__o21ai_1 _13679_ (.A1(_04689_),
    .A2(_04738_),
    .B1(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__a21oi_1 _13680_ (.A1(_04654_),
    .A2(_04740_),
    .B1(_04130_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(\samples_imag[5][3] ),
    .B(_04671_),
    .Y(_04742_));
 sky130_fd_sc_hd__o21ai_1 _13682_ (.A1(_04685_),
    .A2(_04741_),
    .B1(_04742_),
    .Y(_00381_));
 sky130_fd_sc_hd__nor2_1 _13683_ (.A(_04133_),
    .B(_04720_),
    .Y(_04743_));
 sky130_fd_sc_hd__a21oi_1 _13684_ (.A1(\samples_imag[5][4] ),
    .A2(_04706_),
    .B1(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(_04696_),
    .B(_04138_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21ai_1 _13686_ (.A1(_04689_),
    .A2(_04744_),
    .B1(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__a21oi_1 _13687_ (.A1(_04654_),
    .A2(_04746_),
    .B1(_04142_),
    .Y(_04747_));
 sky130_fd_sc_hd__nand2_1 _13688_ (.A(\samples_imag[5][4] ),
    .B(_04671_),
    .Y(_04748_));
 sky130_fd_sc_hd__o21ai_1 _13689_ (.A1(_04685_),
    .A2(_04747_),
    .B1(_04748_),
    .Y(_00382_));
 sky130_fd_sc_hd__clkbuf_4 _13690_ (.A(_04170_),
    .X(_04749_));
 sky130_fd_sc_hd__nor2_1 _13691_ (.A(_04145_),
    .B(_04720_),
    .Y(_04750_));
 sky130_fd_sc_hd__a21oi_1 _13692_ (.A1(\samples_imag[5][5] ),
    .A2(_04706_),
    .B1(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_1 _13693_ (.A(_04696_),
    .B(_04150_),
    .Y(_04752_));
 sky130_fd_sc_hd__o21ai_1 _13694_ (.A1(_04689_),
    .A2(_04751_),
    .B1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__a21oi_1 _13695_ (.A1(_04749_),
    .A2(_04753_),
    .B1(_04154_),
    .Y(_04754_));
 sky130_fd_sc_hd__clkbuf_4 _13696_ (.A(_04670_),
    .X(_04755_));
 sky130_fd_sc_hd__nand2_1 _13697_ (.A(\samples_imag[5][5] ),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__o21ai_1 _13698_ (.A1(_04685_),
    .A2(_04754_),
    .B1(_04756_),
    .Y(_00383_));
 sky130_fd_sc_hd__buf_2 _13699_ (.A(_04669_),
    .X(_04757_));
 sky130_fd_sc_hd__nor2_1 _13700_ (.A(_04720_),
    .B(_04158_),
    .Y(_04758_));
 sky130_fd_sc_hd__a21oi_1 _13701_ (.A1(\samples_imag[5][6] ),
    .A2(_04706_),
    .B1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _13702_ (.A(_04696_),
    .B(_04162_),
    .Y(_04760_));
 sky130_fd_sc_hd__o21ai_1 _13703_ (.A1(_04689_),
    .A2(_04759_),
    .B1(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__a21oi_1 _13704_ (.A1(_04749_),
    .A2(_04761_),
    .B1(_04166_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand2_1 _13705_ (.A(\samples_imag[5][6] ),
    .B(_04755_),
    .Y(_04763_));
 sky130_fd_sc_hd__o21ai_1 _13706_ (.A1(_04757_),
    .A2(_04762_),
    .B1(_04763_),
    .Y(_00384_));
 sky130_fd_sc_hd__nor2_1 _13707_ (.A(_04720_),
    .B(_04173_),
    .Y(_04764_));
 sky130_fd_sc_hd__a21oi_1 _13708_ (.A1(\samples_imag[5][7] ),
    .A2(_04706_),
    .B1(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _13709_ (.A(_04696_),
    .B(_04177_),
    .Y(_04766_));
 sky130_fd_sc_hd__o21ai_1 _13710_ (.A1(_04689_),
    .A2(_04765_),
    .B1(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__a21oi_1 _13711_ (.A1(_04749_),
    .A2(_04767_),
    .B1(_04181_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2_1 _13712_ (.A(\samples_imag[5][7] ),
    .B(_04755_),
    .Y(_04769_));
 sky130_fd_sc_hd__o21ai_1 _13713_ (.A1(_04757_),
    .A2(_04768_),
    .B1(_04769_),
    .Y(_00385_));
 sky130_fd_sc_hd__nor2_1 _13714_ (.A(_04720_),
    .B(_04186_),
    .Y(_04770_));
 sky130_fd_sc_hd__a21oi_1 _13715_ (.A1(\samples_imag[5][8] ),
    .A2(_04706_),
    .B1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_1 _13716_ (.A(_03346_),
    .B(_04190_),
    .Y(_04772_));
 sky130_fd_sc_hd__o21ai_1 _13717_ (.A1(_04689_),
    .A2(_04771_),
    .B1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__a21oi_1 _13718_ (.A1(_04749_),
    .A2(_04773_),
    .B1(_04194_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _13719_ (.A(\samples_imag[5][8] ),
    .B(_04755_),
    .Y(_04775_));
 sky130_fd_sc_hd__o21ai_1 _13720_ (.A1(_04757_),
    .A2(_04774_),
    .B1(_04775_),
    .Y(_00386_));
 sky130_fd_sc_hd__nor2_2 _13721_ (.A(_04720_),
    .B(_04198_),
    .Y(_04776_));
 sky130_fd_sc_hd__a21oi_1 _13722_ (.A1(\samples_imag[5][9] ),
    .A2(_04674_),
    .B1(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_1 _13723_ (.A(_03346_),
    .B(_04202_),
    .Y(_04778_));
 sky130_fd_sc_hd__o21ai_1 _13724_ (.A1(_04689_),
    .A2(_04777_),
    .B1(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__a21oi_1 _13725_ (.A1(_04749_),
    .A2(_04779_),
    .B1(_04206_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _13726_ (.A(\samples_imag[5][9] ),
    .B(_04755_),
    .Y(_04781_));
 sky130_fd_sc_hd__o21ai_1 _13727_ (.A1(_04757_),
    .A2(_04780_),
    .B1(_04781_),
    .Y(_00387_));
 sky130_fd_sc_hd__and3b_1 _13728_ (.A_N(_03835_),
    .B(_03839_),
    .C(_03837_),
    .X(_04782_));
 sky130_fd_sc_hd__o21ai_1 _13729_ (.A1(_03888_),
    .A2(_04782_),
    .B1(_04210_),
    .Y(_04783_));
 sky130_fd_sc_hd__clkbuf_4 _13730_ (.A(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__nand2_4 _13731_ (.A(_03147_),
    .B(net614),
    .Y(_04785_));
 sky130_fd_sc_hd__clkbuf_4 _13732_ (.A(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__nor2_1 _13733_ (.A(_04785_),
    .B(_04784_),
    .Y(_04787_));
 sky130_fd_sc_hd__a22oi_2 _13734_ (.A1(\samples_imag[6][0] ),
    .A2(_04786_),
    .B1(_04787_),
    .B2(_03994_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand2b_1 _13735_ (.A_N(net45),
    .B(_03316_),
    .Y(_04789_));
 sky130_fd_sc_hd__buf_2 _13736_ (.A(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__or2_0 _13737_ (.A(_04790_),
    .B(_04784_),
    .X(_04791_));
 sky130_fd_sc_hd__o22ai_2 _13738_ (.A1(_03676_),
    .A2(_04788_),
    .B1(_04791_),
    .B2(_03925_),
    .Y(_04792_));
 sky130_fd_sc_hd__nor2_1 _13739_ (.A(_04001_),
    .B(_04784_),
    .Y(_04793_));
 sky130_fd_sc_hd__a221o_1 _13740_ (.A1(\samples_imag[6][0] ),
    .A2(_04784_),
    .B1(_04792_),
    .B2(_03999_),
    .C1(_04793_),
    .X(_00388_));
 sky130_fd_sc_hd__buf_4 _13741_ (.A(_04784_),
    .X(_04794_));
 sky130_fd_sc_hd__clkbuf_4 _13742_ (.A(_03676_),
    .X(_04795_));
 sky130_fd_sc_hd__buf_4 _13743_ (.A(_04785_),
    .X(_04796_));
 sky130_fd_sc_hd__clkbuf_4 _13744_ (.A(_04785_),
    .X(_04797_));
 sky130_fd_sc_hd__nor2_2 _13745_ (.A(_04006_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__a21oi_1 _13746_ (.A1(\samples_imag[6][10] ),
    .A2(_04796_),
    .B1(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__clkbuf_4 _13747_ (.A(_03676_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _13748_ (.A(_04800_),
    .B(_04020_),
    .Y(_04801_));
 sky130_fd_sc_hd__o21ai_1 _13749_ (.A1(_04795_),
    .A2(_04799_),
    .B1(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_1 _13750_ (.A1(_04749_),
    .A2(_04802_),
    .B1(_04025_),
    .Y(_04803_));
 sky130_fd_sc_hd__buf_2 _13751_ (.A(_04784_),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _13752_ (.A(\samples_imag[6][10] ),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__o21ai_1 _13753_ (.A1(_04794_),
    .A2(_04803_),
    .B1(_04805_),
    .Y(_00389_));
 sky130_fd_sc_hd__nor2_1 _13754_ (.A(_04031_),
    .B(_04797_),
    .Y(_04806_));
 sky130_fd_sc_hd__a21oi_1 _13755_ (.A1(\samples_imag[6][11] ),
    .A2(_04796_),
    .B1(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__buf_2 _13756_ (.A(_03676_),
    .X(_04808_));
 sky130_fd_sc_hd__nand2_1 _13757_ (.A(_04808_),
    .B(_04036_),
    .Y(_04809_));
 sky130_fd_sc_hd__o21ai_1 _13758_ (.A1(_04795_),
    .A2(_04807_),
    .B1(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__a21oi_1 _13759_ (.A1(_04749_),
    .A2(_04810_),
    .B1(_04040_),
    .Y(_04811_));
 sky130_fd_sc_hd__nand2_1 _13760_ (.A(\samples_imag[6][11] ),
    .B(_04804_),
    .Y(_04812_));
 sky130_fd_sc_hd__o21ai_1 _13761_ (.A1(_04794_),
    .A2(_04811_),
    .B1(_04812_),
    .Y(_00390_));
 sky130_fd_sc_hd__clkbuf_2 _13762_ (.A(_04783_),
    .X(_04813_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_04045_),
    .B(_04797_),
    .Y(_04814_));
 sky130_fd_sc_hd__a21oi_1 _13764_ (.A1(\samples_imag[6][12] ),
    .A2(_04796_),
    .B1(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _13765_ (.A(_04808_),
    .B(_04052_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_1 _13766_ (.A1(_04795_),
    .A2(_04815_),
    .B1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__a21oi_1 _13767_ (.A1(_04749_),
    .A2(_04817_),
    .B1(_04057_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand2_1 _13768_ (.A(\samples_imag[6][12] ),
    .B(_04804_),
    .Y(_04819_));
 sky130_fd_sc_hd__o21ai_1 _13769_ (.A1(_04818_),
    .A2(_04813_),
    .B1(_04819_),
    .Y(_00391_));
 sky130_fd_sc_hd__nor2_1 _13770_ (.A(_04061_),
    .B(_04797_),
    .Y(_04820_));
 sky130_fd_sc_hd__a21oi_1 _13771_ (.A1(\samples_imag[6][13] ),
    .A2(_04796_),
    .B1(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _13772_ (.A(_04808_),
    .B(_04066_),
    .Y(_04822_));
 sky130_fd_sc_hd__o21ai_1 _13773_ (.A1(_04795_),
    .A2(_04821_),
    .B1(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__a21oi_1 _13774_ (.A1(_04749_),
    .A2(_04823_),
    .B1(_04070_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand2_1 _13775_ (.A(\samples_imag[6][13] ),
    .B(_04804_),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ai_1 _13776_ (.A1(_04813_),
    .A2(_04824_),
    .B1(_04825_),
    .Y(_00392_));
 sky130_fd_sc_hd__buf_2 _13777_ (.A(_04785_),
    .X(_04826_));
 sky130_fd_sc_hd__nor2_1 _13778_ (.A(_04073_),
    .B(_04797_),
    .Y(_04827_));
 sky130_fd_sc_hd__a21oi_1 _13779_ (.A1(\samples_imag[6][14] ),
    .A2(_04826_),
    .B1(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_04808_),
    .B(_04080_),
    .Y(_04829_));
 sky130_fd_sc_hd__o21ai_1 _13781_ (.A1(_04795_),
    .A2(_04828_),
    .B1(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__a21oi_1 _13782_ (.A1(_04749_),
    .A2(_04830_),
    .B1(_04084_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand2_1 _13783_ (.A(\samples_imag[6][14] ),
    .B(_04804_),
    .Y(_04832_));
 sky130_fd_sc_hd__o21ai_1 _13784_ (.A1(_04813_),
    .A2(_04831_),
    .B1(_04832_),
    .Y(_00393_));
 sky130_fd_sc_hd__clkbuf_4 _13785_ (.A(_04784_),
    .X(_04833_));
 sky130_fd_sc_hd__nand2_1 _13786_ (.A(\samples_imag[6][15] ),
    .B(_04785_),
    .Y(_04834_));
 sky130_fd_sc_hd__o211ai_1 _13787_ (.A1(_04090_),
    .A2(_04797_),
    .B1(_04834_),
    .C1(_04790_),
    .Y(_04835_));
 sky130_fd_sc_hd__o21ai_0 _13788_ (.A1(_04790_),
    .A2(net525),
    .B1(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__a211oi_1 _13789_ (.A1(_04088_),
    .A2(_04836_),
    .B1(_04833_),
    .C1(_04095_),
    .Y(_04837_));
 sky130_fd_sc_hd__a21o_1 _13790_ (.A1(\samples_imag[6][15] ),
    .A2(_04833_),
    .B1(_04837_),
    .X(_00394_));
 sky130_fd_sc_hd__buf_2 _13791_ (.A(_04170_),
    .X(_04838_));
 sky130_fd_sc_hd__nor2_1 _13792_ (.A(_04097_),
    .B(_04797_),
    .Y(_04839_));
 sky130_fd_sc_hd__a21oi_1 _13793_ (.A1(\samples_imag[6][1] ),
    .A2(_04826_),
    .B1(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_1 _13794_ (.A(_04808_),
    .B(_04101_),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_1 _13795_ (.A1(_04795_),
    .A2(_04840_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__a21oi_1 _13796_ (.A1(_04838_),
    .A2(_04842_),
    .B1(_04105_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _13797_ (.A(\samples_imag[6][1] ),
    .B(_04804_),
    .Y(_04844_));
 sky130_fd_sc_hd__o21ai_1 _13798_ (.A1(_04813_),
    .A2(_04843_),
    .B1(_04844_),
    .Y(_00395_));
 sky130_fd_sc_hd__nor2_1 _13799_ (.A(_04797_),
    .B(_04109_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21oi_1 _13800_ (.A1(\samples_imag[6][2] ),
    .A2(_04826_),
    .B1(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _13801_ (.A(_04808_),
    .B(_04114_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21ai_1 _13802_ (.A1(_04800_),
    .A2(_04846_),
    .B1(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21oi_1 _13803_ (.A1(_04838_),
    .A2(_04848_),
    .B1(_04118_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _13804_ (.A(\samples_imag[6][2] ),
    .B(_04804_),
    .Y(_04850_));
 sky130_fd_sc_hd__o21ai_1 _13805_ (.A1(_04813_),
    .A2(_04849_),
    .B1(_04850_),
    .Y(_00396_));
 sky130_fd_sc_hd__nor2_2 _13806_ (.A(_04121_),
    .B(_04786_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_1 _13807_ (.A1(\samples_imag[6][3] ),
    .A2(_04826_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(_04808_),
    .B(_04126_),
    .Y(_04853_));
 sky130_fd_sc_hd__o21ai_1 _13809_ (.A1(_04800_),
    .A2(_04852_),
    .B1(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__a21oi_1 _13810_ (.A1(_04838_),
    .A2(_04854_),
    .B1(_04130_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _13811_ (.A(\samples_imag[6][3] ),
    .B(_04804_),
    .Y(_04856_));
 sky130_fd_sc_hd__o21ai_1 _13812_ (.A1(_04813_),
    .A2(_04855_),
    .B1(_04856_),
    .Y(_00397_));
 sky130_fd_sc_hd__nor2_1 _13813_ (.A(_04786_),
    .B(_04133_),
    .Y(_04857_));
 sky130_fd_sc_hd__a21oi_1 _13814_ (.A1(\samples_imag[6][4] ),
    .A2(_04826_),
    .B1(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _13815_ (.A(_04808_),
    .B(_04138_),
    .Y(_04859_));
 sky130_fd_sc_hd__o21ai_1 _13816_ (.A1(_04800_),
    .A2(_04858_),
    .B1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__a21oi_1 _13817_ (.A1(_04838_),
    .A2(_04860_),
    .B1(_04142_),
    .Y(_04861_));
 sky130_fd_sc_hd__nand2_1 _13818_ (.A(\samples_imag[6][4] ),
    .B(_04804_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21ai_1 _13819_ (.A1(_04813_),
    .A2(_04861_),
    .B1(_04862_),
    .Y(_00398_));
 sky130_fd_sc_hd__nor2_1 _13820_ (.A(_04786_),
    .B(_04145_),
    .Y(_04863_));
 sky130_fd_sc_hd__a21oi_1 _13821_ (.A1(\samples_imag[6][5] ),
    .A2(_04826_),
    .B1(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_1 _13822_ (.A(_04808_),
    .B(_04150_),
    .Y(_04865_));
 sky130_fd_sc_hd__o21ai_1 _13823_ (.A1(_04800_),
    .A2(_04864_),
    .B1(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__a21oi_1 _13824_ (.A1(_04838_),
    .A2(_04866_),
    .B1(_04154_),
    .Y(_04867_));
 sky130_fd_sc_hd__nand2_1 _13825_ (.A(\samples_imag[6][5] ),
    .B(_04804_),
    .Y(_04868_));
 sky130_fd_sc_hd__o21ai_1 _13826_ (.A1(_04813_),
    .A2(_04867_),
    .B1(_04868_),
    .Y(_00399_));
 sky130_fd_sc_hd__nor2_1 _13827_ (.A(_04158_),
    .B(_04786_),
    .Y(_04869_));
 sky130_fd_sc_hd__a21oi_1 _13828_ (.A1(\samples_imag[6][6] ),
    .A2(_04826_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(_04808_),
    .B(_04162_),
    .Y(_04871_));
 sky130_fd_sc_hd__o21ai_1 _13830_ (.A1(_04800_),
    .A2(_04870_),
    .B1(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21oi_1 _13831_ (.A1(_04838_),
    .A2(_04872_),
    .B1(_04166_),
    .Y(_04873_));
 sky130_fd_sc_hd__buf_4 _13832_ (.A(_04784_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _13833_ (.A(\samples_imag[6][6] ),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_1 _13834_ (.A1(_04813_),
    .A2(_04873_),
    .B1(_04875_),
    .Y(_00400_));
 sky130_fd_sc_hd__nor2_2 _13835_ (.A(_04173_),
    .B(_04786_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_1 _13836_ (.A1(\samples_imag[6][7] ),
    .A2(_04826_),
    .B1(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_1 _13837_ (.A(_03676_),
    .B(_04177_),
    .Y(_04878_));
 sky130_fd_sc_hd__o21ai_1 _13838_ (.A1(_04800_),
    .A2(_04877_),
    .B1(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21oi_1 _13839_ (.A1(_04838_),
    .A2(_04879_),
    .B1(_04181_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _13840_ (.A(\samples_imag[6][7] ),
    .B(_04874_),
    .Y(_04881_));
 sky130_fd_sc_hd__o21ai_1 _13841_ (.A1(_04813_),
    .A2(_04880_),
    .B1(_04881_),
    .Y(_00401_));
 sky130_fd_sc_hd__buf_4 _13842_ (.A(_04783_),
    .X(_04882_));
 sky130_fd_sc_hd__nor2_1 _13843_ (.A(_04186_),
    .B(_04786_),
    .Y(_04883_));
 sky130_fd_sc_hd__a21oi_1 _13844_ (.A1(\samples_imag[6][8] ),
    .A2(_04826_),
    .B1(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_1 _13845_ (.A(_03676_),
    .B(_04190_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_1 _13846_ (.A1(_04800_),
    .A2(_04884_),
    .B1(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_1 _13847_ (.A1(_04838_),
    .A2(_04886_),
    .B1(_04194_),
    .Y(_04887_));
 sky130_fd_sc_hd__nand2_1 _13848_ (.A(\samples_imag[6][8] ),
    .B(_04874_),
    .Y(_04888_));
 sky130_fd_sc_hd__o21ai_1 _13849_ (.A1(_04882_),
    .A2(_04887_),
    .B1(_04888_),
    .Y(_00402_));
 sky130_fd_sc_hd__nor2_2 _13850_ (.A(_04198_),
    .B(_04786_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21oi_1 _13851_ (.A1(\samples_imag[6][9] ),
    .A2(_04826_),
    .B1(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_1 _13852_ (.A(_03676_),
    .B(_04202_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_1 _13853_ (.A1(_04800_),
    .A2(_04890_),
    .B1(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21oi_1 _13854_ (.A1(_04838_),
    .A2(_04892_),
    .B1(_04206_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(\samples_imag[6][9] ),
    .B(_04874_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21ai_1 _13856_ (.A1(_04882_),
    .A2(_04893_),
    .B1(_04894_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand3_1 _13857_ (.A(_03837_),
    .B(_03835_),
    .C(_03839_),
    .Y(_04895_));
 sky130_fd_sc_hd__a21oi_1 _13858_ (.A1(net91),
    .A2(_04895_),
    .B1(_03887_),
    .Y(_04896_));
 sky130_fd_sc_hd__o21ai_2 _13859_ (.A1(_03140_),
    .A2(_04896_),
    .B1(_03891_),
    .Y(_04897_));
 sky130_fd_sc_hd__clkbuf_4 _13860_ (.A(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__clkbuf_4 _13861_ (.A(_03268_),
    .X(_04899_));
 sky130_fd_sc_hd__nand3_4 _13862_ (.A(_03147_),
    .B(net55),
    .C(net642),
    .Y(_04900_));
 sky130_fd_sc_hd__clkbuf_4 _13863_ (.A(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__nor2_1 _13864_ (.A(_04900_),
    .B(_04898_),
    .Y(_04902_));
 sky130_fd_sc_hd__a22oi_1 _13865_ (.A1(\samples_imag[7][0] ),
    .A2(_04901_),
    .B1(_03994_),
    .B2(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_2 _13866_ (.A(_03296_),
    .B(_03291_),
    .Y(_04904_));
 sky130_fd_sc_hd__or2_0 _13867_ (.A(_04904_),
    .B(_04898_),
    .X(_04905_));
 sky130_fd_sc_hd__o22ai_2 _13868_ (.A1(_04899_),
    .A2(_04903_),
    .B1(_04905_),
    .B2(_03925_),
    .Y(_04906_));
 sky130_fd_sc_hd__nor2_1 _13869_ (.A(_04001_),
    .B(_04898_),
    .Y(_04907_));
 sky130_fd_sc_hd__a221o_1 _13870_ (.A1(\samples_imag[7][0] ),
    .A2(_04898_),
    .B1(_04906_),
    .B2(_03999_),
    .C1(_04907_),
    .X(_00404_));
 sky130_fd_sc_hd__buf_4 _13871_ (.A(_04898_),
    .X(_04908_));
 sky130_fd_sc_hd__buf_2 _13872_ (.A(_03268_),
    .X(_04909_));
 sky130_fd_sc_hd__buf_4 _13873_ (.A(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_2 _13874_ (.A(_04900_),
    .X(_04911_));
 sky130_fd_sc_hd__buf_2 _13875_ (.A(_04900_),
    .X(_04912_));
 sky130_fd_sc_hd__nor2_1 _13876_ (.A(_04006_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__a21oi_1 _13877_ (.A1(\samples_imag[7][10] ),
    .A2(_04911_),
    .B1(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__buf_2 _13878_ (.A(_03268_),
    .X(_04915_));
 sky130_fd_sc_hd__nand2_1 _13879_ (.A(_04915_),
    .B(_04020_),
    .Y(_04916_));
 sky130_fd_sc_hd__o21ai_1 _13880_ (.A1(_04910_),
    .A2(_04914_),
    .B1(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__a21oi_1 _13881_ (.A1(_04838_),
    .A2(_04917_),
    .B1(_04025_),
    .Y(_04918_));
 sky130_fd_sc_hd__buf_2 _13882_ (.A(_04898_),
    .X(_04919_));
 sky130_fd_sc_hd__nand2_1 _13883_ (.A(\samples_imag[7][10] ),
    .B(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__o21ai_1 _13884_ (.A1(_04908_),
    .A2(_04918_),
    .B1(_04920_),
    .Y(_00405_));
 sky130_fd_sc_hd__buf_2 _13885_ (.A(_04170_),
    .X(_04921_));
 sky130_fd_sc_hd__nor2_2 _13886_ (.A(_04031_),
    .B(_04912_),
    .Y(_04922_));
 sky130_fd_sc_hd__a21oi_1 _13887_ (.A1(\samples_imag[7][11] ),
    .A2(_04911_),
    .B1(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__buf_2 _13888_ (.A(_03268_),
    .X(_04924_));
 sky130_fd_sc_hd__nand2_1 _13889_ (.A(_04924_),
    .B(_04036_),
    .Y(_04925_));
 sky130_fd_sc_hd__o21ai_1 _13890_ (.A1(_04910_),
    .A2(_04923_),
    .B1(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__a21oi_1 _13891_ (.A1(_04921_),
    .A2(_04926_),
    .B1(_04040_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2_1 _13892_ (.A(\samples_imag[7][11] ),
    .B(_04919_),
    .Y(_04928_));
 sky130_fd_sc_hd__o21ai_1 _13893_ (.A1(_04908_),
    .A2(_04927_),
    .B1(_04928_),
    .Y(_00406_));
 sky130_fd_sc_hd__buf_2 _13894_ (.A(_04897_),
    .X(_04929_));
 sky130_fd_sc_hd__nor2_2 _13895_ (.A(_04912_),
    .B(net646),
    .Y(_04930_));
 sky130_fd_sc_hd__a21oi_1 _13896_ (.A1(\samples_imag[7][12] ),
    .A2(_04911_),
    .B1(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand2_1 _13897_ (.A(_04924_),
    .B(_04052_),
    .Y(_04932_));
 sky130_fd_sc_hd__o21ai_1 _13898_ (.A1(_04910_),
    .A2(_04931_),
    .B1(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__a21oi_1 _13899_ (.A1(_04921_),
    .A2(_04933_),
    .B1(_04057_),
    .Y(_04934_));
 sky130_fd_sc_hd__nand2_1 _13900_ (.A(\samples_imag[7][12] ),
    .B(_04919_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21ai_1 _13901_ (.A1(_04929_),
    .A2(_04934_),
    .B1(_04935_),
    .Y(_00407_));
 sky130_fd_sc_hd__nor2_1 _13902_ (.A(_04912_),
    .B(_04061_),
    .Y(_04936_));
 sky130_fd_sc_hd__a21oi_1 _13903_ (.A1(\samples_imag[7][13] ),
    .A2(_04911_),
    .B1(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2_1 _13904_ (.A(_04924_),
    .B(_04066_),
    .Y(_04938_));
 sky130_fd_sc_hd__o21ai_1 _13905_ (.A1(_04910_),
    .A2(_04937_),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__a21oi_1 _13906_ (.A1(_04921_),
    .A2(_04939_),
    .B1(_04070_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(\samples_imag[7][13] ),
    .B(_04919_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21ai_1 _13908_ (.A1(_04929_),
    .A2(_04940_),
    .B1(_04941_),
    .Y(_00408_));
 sky130_fd_sc_hd__nor2_1 _13909_ (.A(_04912_),
    .B(_04073_),
    .Y(_04942_));
 sky130_fd_sc_hd__a21oi_1 _13910_ (.A1(\samples_imag[7][14] ),
    .A2(_04911_),
    .B1(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_04924_),
    .B(_04080_),
    .Y(_04944_));
 sky130_fd_sc_hd__o21ai_1 _13912_ (.A1(_04910_),
    .A2(_04943_),
    .B1(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__a21oi_1 _13913_ (.A1(_04921_),
    .A2(_04945_),
    .B1(_04084_),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2_1 _13914_ (.A(\samples_imag[7][14] ),
    .B(_04919_),
    .Y(_04947_));
 sky130_fd_sc_hd__o21ai_1 _13915_ (.A1(_04929_),
    .A2(_04946_),
    .B1(_04947_),
    .Y(_00409_));
 sky130_fd_sc_hd__clkbuf_4 _13916_ (.A(_04898_),
    .X(_04948_));
 sky130_fd_sc_hd__buf_4 _13917_ (.A(_04900_),
    .X(_04949_));
 sky130_fd_sc_hd__nand2_1 _13918_ (.A(\samples_imag[7][15] ),
    .B(_04900_),
    .Y(_04950_));
 sky130_fd_sc_hd__o211ai_1 _13919_ (.A1(_04949_),
    .A2(_04090_),
    .B1(_04950_),
    .C1(_04904_),
    .Y(_04951_));
 sky130_fd_sc_hd__o21ai_0 _13920_ (.A1(_04904_),
    .A2(net54),
    .B1(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__a211oi_1 _13921_ (.A1(_04029_),
    .A2(_04952_),
    .B1(_04948_),
    .C1(_04095_),
    .Y(_04953_));
 sky130_fd_sc_hd__a21o_1 _13922_ (.A1(\samples_imag[7][15] ),
    .A2(_04948_),
    .B1(_04953_),
    .X(_00410_));
 sky130_fd_sc_hd__nor2_1 _13923_ (.A(_04912_),
    .B(_04097_),
    .Y(_04954_));
 sky130_fd_sc_hd__a21oi_1 _13924_ (.A1(\samples_imag[7][1] ),
    .A2(_04911_),
    .B1(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _13925_ (.A(_04101_),
    .B(_04924_),
    .Y(_04956_));
 sky130_fd_sc_hd__o21ai_1 _13926_ (.A1(_04910_),
    .A2(_04955_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__a21oi_1 _13927_ (.A1(_04921_),
    .A2(_04957_),
    .B1(_04105_),
    .Y(_04958_));
 sky130_fd_sc_hd__nand2_1 _13928_ (.A(\samples_imag[7][1] ),
    .B(_04919_),
    .Y(_04959_));
 sky130_fd_sc_hd__o21ai_1 _13929_ (.A1(_04929_),
    .A2(_04958_),
    .B1(_04959_),
    .Y(_00411_));
 sky130_fd_sc_hd__nor2_2 _13930_ (.A(_04109_),
    .B(_04912_),
    .Y(_04960_));
 sky130_fd_sc_hd__a21oi_1 _13931_ (.A1(\samples_imag[7][2] ),
    .A2(_04911_),
    .B1(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand2_1 _13932_ (.A(_04924_),
    .B(_04114_),
    .Y(_04962_));
 sky130_fd_sc_hd__o21ai_1 _13933_ (.A1(_04915_),
    .A2(_04961_),
    .B1(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__a21oi_1 _13934_ (.A1(_04921_),
    .A2(_04963_),
    .B1(_04118_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand2_1 _13935_ (.A(\samples_imag[7][2] ),
    .B(_04919_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21ai_1 _13936_ (.A1(_04929_),
    .A2(_04964_),
    .B1(_04965_),
    .Y(_00412_));
 sky130_fd_sc_hd__nor2_1 _13937_ (.A(_04121_),
    .B(_04912_),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_1 _13938_ (.A1(\samples_imag[7][3] ),
    .A2(_04911_),
    .B1(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nand2_1 _13939_ (.A(_04924_),
    .B(_04126_),
    .Y(_04968_));
 sky130_fd_sc_hd__o21ai_1 _13940_ (.A1(_04915_),
    .A2(_04967_),
    .B1(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__a21oi_1 _13941_ (.A1(_04921_),
    .A2(_04969_),
    .B1(_04130_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_1 _13942_ (.A(\samples_imag[7][3] ),
    .B(_04919_),
    .Y(_04971_));
 sky130_fd_sc_hd__o21ai_1 _13943_ (.A1(_04929_),
    .A2(_04970_),
    .B1(_04971_),
    .Y(_00413_));
 sky130_fd_sc_hd__nor2_1 _13944_ (.A(_04133_),
    .B(_04912_),
    .Y(_04972_));
 sky130_fd_sc_hd__a21oi_1 _13945_ (.A1(\samples_imag[7][4] ),
    .A2(_04911_),
    .B1(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_1 _13946_ (.A(_04924_),
    .B(_04138_),
    .Y(_04974_));
 sky130_fd_sc_hd__o21ai_1 _13947_ (.A1(_04915_),
    .A2(_04973_),
    .B1(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__a21oi_1 _13948_ (.A1(_04921_),
    .A2(_04975_),
    .B1(_04142_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _13949_ (.A(\samples_imag[7][4] ),
    .B(_04919_),
    .Y(_04977_));
 sky130_fd_sc_hd__o21ai_1 _13950_ (.A1(_04929_),
    .A2(_04976_),
    .B1(_04977_),
    .Y(_00414_));
 sky130_fd_sc_hd__nor2_1 _13951_ (.A(_04145_),
    .B(_04912_),
    .Y(_04978_));
 sky130_fd_sc_hd__a21oi_1 _13952_ (.A1(\samples_imag[7][5] ),
    .A2(_04911_),
    .B1(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _13953_ (.A(_04924_),
    .B(_04150_),
    .Y(_04980_));
 sky130_fd_sc_hd__o21ai_1 _13954_ (.A1(_04915_),
    .A2(_04979_),
    .B1(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__a21oi_1 _13955_ (.A1(_04921_),
    .A2(_04981_),
    .B1(_04154_),
    .Y(_04982_));
 sky130_fd_sc_hd__nand2_1 _13956_ (.A(\samples_imag[7][5] ),
    .B(_04919_),
    .Y(_04983_));
 sky130_fd_sc_hd__o21ai_1 _13957_ (.A1(_04929_),
    .A2(_04982_),
    .B1(_04983_),
    .Y(_00415_));
 sky130_fd_sc_hd__clkbuf_4 _13958_ (.A(_04900_),
    .X(_04984_));
 sky130_fd_sc_hd__nor2_2 _13959_ (.A(_04949_),
    .B(_04158_),
    .Y(_04985_));
 sky130_fd_sc_hd__a21oi_1 _13960_ (.A1(\samples_imag[7][6] ),
    .A2(_04984_),
    .B1(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _13961_ (.A(_04924_),
    .B(_04162_),
    .Y(_04987_));
 sky130_fd_sc_hd__o21ai_1 _13962_ (.A1(_04915_),
    .A2(_04986_),
    .B1(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__a21oi_1 _13963_ (.A1(_04921_),
    .A2(_04988_),
    .B1(_04166_),
    .Y(_04989_));
 sky130_fd_sc_hd__clkbuf_4 _13964_ (.A(_04898_),
    .X(_04990_));
 sky130_fd_sc_hd__nand2_1 _13965_ (.A(\samples_imag[7][6] ),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__o21ai_1 _13966_ (.A1(_04929_),
    .A2(_04989_),
    .B1(_04991_),
    .Y(_00416_));
 sky130_fd_sc_hd__buf_4 _13967_ (.A(_04170_),
    .X(_04992_));
 sky130_fd_sc_hd__nor2_2 _13968_ (.A(_04949_),
    .B(_04173_),
    .Y(_04993_));
 sky130_fd_sc_hd__a21oi_1 _13969_ (.A1(\samples_imag[7][7] ),
    .A2(_04984_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_1 _13970_ (.A(_04899_),
    .B(_04177_),
    .Y(_04995_));
 sky130_fd_sc_hd__o21ai_1 _13971_ (.A1(_04915_),
    .A2(_04994_),
    .B1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__a21oi_1 _13972_ (.A1(_04992_),
    .A2(_04996_),
    .B1(_04181_),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _13973_ (.A(\samples_imag[7][7] ),
    .B(_04990_),
    .Y(_04998_));
 sky130_fd_sc_hd__o21ai_1 _13974_ (.A1(_04929_),
    .A2(_04997_),
    .B1(_04998_),
    .Y(_00417_));
 sky130_fd_sc_hd__buf_2 _13975_ (.A(_04897_),
    .X(_04999_));
 sky130_fd_sc_hd__nor2_2 _13976_ (.A(_04949_),
    .B(_04186_),
    .Y(_05000_));
 sky130_fd_sc_hd__a21oi_1 _13977_ (.A1(\samples_imag[7][8] ),
    .A2(_04984_),
    .B1(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__nand2_1 _13978_ (.A(_04899_),
    .B(_04190_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21ai_1 _13979_ (.A1(_04915_),
    .A2(_05001_),
    .B1(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__a21oi_1 _13980_ (.A1(_04992_),
    .A2(_05003_),
    .B1(_04194_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_1 _13981_ (.A(\samples_imag[7][8] ),
    .B(_04990_),
    .Y(_05005_));
 sky130_fd_sc_hd__o21ai_1 _13982_ (.A1(_04999_),
    .A2(_05004_),
    .B1(_05005_),
    .Y(_00418_));
 sky130_fd_sc_hd__nor2_2 _13983_ (.A(_04949_),
    .B(_04198_),
    .Y(_05006_));
 sky130_fd_sc_hd__a21oi_1 _13984_ (.A1(\samples_imag[7][9] ),
    .A2(_04984_),
    .B1(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _13985_ (.A(_04899_),
    .B(_04202_),
    .Y(_05008_));
 sky130_fd_sc_hd__o21ai_1 _13986_ (.A1(_04915_),
    .A2(_05007_),
    .B1(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__a21oi_1 _13987_ (.A1(_04992_),
    .A2(_05009_),
    .B1(_04206_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand2_1 _13988_ (.A(\samples_imag[7][9] ),
    .B(_04990_),
    .Y(_05011_));
 sky130_fd_sc_hd__o21ai_1 _13989_ (.A1(_04999_),
    .A2(_05010_),
    .B1(_05011_),
    .Y(_00419_));
 sky130_fd_sc_hd__xnor2_4 _13990_ (.A(_05882_),
    .B(_07736_),
    .Y(_05012_));
 sky130_fd_sc_hd__clkbuf_2 _13991_ (.A(_07728_),
    .X(_05013_));
 sky130_fd_sc_hd__inv_1 _13992_ (.A(_07742_),
    .Y(_05014_));
 sky130_fd_sc_hd__clkbuf_2 _13993_ (.A(_07747_),
    .X(_05015_));
 sky130_fd_sc_hd__inv_1 _13994_ (.A(_07752_),
    .Y(_05016_));
 sky130_fd_sc_hd__buf_2 _13995_ (.A(_07757_),
    .X(_05017_));
 sky130_fd_sc_hd__inv_1 _13996_ (.A(_07762_),
    .Y(_05018_));
 sky130_fd_sc_hd__clkbuf_2 _13997_ (.A(_07767_),
    .X(_05019_));
 sky130_fd_sc_hd__inv_1 _13998_ (.A(_07772_),
    .Y(_05020_));
 sky130_fd_sc_hd__clkbuf_2 _13999_ (.A(_07777_),
    .X(_05021_));
 sky130_fd_sc_hd__clkbuf_2 _14000_ (.A(_07782_),
    .X(_05022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__xor2_4 clone52 (.A(_05012_),
    .B(_05038_),
    .X(net52));
 sky130_fd_sc_hd__a21o_1 _14003_ (.A1(_05888_),
    .A2(_07796_),
    .B1(_07795_),
    .X(_05025_));
 sky130_fd_sc_hd__a21o_1 _14004_ (.A1(_05025_),
    .A2(_07792_),
    .B1(_07791_),
    .X(_05026_));
 sky130_fd_sc_hd__a21o_1 _14005_ (.A1(_05026_),
    .A2(_07787_),
    .B1(_07786_),
    .X(_05027_));
 sky130_fd_sc_hd__a21o_1 _14006_ (.A1(_05027_),
    .A2(_05022_),
    .B1(_07781_),
    .X(_05028_));
 sky130_fd_sc_hd__a21oi_2 _14007_ (.A1(_05028_),
    .A2(_05021_),
    .B1(_07776_),
    .Y(_05029_));
 sky130_fd_sc_hd__o21bai_2 _14008_ (.A1(_05029_),
    .A2(_05020_),
    .B1_N(_07771_),
    .Y(_05030_));
 sky130_fd_sc_hd__a21oi_2 _14009_ (.A1(_05030_),
    .A2(_05019_),
    .B1(_07766_),
    .Y(_05031_));
 sky130_fd_sc_hd__o21bai_1 _14010_ (.A1(_05031_),
    .A2(_05018_),
    .B1_N(_07761_),
    .Y(_05032_));
 sky130_fd_sc_hd__a21oi_1 _14011_ (.A1(_05017_),
    .A2(_05032_),
    .B1(_07756_),
    .Y(_05033_));
 sky130_fd_sc_hd__o21bai_1 _14012_ (.A1(_05016_),
    .A2(_05033_),
    .B1_N(_07751_),
    .Y(_05034_));
 sky130_fd_sc_hd__a21oi_1 _14013_ (.A1(_05015_),
    .A2(_05034_),
    .B1(_07746_),
    .Y(_05035_));
 sky130_fd_sc_hd__o21bai_1 _14014_ (.A1(_05014_),
    .A2(_05035_),
    .B1_N(_07741_),
    .Y(_05036_));
 sky130_fd_sc_hd__a21o_1 _14015_ (.A1(_05036_),
    .A2(_05013_),
    .B1(_07727_),
    .X(_05037_));
 sky130_fd_sc_hd__a21oi_4 _14016_ (.A1(_07723_),
    .A2(_05037_),
    .B1(_07722_),
    .Y(_05038_));
 sky130_fd_sc_hd__xor2_4 _14017_ (.A(_05012_),
    .B(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__nand3_4 _14018_ (.A(\temp_real[0] ),
    .B(_07739_),
    .C(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_8 _14019_ (.A(_05040_),
    .B(_07733_),
    .Y(_05041_));
 sky130_fd_sc_hd__inv_2 _14020_ (.A(_07796_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21oi_4 _14021_ (.A1(_07731_),
    .A2(_05042_),
    .B1(_07797_),
    .Y(_05043_));
 sky130_fd_sc_hd__nor2_4 _14022_ (.A(_05043_),
    .B(_07792_),
    .Y(_05044_));
 sky130_fd_sc_hd__nor2_4 _14023_ (.A(_05044_),
    .B(_07793_),
    .Y(_05045_));
 sky130_fd_sc_hd__nor2_2 _14024_ (.A(_07787_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__nor2_2 _14025_ (.A(_05046_),
    .B(_07788_),
    .Y(_05047_));
 sky130_fd_sc_hd__nor2_1 _14026_ (.A(_05047_),
    .B(_05022_),
    .Y(_05048_));
 sky130_fd_sc_hd__nor2_2 _14027_ (.A(_05048_),
    .B(_07783_),
    .Y(_05049_));
 sky130_fd_sc_hd__o21bai_1 _14028_ (.A1(_05049_),
    .A2(_05021_),
    .B1_N(_07778_),
    .Y(_05050_));
 sky130_fd_sc_hd__a21oi_2 _14029_ (.A1(_05020_),
    .A2(_05050_),
    .B1(_07773_),
    .Y(_05051_));
 sky130_fd_sc_hd__o21bai_1 _14030_ (.A1(_05051_),
    .A2(_05019_),
    .B1_N(_07768_),
    .Y(_05052_));
 sky130_fd_sc_hd__a21oi_2 _14031_ (.A1(_05052_),
    .A2(_05018_),
    .B1(_07763_),
    .Y(_05053_));
 sky130_fd_sc_hd__o21bai_1 _14032_ (.A1(_05053_),
    .A2(_05017_),
    .B1_N(_07758_),
    .Y(_05054_));
 sky130_fd_sc_hd__a21oi_2 _14033_ (.A1(_05016_),
    .A2(_05054_),
    .B1(_07753_),
    .Y(_05055_));
 sky130_fd_sc_hd__o21bai_1 _14034_ (.A1(_05055_),
    .A2(_05015_),
    .B1_N(_07748_),
    .Y(_05056_));
 sky130_fd_sc_hd__a21oi_2 _14035_ (.A1(_05014_),
    .A2(_05056_),
    .B1(_07743_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_1 _14036_ (.A(_05057_),
    .B(_05013_),
    .Y(_05058_));
 sky130_fd_sc_hd__nor2_1 _14037_ (.A(_05058_),
    .B(_07729_),
    .Y(_05059_));
 sky130_fd_sc_hd__nor2_1 _14038_ (.A(_07723_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nor2_1 _14039_ (.A(_05060_),
    .B(_07724_),
    .Y(_05061_));
 sky130_fd_sc_hd__xnor2_2 _14040_ (.A(_05061_),
    .B(_05012_),
    .Y(_05062_));
 sky130_fd_sc_hd__nor2_1 _14041_ (.A(_07792_),
    .B(_05885_),
    .Y(_05063_));
 sky130_fd_sc_hd__nor2_1 _14042_ (.A(_07793_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _14043_ (.A(_07787_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nor2_2 _14044_ (.A(_05065_),
    .B(_07788_),
    .Y(_05066_));
 sky130_fd_sc_hd__nor2_2 _14045_ (.A(_05022_),
    .B(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_1 _14046_ (.A(_07783_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__nor2_1 _14047_ (.A(_05068_),
    .B(_05021_),
    .Y(_05069_));
 sky130_fd_sc_hd__nor2_2 _14048_ (.A(_05069_),
    .B(_07778_),
    .Y(_05070_));
 sky130_fd_sc_hd__nor2_1 _14049_ (.A(_07772_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nor2_1 _14050_ (.A(_07773_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__nor2_1 _14051_ (.A(_05072_),
    .B(_05019_),
    .Y(_05073_));
 sky130_fd_sc_hd__nor2_2 _14052_ (.A(_05073_),
    .B(_07768_),
    .Y(_05074_));
 sky130_fd_sc_hd__nor2_2 _14053_ (.A(_05074_),
    .B(_07762_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _14054_ (.A(_07763_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nor2_1 _14055_ (.A(_05017_),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__nor2_2 _14056_ (.A(_05077_),
    .B(_07758_),
    .Y(_05078_));
 sky130_fd_sc_hd__nor2_1 _14057_ (.A(_07752_),
    .B(_05078_),
    .Y(_05079_));
 sky130_fd_sc_hd__nor2_1 _14058_ (.A(_05079_),
    .B(_07753_),
    .Y(_05080_));
 sky130_fd_sc_hd__nor2_1 _14059_ (.A(_05080_),
    .B(_05015_),
    .Y(_05081_));
 sky130_fd_sc_hd__nor2_1 _14060_ (.A(_05081_),
    .B(_07748_),
    .Y(_05082_));
 sky130_fd_sc_hd__nor2_1 _14061_ (.A(_07742_),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__nor2_1 _14062_ (.A(_05083_),
    .B(_07743_),
    .Y(_05084_));
 sky130_fd_sc_hd__nor2_1 _14063_ (.A(_05084_),
    .B(_05013_),
    .Y(_05085_));
 sky130_fd_sc_hd__nor2_2 _14064_ (.A(_07729_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__xnor2_2 _14065_ (.A(_05086_),
    .B(_07723_),
    .Y(_05087_));
 sky130_fd_sc_hd__xnor2_1 _14066_ (.A(_05013_),
    .B(net564),
    .Y(_05088_));
 sky130_fd_sc_hd__xnor2_2 _14067_ (.A(net581),
    .B(_07742_),
    .Y(_05089_));
 sky130_fd_sc_hd__xor2_2 _14068_ (.A(_05017_),
    .B(_05053_),
    .X(_05090_));
 sky130_fd_sc_hd__xor2_2 _14069_ (.A(_05015_),
    .B(_05055_),
    .X(_05091_));
 sky130_fd_sc_hd__xnor2_2 _14070_ (.A(_05016_),
    .B(net599),
    .Y(_05092_));
 sky130_fd_sc_hd__xnor2_1 _14071_ (.A(_07772_),
    .B(net592),
    .Y(_05093_));
 sky130_fd_sc_hd__xnor2_1 _14072_ (.A(_05021_),
    .B(_05049_),
    .Y(_05094_));
 sky130_fd_sc_hd__xnor2_1 _14073_ (.A(_07787_),
    .B(net513),
    .Y(_05095_));
 sky130_fd_sc_hd__xor2_2 _14074_ (.A(net617),
    .B(net578),
    .X(_05096_));
 sky130_fd_sc_hd__xor2_2 _14075_ (.A(_05022_),
    .B(_05066_),
    .X(_05097_));
 sky130_fd_sc_hd__nor4b_1 _14076_ (.A(_07733_),
    .B(_05096_),
    .C(_05097_),
    .D_N(_05886_),
    .Y(_05098_));
 sky130_fd_sc_hd__nand4_1 _14077_ (.A(_05093_),
    .B(_05094_),
    .C(_05095_),
    .D(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_4 _14078_ (.A(_05018_),
    .B(net597),
    .Y(_05100_));
 sky130_fd_sc_hd__xor2_1 _14079_ (.A(_05019_),
    .B(_05051_),
    .X(_05101_));
 sky130_fd_sc_hd__or4_4 _14080_ (.A(_05092_),
    .B(_05099_),
    .C(_05100_),
    .D(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__nor3_4 _14081_ (.A(_05090_),
    .B(_05091_),
    .C(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _14082_ (.A(net53),
    .B(_07738_),
    .Y(_05104_));
 sky130_fd_sc_hd__a41oi_4 _14083_ (.A1(_05103_),
    .A2(_05088_),
    .A3(_05089_),
    .A4(_05087_),
    .B1(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2b_4 _14084_ (.A_N(_05062_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__and2_4 _14085_ (.A(_05106_),
    .B(_07733_),
    .X(_05107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__a22o_1 _14087_ (.A1(\samples_real[0][0] ),
    .A2(_03176_),
    .B1(_03995_),
    .B2(_05107_),
    .X(_05109_));
 sky130_fd_sc_hd__nand2_1 _14088_ (.A(_03449_),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__o31ai_1 _14089_ (.A1(_03894_),
    .A2(_03893_),
    .A3(_05041_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2b_1 _14090_ (.A_N(_03141_),
    .B(net74),
    .Y(_05112_));
 sky130_fd_sc_hd__buf_4 _14091_ (.A(_05112_),
    .X(_05113_));
 sky130_fd_sc_hd__nor2_1 _14092_ (.A(_03893_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__a221o_1 _14093_ (.A1(\samples_real[0][0] ),
    .A2(_03893_),
    .B1(_05111_),
    .B2(_03999_),
    .C1(_05114_),
    .X(_00420_));
 sky130_fd_sc_hd__buf_12 _14094_ (.A(_05040_),
    .X(_05115_));
 sky130_fd_sc_hd__a21o_1 _14095_ (.A1(net612),
    .A2(_05889_),
    .B1(_07791_),
    .X(_05116_));
 sky130_fd_sc_hd__a21o_1 _14096_ (.A1(_07787_),
    .A2(_05116_),
    .B1(_07786_),
    .X(_05117_));
 sky130_fd_sc_hd__a21o_1 _14097_ (.A1(_05022_),
    .A2(_05117_),
    .B1(_07781_),
    .X(_05118_));
 sky130_fd_sc_hd__a21oi_1 _14098_ (.A1(_05021_),
    .A2(_05118_),
    .B1(_07776_),
    .Y(_05119_));
 sky130_fd_sc_hd__o21bai_1 _14099_ (.A1(_05020_),
    .A2(_05119_),
    .B1_N(_07771_),
    .Y(_05120_));
 sky130_fd_sc_hd__a21oi_1 _14100_ (.A1(_05019_),
    .A2(_05120_),
    .B1(_07766_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21bai_1 _14101_ (.A1(_05018_),
    .A2(_05121_),
    .B1_N(_07761_),
    .Y(_05122_));
 sky130_fd_sc_hd__a21oi_2 _14102_ (.A1(_05017_),
    .A2(_05122_),
    .B1(_07756_),
    .Y(_05123_));
 sky130_fd_sc_hd__xnor2_2 _14103_ (.A(_07752_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_8 _14104_ (.A(net568),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__buf_12 _14105_ (.A(_05106_),
    .X(_05126_));
 sky130_fd_sc_hd__nand2_8 _14106_ (.A(net577),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _14107_ (.A(\samples_real[0][10] ),
    .B(_04089_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_2 _14108_ (.A1(_03715_),
    .A2(_05127_),
    .B1(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _14109_ (.A(_03466_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_2 _14110_ (.A1(_04108_),
    .A2(_05125_),
    .B1(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__nor2b_1 _14111_ (.A(_04055_),
    .B_N(net75),
    .Y(_05132_));
 sky130_fd_sc_hd__buf_4 _14112_ (.A(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__a21oi_2 _14113_ (.A1(_04992_),
    .A2(_05131_),
    .B1(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _14114_ (.A(\samples_real[0][10] ),
    .B(_04168_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21ai_2 _14115_ (.A1(_04184_),
    .A2(_05134_),
    .B1(_05135_),
    .Y(_00421_));
 sky130_fd_sc_hd__buf_2 _14116_ (.A(_03309_),
    .X(_05136_));
 sky130_fd_sc_hd__xor2_1 _14117_ (.A(_05015_),
    .B(_05034_),
    .X(_05137_));
 sky130_fd_sc_hd__nand2_8 _14118_ (.A(net568),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_8 _14119_ (.A(_05091_),
    .B(_05126_),
    .Y(_05139_));
 sky130_fd_sc_hd__nand2_1 _14120_ (.A(\samples_real[0][11] ),
    .B(_04089_),
    .Y(_05140_));
 sky130_fd_sc_hd__o21ai_2 _14121_ (.A1(_03715_),
    .A2(_05139_),
    .B1(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _14122_ (.A(_03466_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_2 _14123_ (.A1(_05136_),
    .A2(_05138_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2b_1 _14124_ (.A(_04055_),
    .B_N(net76),
    .Y(_05144_));
 sky130_fd_sc_hd__clkbuf_4 _14125_ (.A(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a21oi_2 _14126_ (.A1(_05143_),
    .A2(_04992_),
    .B1(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_1 _14127_ (.A(\samples_real[0][11] ),
    .B(_04168_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_1 _14128_ (.A1(_04184_),
    .A2(_05146_),
    .B1(_05147_),
    .Y(_00422_));
 sky130_fd_sc_hd__o21bai_1 _14129_ (.A1(_05016_),
    .A2(_05123_),
    .B1_N(_07751_),
    .Y(_05148_));
 sky130_fd_sc_hd__a21oi_1 _14130_ (.A1(_05015_),
    .A2(_05148_),
    .B1(_07746_),
    .Y(_05149_));
 sky130_fd_sc_hd__xnor2_1 _14131_ (.A(_07742_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_8 _14132_ (.A(_05115_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2b_4 _14133_ (.A_N(_05089_),
    .B(net64),
    .Y(_05152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__nand2_1 _14135_ (.A(\samples_real[0][12] ),
    .B(_04089_),
    .Y(_05154_));
 sky130_fd_sc_hd__o21ai_2 _14136_ (.A1(_03715_),
    .A2(_05152_),
    .B1(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _14137_ (.A(_03466_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_1 _14138_ (.A1(_05136_),
    .A2(_05151_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nor2b_1 _14139_ (.A(_04055_),
    .B_N(net78),
    .Y(_05158_));
 sky130_fd_sc_hd__clkbuf_4 _14140_ (.A(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a21oi_1 _14141_ (.A1(_04992_),
    .A2(_05157_),
    .B1(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_1 _14142_ (.A(\samples_real[0][12] ),
    .B(_04168_),
    .Y(_05161_));
 sky130_fd_sc_hd__o21ai_1 _14143_ (.A1(_04184_),
    .A2(_05160_),
    .B1(_05161_),
    .Y(_00423_));
 sky130_fd_sc_hd__xor2_1 _14144_ (.A(_05013_),
    .B(_05036_),
    .X(_05162_));
 sky130_fd_sc_hd__nand2_8 _14145_ (.A(_05115_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2b_4 _14146_ (.A_N(_05088_),
    .B(net64),
    .Y(_05164_));
 sky130_fd_sc_hd__buf_6 clone56 (.A(_03149_),
    .X(net56));
 sky130_fd_sc_hd__nand2_1 _14148_ (.A(\samples_real[0][13] ),
    .B(_04089_),
    .Y(_05166_));
 sky130_fd_sc_hd__o21ai_2 _14149_ (.A1(_03715_),
    .A2(_05164_),
    .B1(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_1 _14150_ (.A(_03466_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ai_1 _14151_ (.A1(_05136_),
    .A2(_05163_),
    .B1(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__nor2b_1 _14152_ (.A(_04055_),
    .B_N(net79),
    .Y(_05170_));
 sky130_fd_sc_hd__clkbuf_4 _14153_ (.A(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__a21oi_1 _14154_ (.A1(_04992_),
    .A2(_05169_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _14155_ (.A(\samples_real[0][13] ),
    .B(_04168_),
    .Y(_05173_));
 sky130_fd_sc_hd__o21ai_1 _14156_ (.A1(_04184_),
    .A2(_05172_),
    .B1(_05173_),
    .Y(_00424_));
 sky130_fd_sc_hd__o21bai_1 _14157_ (.A1(_05014_),
    .A2(_05149_),
    .B1_N(_07741_),
    .Y(_05174_));
 sky130_fd_sc_hd__a21oi_1 _14158_ (.A1(_05013_),
    .A2(_05174_),
    .B1(_07727_),
    .Y(_05175_));
 sky130_fd_sc_hd__xnor2_1 _14159_ (.A(_07723_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__nand2_4 _14160_ (.A(_05040_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2b_4 _14161_ (.A_N(_05087_),
    .B(_05106_),
    .Y(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net601));
 sky130_fd_sc_hd__nand2_1 _14163_ (.A(\samples_real[0][14] ),
    .B(_04089_),
    .Y(_05180_));
 sky130_fd_sc_hd__o21ai_2 _14164_ (.A1(_03715_),
    .A2(_05178_),
    .B1(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _14165_ (.A(_03466_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_1 _14166_ (.A1(_05136_),
    .A2(_05177_),
    .B1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__nor2b_1 _14167_ (.A(_04055_),
    .B_N(net80),
    .Y(_05184_));
 sky130_fd_sc_hd__buf_4 _14168_ (.A(_05184_),
    .X(_05185_));
 sky130_fd_sc_hd__a21oi_1 _14169_ (.A1(_04992_),
    .A2(_05183_),
    .B1(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _14170_ (.A(\samples_real[0][14] ),
    .B(_04168_),
    .Y(_05187_));
 sky130_fd_sc_hd__o21ai_1 _14171_ (.A1(_04184_),
    .A2(_05186_),
    .B1(_05187_),
    .Y(_00425_));
 sky130_fd_sc_hd__nor2_4 _14172_ (.A(_05062_),
    .B(net567),
    .Y(_05188_));
 sky130_fd_sc_hd__nand2_1 _14173_ (.A(\samples_real[0][15] ),
    .B(_04091_),
    .Y(_05189_));
 sky130_fd_sc_hd__o211ai_1 _14174_ (.A1(_04089_),
    .A2(_05188_),
    .B1(_05189_),
    .C1(_03309_),
    .Y(_05190_));
 sky130_fd_sc_hd__o21ai_0 _14175_ (.A1(_03894_),
    .A2(net566),
    .B1(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__nor2_4 _14176_ (.A(_03142_),
    .B(net81),
    .Y(_05192_));
 sky130_fd_sc_hd__a211oi_1 _14177_ (.A1(_04029_),
    .A2(_05191_),
    .B1(_05192_),
    .C1(_04087_),
    .Y(_05193_));
 sky130_fd_sc_hd__a21o_1 _14178_ (.A1(\samples_real[0][15] ),
    .A2(_04087_),
    .B1(_05193_),
    .X(_00426_));
 sky130_fd_sc_hd__nand2b_4 _14179_ (.A_N(_05886_),
    .B(_05106_),
    .Y(_05194_));
 sky130_fd_sc_hd__buf_6 rebuffer244 (.A(_05219_),
    .X(net619));
 sky130_fd_sc_hd__nor2_4 _14181_ (.A(_04089_),
    .B(_05194_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_2 _14182_ (.A1(\samples_real[0][1] ),
    .A2(_03715_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a31oi_4 _14183_ (.A1(net53),
    .A2(net565),
    .A3(_07739_),
    .B1(_05890_),
    .Y(_05198_));
 sky130_fd_sc_hd__nor2_1 _14184_ (.A(_03894_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__a21oi_1 _14185_ (.A1(_05197_),
    .A2(_04108_),
    .B1(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__nor2b_2 _14186_ (.A(_04023_),
    .B_N(net82),
    .Y(_05201_));
 sky130_fd_sc_hd__buf_4 _14187_ (.A(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__a21oi_1 _14188_ (.A1(_05200_),
    .A2(_04992_),
    .B1(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_1 _14189_ (.A(\samples_real[0][1] ),
    .B(_04168_),
    .Y(_05204_));
 sky130_fd_sc_hd__o21ai_1 _14190_ (.A1(_05203_),
    .A2(_04184_),
    .B1(_05204_),
    .Y(_00427_));
 sky130_fd_sc_hd__xor2_1 _14191_ (.A(net612),
    .B(_05889_),
    .X(_05205_));
 sky130_fd_sc_hd__nand2_8 _14192_ (.A(_05115_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_8 _14193_ (.A(_05096_),
    .B(_05126_),
    .Y(_05207_));
 sky130_fd_sc_hd__nand2_1 _14194_ (.A(\samples_real[0][2] ),
    .B(_04091_),
    .Y(_05208_));
 sky130_fd_sc_hd__o21ai_2 _14195_ (.A1(_03715_),
    .A2(_05207_),
    .B1(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand2_1 _14196_ (.A(_03466_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__o21ai_2 _14197_ (.A1(_05136_),
    .A2(_05206_),
    .B1(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nor2b_1 _14198_ (.A(_03141_),
    .B_N(net83),
    .Y(_05212_));
 sky130_fd_sc_hd__buf_4 _14199_ (.A(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__a21oi_2 _14200_ (.A1(_05211_),
    .A2(_04992_),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(\samples_real[0][2] ),
    .B(_04003_),
    .Y(_05215_));
 sky130_fd_sc_hd__o21ai_2 _14202_ (.A1(_04184_),
    .A2(_05214_),
    .B1(_05215_),
    .Y(_00428_));
 sky130_fd_sc_hd__clkbuf_4 _14203_ (.A(_04236_),
    .X(_05216_));
 sky130_fd_sc_hd__xor2_1 _14204_ (.A(_07787_),
    .B(_05026_),
    .X(_05217_));
 sky130_fd_sc_hd__nand2_8 _14205_ (.A(net568),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand2b_4 _14206_ (.A_N(_05095_),
    .B(net64),
    .Y(_05219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__nand2_1 _14208_ (.A(\samples_real[0][3] ),
    .B(_04091_),
    .Y(_05221_));
 sky130_fd_sc_hd__o21ai_2 _14209_ (.A1(_03177_),
    .A2(_05219_),
    .B1(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__nand2_1 _14210_ (.A(_03466_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_2 _14211_ (.A1(_05218_),
    .A2(_05136_),
    .B1(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__nor2b_1 _14212_ (.A(_03141_),
    .B_N(net84),
    .Y(_05225_));
 sky130_fd_sc_hd__buf_4 _14213_ (.A(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__a21oi_2 _14214_ (.A1(_05224_),
    .A2(_05216_),
    .B1(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2_1 _14215_ (.A(\samples_real[0][3] ),
    .B(_04003_),
    .Y(_05228_));
 sky130_fd_sc_hd__o21ai_2 _14216_ (.A1(_04184_),
    .A2(_05227_),
    .B1(_05228_),
    .Y(_00429_));
 sky130_fd_sc_hd__xor2_1 _14217_ (.A(_05022_),
    .B(_05117_),
    .X(_05229_));
 sky130_fd_sc_hd__nand2_4 _14218_ (.A(_05115_),
    .B(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand2_8 _14219_ (.A(_05097_),
    .B(_05126_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _14220_ (.A(\samples_real[0][4] ),
    .B(_04091_),
    .Y(_05232_));
 sky130_fd_sc_hd__o21ai_2 _14221_ (.A1(_05231_),
    .A2(_03177_),
    .B1(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hd__nand2_1 _14222_ (.A(_03449_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_2 _14223_ (.A1(_05136_),
    .A2(_05230_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__nor2b_1 _14224_ (.A(_03141_),
    .B_N(net85),
    .Y(_05236_));
 sky130_fd_sc_hd__buf_4 _14225_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__a21oi_2 _14226_ (.A1(_05216_),
    .A2(_05235_),
    .B1(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__nand2_1 _14227_ (.A(\samples_real[0][4] ),
    .B(_04003_),
    .Y(_05239_));
 sky130_fd_sc_hd__o21ai_1 _14228_ (.A1(_05238_),
    .A2(_04087_),
    .B1(_05239_),
    .Y(_00430_));
 sky130_fd_sc_hd__xor2_1 _14229_ (.A(_05021_),
    .B(_05028_),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_8 _14230_ (.A(net568),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__nand2b_4 _14231_ (.A_N(_05094_),
    .B(_05106_),
    .Y(_05242_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(data_valid_in),
    .X(net649));
 sky130_fd_sc_hd__nand2_1 _14233_ (.A(\samples_real[0][5] ),
    .B(_04091_),
    .Y(_05244_));
 sky130_fd_sc_hd__o21ai_1 _14234_ (.A1(_03177_),
    .A2(_05242_),
    .B1(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_1 _14235_ (.A(_03449_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__o21ai_2 _14236_ (.A1(_05136_),
    .A2(_05241_),
    .B1(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__nor2b_1 _14237_ (.A(_03141_),
    .B_N(net86),
    .Y(_05248_));
 sky130_fd_sc_hd__buf_4 _14238_ (.A(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__a21oi_2 _14239_ (.A1(_05247_),
    .A2(_05216_),
    .B1(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_1 _14240_ (.A(\samples_real[0][5] ),
    .B(_04003_),
    .Y(_05251_));
 sky130_fd_sc_hd__o21ai_1 _14241_ (.A1(_05250_),
    .A2(_04087_),
    .B1(_05251_),
    .Y(_00431_));
 sky130_fd_sc_hd__xnor2_2 _14242_ (.A(_07772_),
    .B(_05119_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_8 _14243_ (.A(_05040_),
    .B(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2b_4 _14244_ (.A_N(_05093_),
    .B(_05106_),
    .Y(_05254_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(rst_n),
    .X(net648));
 sky130_fd_sc_hd__nand2_1 _14246_ (.A(\samples_real[0][6] ),
    .B(_04091_),
    .Y(_05256_));
 sky130_fd_sc_hd__o21ai_2 _14247_ (.A1(_05254_),
    .A2(_03177_),
    .B1(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__nand2_1 _14248_ (.A(_03449_),
    .B(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__o21ai_1 _14249_ (.A1(_05136_),
    .A2(_05253_),
    .B1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__nor2b_1 _14250_ (.A(_03141_),
    .B_N(net87),
    .Y(_05260_));
 sky130_fd_sc_hd__clkbuf_8 _14251_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__a21oi_1 _14252_ (.A1(_05259_),
    .A2(_05216_),
    .B1(_05261_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_1 _14253_ (.A(\samples_real[0][6] ),
    .B(_04003_),
    .Y(_05263_));
 sky130_fd_sc_hd__o21ai_1 _14254_ (.A1(_04087_),
    .A2(_05262_),
    .B1(_05263_),
    .Y(_00432_));
 sky130_fd_sc_hd__xor2_2 _14255_ (.A(_05019_),
    .B(_05030_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_8 _14256_ (.A(net568),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_8 _14257_ (.A(_05101_),
    .B(net64),
    .Y(_05266_));
 sky130_fd_sc_hd__nand2_1 _14258_ (.A(\samples_real[0][7] ),
    .B(_04091_),
    .Y(_05267_));
 sky130_fd_sc_hd__o21ai_2 _14259_ (.A1(_03177_),
    .A2(_05266_),
    .B1(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _14260_ (.A(_03449_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_1 _14261_ (.A1(_05136_),
    .A2(_05265_),
    .B1(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__nor2b_1 _14262_ (.A(_03141_),
    .B_N(net88),
    .Y(_05271_));
 sky130_fd_sc_hd__buf_4 _14263_ (.A(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__a21oi_1 _14264_ (.A1(_05270_),
    .A2(_05216_),
    .B1(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__nand2_1 _14265_ (.A(\samples_real[0][7] ),
    .B(_04003_),
    .Y(_05274_));
 sky130_fd_sc_hd__o21ai_1 _14266_ (.A1(_04087_),
    .A2(_05273_),
    .B1(_05274_),
    .Y(_00433_));
 sky130_fd_sc_hd__xnor2_1 _14267_ (.A(_07762_),
    .B(_05121_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_8 _14268_ (.A(_05115_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_8 _14269_ (.A(_05100_),
    .B(net64),
    .Y(_05277_));
 sky130_fd_sc_hd__nand2_1 _14270_ (.A(\samples_real[0][8] ),
    .B(_04091_),
    .Y(_05278_));
 sky130_fd_sc_hd__o21ai_2 _14271_ (.A1(_03177_),
    .A2(_05277_),
    .B1(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _14272_ (.A(_03449_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21ai_1 _14273_ (.A1(_03466_),
    .A2(_05276_),
    .B1(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nor2b_1 _14274_ (.A(_03141_),
    .B_N(net89),
    .Y(_05282_));
 sky130_fd_sc_hd__buf_4 _14275_ (.A(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__a21oi_1 _14276_ (.A1(_05216_),
    .A2(_05281_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2_1 _14277_ (.A(\samples_real[0][8] ),
    .B(_04003_),
    .Y(_05285_));
 sky130_fd_sc_hd__o21ai_1 _14278_ (.A1(_04087_),
    .A2(_05284_),
    .B1(_05285_),
    .Y(_00434_));
 sky130_fd_sc_hd__xor2_2 _14279_ (.A(_05017_),
    .B(net573),
    .X(_05286_));
 sky130_fd_sc_hd__nand2_4 _14280_ (.A(_05040_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__nand2_8 _14281_ (.A(_05090_),
    .B(_05126_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(\samples_real[0][9] ),
    .B(_04091_),
    .Y(_05289_));
 sky130_fd_sc_hd__o21ai_2 _14283_ (.A1(_03177_),
    .A2(_05288_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_1 _14284_ (.A(_03449_),
    .B(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__o21ai_1 _14285_ (.A1(_03466_),
    .A2(_05287_),
    .B1(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nor2b_1 _14286_ (.A(\state[1] ),
    .B_N(net90),
    .Y(_05293_));
 sky130_fd_sc_hd__buf_4 _14287_ (.A(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a21oi_1 _14288_ (.A1(_05216_),
    .A2(_05292_),
    .B1(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_1 _14289_ (.A(\samples_real[0][9] ),
    .B(_04003_),
    .Y(_05296_));
 sky130_fd_sc_hd__o21ai_1 _14290_ (.A1(_04087_),
    .A2(_05295_),
    .B1(_05296_),
    .Y(_00435_));
 sky130_fd_sc_hd__a22oi_2 _14291_ (.A1(\samples_real[1][0] ),
    .A2(_04217_),
    .B1(_05107_),
    .B2(_04219_),
    .Y(_05297_));
 sky130_fd_sc_hd__nor2_1 _14292_ (.A(_05297_),
    .B(_04214_),
    .Y(_05298_));
 sky130_fd_sc_hd__nor3_1 _14293_ (.A(_04222_),
    .B(_04212_),
    .C(_05041_),
    .Y(_05299_));
 sky130_fd_sc_hd__o21ai_1 _14294_ (.A1(_05299_),
    .A2(_05298_),
    .B1(_04004_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _14295_ (.A(\samples_real[1][0] ),
    .B(_04227_),
    .Y(_05301_));
 sky130_fd_sc_hd__o211ai_1 _14296_ (.A1(_04246_),
    .A2(_05113_),
    .B1(_05301_),
    .C1(_05300_),
    .Y(_00436_));
 sky130_fd_sc_hd__nor2_4 _14297_ (.A(_04265_),
    .B(_05127_),
    .Y(_05302_));
 sky130_fd_sc_hd__a211oi_2 _14298_ (.A1(\samples_real[1][10] ),
    .A2(_04239_),
    .B1(_04243_),
    .C1(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__a21oi_1 _14299_ (.A1(_04214_),
    .A2(_05125_),
    .B1(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21oi_1 _14300_ (.A1(_05216_),
    .A2(_05304_),
    .B1(_05133_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _14301_ (.A(\samples_real[1][10] ),
    .B(_04286_),
    .Y(_05306_));
 sky130_fd_sc_hd__o21ai_1 _14302_ (.A1(_04318_),
    .A2(_05305_),
    .B1(_05306_),
    .Y(_00437_));
 sky130_fd_sc_hd__clkbuf_4 _14303_ (.A(_04216_),
    .X(_05307_));
 sky130_fd_sc_hd__nor2_4 _14304_ (.A(_04265_),
    .B(_05139_),
    .Y(_05308_));
 sky130_fd_sc_hd__a211oi_2 _14305_ (.A1(\samples_real[1][11] ),
    .A2(_05307_),
    .B1(_04243_),
    .C1(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _14306_ (.A1(_04214_),
    .A2(_05138_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__a21oi_2 _14307_ (.A1(_05310_),
    .A2(_05216_),
    .B1(_05145_),
    .Y(_05311_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(\samples_real[1][11] ),
    .B(_04286_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_1 _14309_ (.A1(_04318_),
    .A2(_05311_),
    .B1(_05312_),
    .Y(_00438_));
 sky130_fd_sc_hd__nor2_2 _14310_ (.A(_04265_),
    .B(_05152_),
    .Y(_05313_));
 sky130_fd_sc_hd__a211oi_2 _14311_ (.A1(\samples_real[1][12] ),
    .A2(_05307_),
    .B1(_04243_),
    .C1(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__a21oi_2 _14312_ (.A1(_04214_),
    .A2(_05151_),
    .B1(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__a21oi_2 _14313_ (.A1(_05315_),
    .A2(_05216_),
    .B1(_05159_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _14314_ (.A(\samples_real[1][12] ),
    .B(_04286_),
    .Y(_05317_));
 sky130_fd_sc_hd__o21ai_2 _14315_ (.A1(_04318_),
    .A2(_05316_),
    .B1(_05317_),
    .Y(_00439_));
 sky130_fd_sc_hd__clkbuf_4 _14316_ (.A(_04236_),
    .X(_05318_));
 sky130_fd_sc_hd__nor2_4 _14317_ (.A(_04265_),
    .B(_05164_),
    .Y(_05319_));
 sky130_fd_sc_hd__a211oi_2 _14318_ (.A1(\samples_real[1][13] ),
    .A2(_05307_),
    .B1(_04243_),
    .C1(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__a21oi_2 _14319_ (.A1(_04214_),
    .A2(_05163_),
    .B1(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__a21oi_2 _14320_ (.A1(_05321_),
    .A2(_05318_),
    .B1(_05171_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2_1 _14321_ (.A(\samples_real[1][13] ),
    .B(_04286_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21ai_1 _14322_ (.A1(_04318_),
    .A2(_05322_),
    .B1(_05323_),
    .Y(_00440_));
 sky130_fd_sc_hd__buf_4 _14323_ (.A(_03142_),
    .X(_05324_));
 sky130_fd_sc_hd__nand2_1 _14324_ (.A(_04214_),
    .B(_05177_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _14325_ (.A(\samples_real[1][14] ),
    .B(_04217_),
    .Y(_05326_));
 sky130_fd_sc_hd__o211ai_1 _14326_ (.A1(_04217_),
    .A2(_05178_),
    .B1(_05326_),
    .C1(_04222_),
    .Y(_05327_));
 sky130_fd_sc_hd__a311oi_1 _14327_ (.A1(_05324_),
    .A2(_05325_),
    .A3(_05327_),
    .B1(_04212_),
    .C1(_05185_),
    .Y(_05328_));
 sky130_fd_sc_hd__a21oi_1 _14328_ (.A1(_03692_),
    .A2(_04213_),
    .B1(_05328_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _14329_ (.A(\samples_real[1][15] ),
    .B(_04216_),
    .Y(_05329_));
 sky130_fd_sc_hd__o211ai_1 _14330_ (.A1(_04265_),
    .A2(_05188_),
    .B1(_05329_),
    .C1(_04222_),
    .Y(_05330_));
 sky130_fd_sc_hd__o21ai_0 _14331_ (.A1(_04222_),
    .A2(net52),
    .B1(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a211oi_2 _14332_ (.A1(_04029_),
    .A2(_05331_),
    .B1(_05192_),
    .C1(_04212_),
    .Y(_05332_));
 sky130_fd_sc_hd__a21o_1 _14333_ (.A1(\samples_real[1][15] ),
    .A2(_04246_),
    .B1(_05332_),
    .X(_00442_));
 sky130_fd_sc_hd__nor2_2 _14334_ (.A(_04265_),
    .B(_05194_),
    .Y(_05333_));
 sky130_fd_sc_hd__a21oi_1 _14335_ (.A1(\samples_real[1][1] ),
    .A2(_04239_),
    .B1(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__nand2_1 _14336_ (.A(_04238_),
    .B(_05198_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21ai_2 _14337_ (.A1(_04231_),
    .A2(_05334_),
    .B1(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__a21oi_2 _14338_ (.A1(_05336_),
    .A2(_05318_),
    .B1(_05202_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _14339_ (.A(\samples_real[1][1] ),
    .B(_04225_),
    .Y(_05338_));
 sky130_fd_sc_hd__o21ai_1 _14340_ (.A1(_04318_),
    .A2(_05337_),
    .B1(_05338_),
    .Y(_00443_));
 sky130_fd_sc_hd__nor2_4 _14341_ (.A(_04265_),
    .B(_05207_),
    .Y(_05339_));
 sky130_fd_sc_hd__a211oi_1 _14342_ (.A1(\samples_real[1][2] ),
    .A2(_05307_),
    .B1(_04243_),
    .C1(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21oi_1 _14343_ (.A1(_04214_),
    .A2(_05206_),
    .B1(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__a21oi_1 _14344_ (.A1(_05318_),
    .A2(_05341_),
    .B1(_05213_),
    .Y(_05342_));
 sky130_fd_sc_hd__nand2_1 _14345_ (.A(\samples_real[1][2] ),
    .B(_04225_),
    .Y(_05343_));
 sky130_fd_sc_hd__o21ai_1 _14346_ (.A1(_04318_),
    .A2(_05342_),
    .B1(_05343_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2_1 _14347_ (.A(_04240_),
    .B(_05219_),
    .Y(_05344_));
 sky130_fd_sc_hd__a211oi_1 _14348_ (.A1(\samples_real[1][3] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__a21oi_1 _14349_ (.A1(_04214_),
    .A2(_05218_),
    .B1(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__a21oi_1 _14350_ (.A1(_05346_),
    .A2(_05318_),
    .B1(_05226_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand2_1 _14351_ (.A(\samples_real[1][3] ),
    .B(_04225_),
    .Y(_05348_));
 sky130_fd_sc_hd__o21ai_1 _14352_ (.A1(_04318_),
    .A2(_05347_),
    .B1(_05348_),
    .Y(_00445_));
 sky130_fd_sc_hd__nor2_2 _14353_ (.A(_04240_),
    .B(_05231_),
    .Y(_05349_));
 sky130_fd_sc_hd__a211oi_1 _14354_ (.A1(\samples_real[1][4] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__a21oi_1 _14355_ (.A1(_04214_),
    .A2(_05230_),
    .B1(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a21oi_1 _14356_ (.A1(_05351_),
    .A2(_05318_),
    .B1(_05237_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _14357_ (.A(\samples_real[1][4] ),
    .B(_04225_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21ai_1 _14358_ (.A1(_05352_),
    .A2(_04318_),
    .B1(_05353_),
    .Y(_00446_));
 sky130_fd_sc_hd__nor2_1 _14359_ (.A(_04240_),
    .B(_05242_),
    .Y(_05354_));
 sky130_fd_sc_hd__a211oi_1 _14360_ (.A1(\samples_real[1][5] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__a21oi_1 _14361_ (.A1(_04228_),
    .A2(_05241_),
    .B1(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__a21oi_1 _14362_ (.A1(_05318_),
    .A2(_05356_),
    .B1(_05249_),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_1 _14363_ (.A(\samples_real[1][5] ),
    .B(_04225_),
    .Y(_05358_));
 sky130_fd_sc_hd__o21ai_0 _14364_ (.A1(_04318_),
    .A2(_05357_),
    .B1(_05358_),
    .Y(_00447_));
 sky130_fd_sc_hd__nor2_1 _14365_ (.A(_04240_),
    .B(_05254_),
    .Y(_05359_));
 sky130_fd_sc_hd__a211oi_1 _14366_ (.A1(\samples_real[1][6] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__a21oi_1 _14367_ (.A1(_04228_),
    .A2(_05253_),
    .B1(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__a21oi_1 _14368_ (.A1(_05318_),
    .A2(_05361_),
    .B1(_05261_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _14369_ (.A(\samples_real[1][6] ),
    .B(_04225_),
    .Y(_05363_));
 sky130_fd_sc_hd__o21ai_1 _14370_ (.A1(_04246_),
    .A2(_05362_),
    .B1(_05363_),
    .Y(_00448_));
 sky130_fd_sc_hd__nor2_2 _14371_ (.A(_04240_),
    .B(_05266_),
    .Y(_05364_));
 sky130_fd_sc_hd__a211oi_1 _14372_ (.A1(\samples_real[1][7] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__a21oi_1 _14373_ (.A1(_04228_),
    .A2(_05265_),
    .B1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a21oi_1 _14374_ (.A1(_05318_),
    .A2(_05366_),
    .B1(_05272_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _14375_ (.A(\samples_real[1][7] ),
    .B(_04225_),
    .Y(_05368_));
 sky130_fd_sc_hd__o21ai_1 _14376_ (.A1(_04246_),
    .A2(_05367_),
    .B1(_05368_),
    .Y(_00449_));
 sky130_fd_sc_hd__nor2_4 _14377_ (.A(_04240_),
    .B(_05277_),
    .Y(_05369_));
 sky130_fd_sc_hd__a211oi_2 _14378_ (.A1(\samples_real[1][8] ),
    .A2(_05307_),
    .B1(_03469_),
    .C1(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__a21oi_1 _14379_ (.A1(_04228_),
    .A2(_05276_),
    .B1(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__a21oi_1 _14380_ (.A1(_05371_),
    .A2(_05318_),
    .B1(_05283_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _14381_ (.A(\samples_real[1][8] ),
    .B(_04225_),
    .Y(_05373_));
 sky130_fd_sc_hd__o21ai_1 _14382_ (.A1(_05372_),
    .A2(_04246_),
    .B1(_05373_),
    .Y(_00450_));
 sky130_fd_sc_hd__nor2_4 _14383_ (.A(_04240_),
    .B(_05288_),
    .Y(_05374_));
 sky130_fd_sc_hd__a211oi_2 _14384_ (.A1(\samples_real[1][9] ),
    .A2(_04218_),
    .B1(_03469_),
    .C1(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__a21oi_1 _14385_ (.A1(_04228_),
    .A2(_05287_),
    .B1(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a21oi_1 _14386_ (.A1(_05376_),
    .A2(_05318_),
    .B1(_05294_),
    .Y(_05377_));
 sky130_fd_sc_hd__nand2_1 _14387_ (.A(\samples_real[1][9] ),
    .B(_04225_),
    .Y(_05378_));
 sky130_fd_sc_hd__o21ai_1 _14388_ (.A1(_04246_),
    .A2(_05377_),
    .B1(_05378_),
    .Y(_00451_));
 sky130_fd_sc_hd__a22oi_2 _14389_ (.A1(\samples_real[2][0] ),
    .A2(_04332_),
    .B1(_04334_),
    .B2(_05107_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor2_1 _14390_ (.A(_04329_),
    .B(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__nor3_1 _14391_ (.A(_04337_),
    .B(_04327_),
    .C(_05041_),
    .Y(_05381_));
 sky130_fd_sc_hd__o21ai_1 _14392_ (.A1(_05381_),
    .A2(_05380_),
    .B1(_04004_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand2_1 _14393_ (.A(\samples_real[2][0] ),
    .B(_04342_),
    .Y(_05383_));
 sky130_fd_sc_hd__o211ai_2 _14394_ (.A1(_04377_),
    .A2(_05113_),
    .B1(_05383_),
    .C1(_05382_),
    .Y(_00452_));
 sky130_fd_sc_hd__buf_2 _14395_ (.A(_04236_),
    .X(_05384_));
 sky130_fd_sc_hd__buf_2 _14396_ (.A(_04331_),
    .X(_05385_));
 sky130_fd_sc_hd__nor2_4 _14397_ (.A(_05385_),
    .B(_05127_),
    .Y(_05386_));
 sky130_fd_sc_hd__a211oi_2 _14398_ (.A1(\samples_real[2][10] ),
    .A2(_04429_),
    .B1(_04424_),
    .C1(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__a21oi_2 _14399_ (.A1(_04329_),
    .A2(_05125_),
    .B1(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__a21oi_2 _14400_ (.A1(_05388_),
    .A2(_05384_),
    .B1(_05133_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _14401_ (.A(\samples_real[2][10] ),
    .B(_04388_),
    .Y(_05390_));
 sky130_fd_sc_hd__o21ai_1 _14402_ (.A1(_04409_),
    .A2(_05389_),
    .B1(_05390_),
    .Y(_00453_));
 sky130_fd_sc_hd__nor2_4 _14403_ (.A(_05139_),
    .B(_05385_),
    .Y(_05391_));
 sky130_fd_sc_hd__a211oi_2 _14404_ (.A1(\samples_real[2][11] ),
    .A2(_04429_),
    .B1(_04424_),
    .C1(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__a21oi_2 _14405_ (.A1(_04329_),
    .A2(_05138_),
    .B1(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__a21oi_2 _14406_ (.A1(_05384_),
    .A2(_05393_),
    .B1(_05145_),
    .Y(_05394_));
 sky130_fd_sc_hd__nand2_1 _14407_ (.A(\samples_real[2][11] ),
    .B(_04388_),
    .Y(_05395_));
 sky130_fd_sc_hd__o21ai_1 _14408_ (.A1(_05394_),
    .A2(_04409_),
    .B1(_05395_),
    .Y(_00454_));
 sky130_fd_sc_hd__nor2_4 _14409_ (.A(_05152_),
    .B(_05385_),
    .Y(_05396_));
 sky130_fd_sc_hd__a211oi_2 _14410_ (.A1(\samples_real[2][12] ),
    .A2(_04429_),
    .B1(_04424_),
    .C1(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a21oi_2 _14411_ (.A1(_04329_),
    .A2(_05151_),
    .B1(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__a21oi_2 _14412_ (.A1(_05398_),
    .A2(_05384_),
    .B1(_05159_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2_1 _14413_ (.A(\samples_real[2][12] ),
    .B(_04340_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_1 _14414_ (.A1(_05399_),
    .A2(_04409_),
    .B1(_05400_),
    .Y(_00455_));
 sky130_fd_sc_hd__nor2_4 _14415_ (.A(_05385_),
    .B(_05164_),
    .Y(_05401_));
 sky130_fd_sc_hd__a211oi_2 _14416_ (.A1(\samples_real[2][13] ),
    .A2(_04429_),
    .B1(_04424_),
    .C1(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__a21oi_2 _14417_ (.A1(_04329_),
    .A2(_05163_),
    .B1(_05402_),
    .Y(_05403_));
 sky130_fd_sc_hd__a21oi_2 _14418_ (.A1(_05384_),
    .A2(_05403_),
    .B1(_05171_),
    .Y(_05404_));
 sky130_fd_sc_hd__nand2_1 _14419_ (.A(\samples_real[2][13] ),
    .B(_04340_),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ai_1 _14420_ (.A1(_04409_),
    .A2(_05404_),
    .B1(_05405_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_04329_),
    .B(_05177_),
    .Y(_05406_));
 sky130_fd_sc_hd__nand2_1 _14422_ (.A(\samples_real[2][14] ),
    .B(_04332_),
    .Y(_05407_));
 sky130_fd_sc_hd__o211ai_1 _14423_ (.A1(_04332_),
    .A2(_05178_),
    .B1(_05407_),
    .C1(_04337_),
    .Y(_05408_));
 sky130_fd_sc_hd__a311oi_1 _14424_ (.A1(_03999_),
    .A2(_05406_),
    .A3(_05408_),
    .B1(_04377_),
    .C1(_05185_),
    .Y(_05409_));
 sky130_fd_sc_hd__a21oi_1 _14425_ (.A1(_03527_),
    .A2(_04328_),
    .B1(_05409_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _14426_ (.A(\samples_real[2][15] ),
    .B(_04331_),
    .Y(_05410_));
 sky130_fd_sc_hd__o211ai_1 _14427_ (.A1(_04378_),
    .A2(_05188_),
    .B1(_05410_),
    .C1(_04337_),
    .Y(_05411_));
 sky130_fd_sc_hd__o21ai_0 _14428_ (.A1(_04337_),
    .A2(net52),
    .B1(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__a211oi_2 _14429_ (.A1(_04029_),
    .A2(_05412_),
    .B1(_05192_),
    .C1(_04327_),
    .Y(_05413_));
 sky130_fd_sc_hd__a21o_1 _14430_ (.A1(\samples_real[2][15] ),
    .A2(_04377_),
    .B1(_05413_),
    .X(_00458_));
 sky130_fd_sc_hd__nor2_4 _14431_ (.A(_05194_),
    .B(_04378_),
    .Y(_05414_));
 sky130_fd_sc_hd__a21oi_2 _14432_ (.A1(\samples_real[2][1] ),
    .A2(_04429_),
    .B1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _14433_ (.A(_04424_),
    .B(_05198_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21ai_2 _14434_ (.A1(_04346_),
    .A2(_05415_),
    .B1(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__a21oi_2 _14435_ (.A1(_05384_),
    .A2(_05417_),
    .B1(_05202_),
    .Y(_05418_));
 sky130_fd_sc_hd__nand2_1 _14436_ (.A(\samples_real[2][1] ),
    .B(_04340_),
    .Y(_05419_));
 sky130_fd_sc_hd__o21ai_1 _14437_ (.A1(_05418_),
    .A2(_04409_),
    .B1(_05419_),
    .Y(_00459_));
 sky130_fd_sc_hd__nor2_4 _14438_ (.A(_05207_),
    .B(_05385_),
    .Y(_05420_));
 sky130_fd_sc_hd__a211oi_2 _14439_ (.A1(\samples_real[2][2] ),
    .A2(_04429_),
    .B1(_04424_),
    .C1(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21oi_2 _14440_ (.A1(_04329_),
    .A2(_05206_),
    .B1(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__a21oi_2 _14441_ (.A1(_05422_),
    .A2(_05384_),
    .B1(_05213_),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_1 _14442_ (.A(\samples_real[2][2] ),
    .B(_04340_),
    .Y(_05424_));
 sky130_fd_sc_hd__o21ai_1 _14443_ (.A1(_05423_),
    .A2(_04409_),
    .B1(_05424_),
    .Y(_00460_));
 sky130_fd_sc_hd__nor2_2 _14444_ (.A(_05385_),
    .B(_05219_),
    .Y(_05425_));
 sky130_fd_sc_hd__a211oi_2 _14445_ (.A1(\samples_real[2][3] ),
    .A2(_04429_),
    .B1(_05425_),
    .C1(_03437_),
    .Y(_05426_));
 sky130_fd_sc_hd__a21oi_2 _14446_ (.A1(_04343_),
    .A2(_05218_),
    .B1(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__a21oi_2 _14447_ (.A1(_05384_),
    .A2(_05427_),
    .B1(_05226_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_1 _14448_ (.A(\samples_real[2][3] ),
    .B(_04340_),
    .Y(_05429_));
 sky130_fd_sc_hd__o21ai_1 _14449_ (.A1(_04377_),
    .A2(_05428_),
    .B1(_05429_),
    .Y(_00461_));
 sky130_fd_sc_hd__nor2_4 _14450_ (.A(_05231_),
    .B(_05385_),
    .Y(_05430_));
 sky130_fd_sc_hd__a211oi_2 _14451_ (.A1(\samples_real[2][4] ),
    .A2(_04429_),
    .B1(_03437_),
    .C1(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21oi_2 _14452_ (.A1(_04343_),
    .A2(_05230_),
    .B1(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21oi_2 _14453_ (.A1(_05432_),
    .A2(_05384_),
    .B1(_05237_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand2_1 _14454_ (.A(\samples_real[2][4] ),
    .B(_04340_),
    .Y(_05434_));
 sky130_fd_sc_hd__o21ai_1 _14455_ (.A1(_05433_),
    .A2(_04377_),
    .B1(_05434_),
    .Y(_00462_));
 sky130_fd_sc_hd__nor2_1 _14456_ (.A(_05385_),
    .B(_05242_),
    .Y(_05435_));
 sky130_fd_sc_hd__a211oi_1 _14457_ (.A1(\samples_real[2][5] ),
    .A2(_04333_),
    .B1(_03437_),
    .C1(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__a21oi_1 _14458_ (.A1(_04343_),
    .A2(_05241_),
    .B1(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__a21oi_1 _14459_ (.A1(_05384_),
    .A2(_05437_),
    .B1(_05249_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _14460_ (.A(\samples_real[2][5] ),
    .B(_04340_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_0 _14461_ (.A1(_04377_),
    .A2(_05438_),
    .B1(_05439_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _14462_ (.A(_04329_),
    .B(_05253_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _14463_ (.A(\samples_real[2][6] ),
    .B(_04332_),
    .Y(_05441_));
 sky130_fd_sc_hd__o211ai_1 _14464_ (.A1(_04332_),
    .A2(_05254_),
    .B1(_05441_),
    .C1(_04337_),
    .Y(_05442_));
 sky130_fd_sc_hd__a311oi_1 _14465_ (.A1(_03999_),
    .A2(_05440_),
    .A3(_05442_),
    .B1(_04327_),
    .C1(_05261_),
    .Y(_05443_));
 sky130_fd_sc_hd__a21oi_1 _14466_ (.A1(_03734_),
    .A2(_04328_),
    .B1(_05443_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_4 _14467_ (.A(_05385_),
    .B(_05266_),
    .Y(_05444_));
 sky130_fd_sc_hd__a211oi_2 _14468_ (.A1(\samples_real[2][7] ),
    .A2(_04333_),
    .B1(_03437_),
    .C1(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__a21oi_1 _14469_ (.A1(_04343_),
    .A2(_05265_),
    .B1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__a21oi_1 _14470_ (.A1(_05384_),
    .A2(_05446_),
    .B1(_05272_),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(\samples_real[2][7] ),
    .B(_04340_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_1 _14472_ (.A1(_04377_),
    .A2(_05447_),
    .B1(_05448_),
    .Y(_00465_));
 sky130_fd_sc_hd__buf_6 _14473_ (.A(_04236_),
    .X(_05449_));
 sky130_fd_sc_hd__nor2_2 _14474_ (.A(_05277_),
    .B(_05385_),
    .Y(_05450_));
 sky130_fd_sc_hd__a211oi_2 _14475_ (.A1(\samples_real[2][8] ),
    .A2(_04333_),
    .B1(_03437_),
    .C1(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__a21oi_1 _14476_ (.A1(_04343_),
    .A2(_05276_),
    .B1(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__a21oi_1 _14477_ (.A1(_05449_),
    .A2(_05452_),
    .B1(_05283_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _14478_ (.A(\samples_real[2][8] ),
    .B(_04340_),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_1 _14479_ (.A1(_04377_),
    .A2(_05453_),
    .B1(_05454_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _14480_ (.A(_04329_),
    .B(_05287_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_1 _14481_ (.A(\samples_real[2][9] ),
    .B(_04332_),
    .Y(_05456_));
 sky130_fd_sc_hd__o211ai_2 _14482_ (.A1(_05288_),
    .A2(_04332_),
    .B1(_05456_),
    .C1(_04337_),
    .Y(_05457_));
 sky130_fd_sc_hd__a311oi_1 _14483_ (.A1(_03999_),
    .A2(_05455_),
    .A3(_05457_),
    .B1(_04327_),
    .C1(_05294_),
    .Y(_05458_));
 sky130_fd_sc_hd__a21oi_1 _14484_ (.A1(_03380_),
    .A2(_04328_),
    .B1(_05458_),
    .Y(_00467_));
 sky130_fd_sc_hd__a22oi_2 _14485_ (.A1(\samples_real[3][0] ),
    .A2(_04447_),
    .B1(_05107_),
    .B2(_04448_),
    .Y(_05459_));
 sky130_fd_sc_hd__o22ai_1 _14486_ (.A1(_04451_),
    .A2(_05041_),
    .B1(_04455_),
    .B2(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__nor2_1 _14487_ (.A(_04444_),
    .B(_05113_),
    .Y(_05461_));
 sky130_fd_sc_hd__a221o_1 _14488_ (.A1(\samples_real[3][0] ),
    .A2(_04444_),
    .B1(_05460_),
    .B2(_03999_),
    .C1(_05461_),
    .X(_00468_));
 sky130_fd_sc_hd__clkbuf_4 _14489_ (.A(_04236_),
    .X(_05462_));
 sky130_fd_sc_hd__buf_2 _14490_ (.A(_03439_),
    .X(_05463_));
 sky130_fd_sc_hd__nand2_1 _14491_ (.A(_05463_),
    .B(_05125_),
    .Y(_05464_));
 sky130_fd_sc_hd__buf_2 _14492_ (.A(_04446_),
    .X(_05465_));
 sky130_fd_sc_hd__buf_2 _14493_ (.A(_04446_),
    .X(_05466_));
 sky130_fd_sc_hd__nand2_1 _14494_ (.A(\samples_real[3][10] ),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__buf_2 _14495_ (.A(_04450_),
    .X(_05468_));
 sky130_fd_sc_hd__o211ai_2 _14496_ (.A1(_05465_),
    .A2(_05127_),
    .B1(_05467_),
    .C1(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__a31oi_1 _14497_ (.A1(_05464_),
    .A2(_05469_),
    .A3(_05462_),
    .B1(_05133_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _14498_ (.A(\samples_real[3][10] ),
    .B(_04534_),
    .Y(_05471_));
 sky130_fd_sc_hd__o21ai_1 _14499_ (.A1(_05470_),
    .A2(_04542_),
    .B1(_05471_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _14500_ (.A(_05463_),
    .B(_05138_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _14501_ (.A(\samples_real[3][11] ),
    .B(_05466_),
    .Y(_05473_));
 sky130_fd_sc_hd__o211ai_2 _14502_ (.A1(_05465_),
    .A2(_05139_),
    .B1(_05473_),
    .C1(_05468_),
    .Y(_05474_));
 sky130_fd_sc_hd__a31oi_2 _14503_ (.A1(_05472_),
    .A2(_05474_),
    .A3(_05462_),
    .B1(_05145_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_1 _14504_ (.A(\samples_real[3][11] ),
    .B(_04534_),
    .Y(_05476_));
 sky130_fd_sc_hd__o21ai_1 _14505_ (.A1(_04542_),
    .A2(_05475_),
    .B1(_05476_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _14506_ (.A(_05463_),
    .B(_05151_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_1 _14507_ (.A(\samples_real[3][12] ),
    .B(_05466_),
    .Y(_05478_));
 sky130_fd_sc_hd__o211ai_2 _14508_ (.A1(_05465_),
    .A2(_05152_),
    .B1(_05478_),
    .C1(_05468_),
    .Y(_05479_));
 sky130_fd_sc_hd__a31oi_2 _14509_ (.A1(_05477_),
    .A2(_05479_),
    .A3(_05462_),
    .B1(_05159_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _14510_ (.A(\samples_real[3][12] ),
    .B(_04534_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_1 _14511_ (.A1(_04542_),
    .A2(_05480_),
    .B1(_05481_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _14512_ (.A(_05463_),
    .B(_05163_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(\samples_real[3][13] ),
    .B(_05466_),
    .Y(_05483_));
 sky130_fd_sc_hd__o211ai_2 _14514_ (.A1(_05465_),
    .A2(_05164_),
    .B1(_05483_),
    .C1(_05468_),
    .Y(_05484_));
 sky130_fd_sc_hd__a31oi_2 _14515_ (.A1(_05482_),
    .A2(_05484_),
    .A3(_05462_),
    .B1(_05171_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _14516_ (.A(\samples_real[3][13] ),
    .B(_04534_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_1 _14517_ (.A1(_04542_),
    .A2(_05485_),
    .B1(_05486_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _14518_ (.A(_05463_),
    .B(_05177_),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _14519_ (.A(\samples_real[3][14] ),
    .B(_05466_),
    .Y(_05488_));
 sky130_fd_sc_hd__o211ai_2 _14520_ (.A1(_05465_),
    .A2(_05178_),
    .B1(_05488_),
    .C1(_05468_),
    .Y(_05489_));
 sky130_fd_sc_hd__a31oi_2 _14521_ (.A1(_05462_),
    .A2(_05487_),
    .A3(_05489_),
    .B1(_05185_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _14522_ (.A(\samples_real[3][14] ),
    .B(_04534_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_1 _14523_ (.A1(_04542_),
    .A2(_05490_),
    .B1(_05491_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _14524_ (.A(\samples_real[3][15] ),
    .B(_04446_),
    .Y(_05492_));
 sky130_fd_sc_hd__o211ai_1 _14525_ (.A1(_04494_),
    .A2(_05188_),
    .B1(_05492_),
    .C1(_04450_),
    .Y(_05493_));
 sky130_fd_sc_hd__o21ai_0 _14526_ (.A1(_04450_),
    .A2(net52),
    .B1(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__a211oi_1 _14527_ (.A1(_04029_),
    .A2(_05494_),
    .B1(_05192_),
    .C1(_04493_),
    .Y(_05495_));
 sky130_fd_sc_hd__a21o_1 _14528_ (.A1(\samples_real[3][15] ),
    .A2(_04493_),
    .B1(_05495_),
    .X(_00474_));
 sky130_fd_sc_hd__nor2_2 _14529_ (.A(_04494_),
    .B(_05194_),
    .Y(_05496_));
 sky130_fd_sc_hd__a21oi_1 _14530_ (.A1(\samples_real[3][1] ),
    .A2(_04447_),
    .B1(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_1 _14531_ (.A(_03439_),
    .B(_05198_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_1 _14532_ (.A1(_04459_),
    .A2(_05497_),
    .B1(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__a21oi_1 _14533_ (.A1(_05449_),
    .A2(_05499_),
    .B1(_05202_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _14534_ (.A(\samples_real[3][1] ),
    .B(_04534_),
    .Y(_05501_));
 sky130_fd_sc_hd__o21ai_1 _14535_ (.A1(_04542_),
    .A2(_05500_),
    .B1(_05501_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _14536_ (.A(_05463_),
    .B(_05206_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(\samples_real[3][2] ),
    .B(_05466_),
    .Y(_05503_));
 sky130_fd_sc_hd__o211ai_2 _14538_ (.A1(_05465_),
    .A2(_05207_),
    .B1(_05503_),
    .C1(_05468_),
    .Y(_05504_));
 sky130_fd_sc_hd__a31oi_1 _14539_ (.A1(_05462_),
    .A2(_05504_),
    .A3(_05502_),
    .B1(_05213_),
    .Y(_05505_));
 sky130_fd_sc_hd__nand2_1 _14540_ (.A(\samples_real[3][2] ),
    .B(_04454_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_1 _14541_ (.A1(_04542_),
    .A2(_05505_),
    .B1(_05506_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _14542_ (.A(_05463_),
    .B(_05218_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _14543_ (.A(\samples_real[3][3] ),
    .B(_05466_),
    .Y(_05508_));
 sky130_fd_sc_hd__o211ai_2 _14544_ (.A1(_05465_),
    .A2(_05219_),
    .B1(_05508_),
    .C1(_05468_),
    .Y(_05509_));
 sky130_fd_sc_hd__a31oi_1 _14545_ (.A1(_05507_),
    .A2(_05509_),
    .A3(_05462_),
    .B1(_05226_),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _14546_ (.A(\samples_real[3][3] ),
    .B(_04454_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_1 _14547_ (.A1(_05510_),
    .A2(_04542_),
    .B1(_05511_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _14548_ (.A(_05463_),
    .B(_05230_),
    .Y(_05512_));
 sky130_fd_sc_hd__nand2_1 _14549_ (.A(\samples_real[3][4] ),
    .B(_04456_),
    .Y(_05513_));
 sky130_fd_sc_hd__o211ai_2 _14550_ (.A1(_05465_),
    .A2(_05231_),
    .B1(_05513_),
    .C1(_05468_),
    .Y(_05514_));
 sky130_fd_sc_hd__a31oi_1 _14551_ (.A1(_05462_),
    .A2(_05514_),
    .A3(_05512_),
    .B1(_05237_),
    .Y(_05515_));
 sky130_fd_sc_hd__nand2_1 _14552_ (.A(\samples_real[3][4] ),
    .B(_04454_),
    .Y(_05516_));
 sky130_fd_sc_hd__o21ai_1 _14553_ (.A1(_04493_),
    .A2(_05515_),
    .B1(_05516_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _14554_ (.A(_05463_),
    .B(_05241_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _14555_ (.A(\samples_real[3][5] ),
    .B(_04456_),
    .Y(_05518_));
 sky130_fd_sc_hd__o211ai_1 _14556_ (.A1(_05465_),
    .A2(_05242_),
    .B1(_05518_),
    .C1(_05468_),
    .Y(_05519_));
 sky130_fd_sc_hd__a31oi_1 _14557_ (.A1(_05462_),
    .A2(_05517_),
    .A3(_05519_),
    .B1(_05249_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_1 _14558_ (.A(\samples_real[3][5] ),
    .B(_04454_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_0 _14559_ (.A1(_04493_),
    .A2(_05520_),
    .B1(_05521_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _14560_ (.A(_05463_),
    .B(_05253_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _14561_ (.A(\samples_real[3][6] ),
    .B(_04456_),
    .Y(_05523_));
 sky130_fd_sc_hd__o211ai_1 _14562_ (.A1(_05465_),
    .A2(_05254_),
    .B1(_05523_),
    .C1(_05468_),
    .Y(_05524_));
 sky130_fd_sc_hd__a31oi_1 _14563_ (.A1(_05462_),
    .A2(_05522_),
    .A3(_05524_),
    .B1(_05261_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _14564_ (.A(\samples_real[3][6] ),
    .B(_04454_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21ai_0 _14565_ (.A1(_04493_),
    .A2(_05525_),
    .B1(_05526_),
    .Y(_00480_));
 sky130_fd_sc_hd__buf_4 _14566_ (.A(_04236_),
    .X(_05527_));
 sky130_fd_sc_hd__nand2_2 _14567_ (.A(_05265_),
    .B(_04455_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _14568_ (.A(\samples_real[3][7] ),
    .B(_04456_),
    .Y(_05529_));
 sky130_fd_sc_hd__o211ai_2 _14569_ (.A1(_05466_),
    .A2(_05266_),
    .B1(_05529_),
    .C1(_04450_),
    .Y(_05530_));
 sky130_fd_sc_hd__a31oi_1 _14570_ (.A1(_05527_),
    .A2(_05528_),
    .A3(_05530_),
    .B1(_05272_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(\samples_real[3][7] ),
    .B(_04454_),
    .Y(_05532_));
 sky130_fd_sc_hd__o21ai_1 _14572_ (.A1(_05531_),
    .A2(_04493_),
    .B1(_05532_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _14573_ (.A(_04455_),
    .B(_05276_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(\samples_real[3][8] ),
    .B(_04456_),
    .Y(_05534_));
 sky130_fd_sc_hd__o211ai_2 _14575_ (.A1(_05277_),
    .A2(_05466_),
    .B1(_05534_),
    .C1(_04450_),
    .Y(_05535_));
 sky130_fd_sc_hd__a31oi_1 _14576_ (.A1(_05527_),
    .A2(_05533_),
    .A3(_05535_),
    .B1(_05283_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand2_1 _14577_ (.A(\samples_real[3][8] ),
    .B(_04454_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_1 _14578_ (.A1(_04493_),
    .A2(_05536_),
    .B1(_05537_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _14579_ (.A(_04455_),
    .B(_05287_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(\samples_real[3][9] ),
    .B(_04456_),
    .Y(_05539_));
 sky130_fd_sc_hd__o211ai_2 _14581_ (.A1(_05466_),
    .A2(_05288_),
    .B1(_05539_),
    .C1(_04450_),
    .Y(_05540_));
 sky130_fd_sc_hd__a31oi_1 _14582_ (.A1(_05527_),
    .A2(_05540_),
    .A3(_05538_),
    .B1(_05294_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _14583_ (.A(\samples_real[3][9] ),
    .B(_04454_),
    .Y(_05542_));
 sky130_fd_sc_hd__o21ai_1 _14584_ (.A1(_04493_),
    .A2(_05541_),
    .B1(_05542_),
    .Y(_00483_));
 sky130_fd_sc_hd__a22oi_1 _14585_ (.A1(\samples_real[4][0] ),
    .A2(_04560_),
    .B1(_04562_),
    .B2(_05107_),
    .Y(_05543_));
 sky130_fd_sc_hd__nor2_1 _14586_ (.A(_04557_),
    .B(_05041_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_1 _14587_ (.A(_04564_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21ai_0 _14588_ (.A1(_04564_),
    .A2(_05543_),
    .B1(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__nor2_1 _14589_ (.A(_04557_),
    .B(_05113_),
    .Y(_05547_));
 sky130_fd_sc_hd__a221o_1 _14590_ (.A1(\samples_real[4][0] ),
    .A2(_04557_),
    .B1(_05546_),
    .B2(_04088_),
    .C1(_05547_),
    .X(_00484_));
 sky130_fd_sc_hd__buf_2 _14591_ (.A(_04556_),
    .X(_05548_));
 sky130_fd_sc_hd__buf_2 _14592_ (.A(_03467_),
    .X(_05549_));
 sky130_fd_sc_hd__nor2_4 _14593_ (.A(_05127_),
    .B(_04655_),
    .Y(_05550_));
 sky130_fd_sc_hd__a211oi_2 _14594_ (.A1(\samples_real[4][10] ),
    .A2(_04588_),
    .B1(_04564_),
    .C1(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__a21oi_2 _14595_ (.A1(_05549_),
    .A2(_05125_),
    .B1(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__a21oi_1 _14596_ (.A1(_05552_),
    .A2(_05449_),
    .B1(_05133_),
    .Y(_05553_));
 sky130_fd_sc_hd__nand2_1 _14597_ (.A(\samples_real[4][10] ),
    .B(_04646_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_1 _14598_ (.A1(_05553_),
    .A2(_05548_),
    .B1(_05554_),
    .Y(_00485_));
 sky130_fd_sc_hd__buf_2 _14599_ (.A(_03272_),
    .X(_05555_));
 sky130_fd_sc_hd__nor2_4 _14600_ (.A(_04655_),
    .B(_05139_),
    .Y(_05556_));
 sky130_fd_sc_hd__a211oi_2 _14601_ (.A1(\samples_real[4][11] ),
    .A2(_04588_),
    .B1(_05555_),
    .C1(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__a21oi_2 _14602_ (.A1(_05549_),
    .A2(_05138_),
    .B1(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a21oi_1 _14603_ (.A1(_05449_),
    .A2(_05558_),
    .B1(_05145_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _14604_ (.A(\samples_real[4][11] ),
    .B(_04646_),
    .Y(_05560_));
 sky130_fd_sc_hd__o21ai_1 _14605_ (.A1(_05559_),
    .A2(_05548_),
    .B1(_05560_),
    .Y(_00486_));
 sky130_fd_sc_hd__nor2_4 _14606_ (.A(_04655_),
    .B(_05152_),
    .Y(_05561_));
 sky130_fd_sc_hd__a211oi_1 _14607_ (.A1(\samples_real[4][12] ),
    .A2(_04588_),
    .B1(_05555_),
    .C1(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__a21oi_1 _14608_ (.A1(_05549_),
    .A2(_05151_),
    .B1(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__a21oi_1 _14609_ (.A1(_05563_),
    .A2(_05449_),
    .B1(_05159_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _14610_ (.A(\samples_real[4][12] ),
    .B(_04646_),
    .Y(_05565_));
 sky130_fd_sc_hd__o21ai_1 _14611_ (.A1(_05548_),
    .A2(_05564_),
    .B1(_05565_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_4 _14612_ (.A(_04655_),
    .B(_05164_),
    .Y(_05566_));
 sky130_fd_sc_hd__a211oi_2 _14613_ (.A1(\samples_real[4][13] ),
    .A2(_04588_),
    .B1(_05555_),
    .C1(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__a21oi_1 _14614_ (.A1(_05549_),
    .A2(_05163_),
    .B1(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__a21oi_1 _14615_ (.A1(_05449_),
    .A2(_05568_),
    .B1(_05171_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(\samples_real[4][13] ),
    .B(_04646_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21ai_1 _14617_ (.A1(_05548_),
    .A2(_05569_),
    .B1(_05570_),
    .Y(_00488_));
 sky130_fd_sc_hd__nor2_2 _14618_ (.A(_04655_),
    .B(_05178_),
    .Y(_05571_));
 sky130_fd_sc_hd__a211oi_1 _14619_ (.A1(\samples_real[4][14] ),
    .A2(_04588_),
    .B1(_05555_),
    .C1(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__a21oi_1 _14620_ (.A1(_05549_),
    .A2(_05177_),
    .B1(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__a21oi_1 _14621_ (.A1(_05573_),
    .A2(_05449_),
    .B1(_05185_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_1 _14622_ (.A(\samples_real[4][14] ),
    .B(_04646_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_1 _14623_ (.A1(_05548_),
    .A2(_05574_),
    .B1(_05575_),
    .Y(_00489_));
 sky130_fd_sc_hd__nor2_1 _14624_ (.A(\samples_real[4][15] ),
    .B(net549),
    .Y(_05576_));
 sky130_fd_sc_hd__a211oi_1 _14625_ (.A1(net551),
    .A2(_05188_),
    .B1(_05576_),
    .C1(_03467_),
    .Y(_05577_));
 sky130_fd_sc_hd__a21oi_1 _14626_ (.A1(_04564_),
    .A2(net52),
    .B1(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__a211oi_1 _14627_ (.A1(_04029_),
    .A2(_05578_),
    .B1(_05192_),
    .C1(_04593_),
    .Y(_05579_));
 sky130_fd_sc_hd__a21o_1 _14628_ (.A1(\samples_real[4][15] ),
    .A2(_04593_),
    .B1(_05579_),
    .X(_00490_));
 sky130_fd_sc_hd__nor2_2 _14629_ (.A(_04655_),
    .B(_05194_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21oi_1 _14630_ (.A1(\samples_real[4][1] ),
    .A2(_04588_),
    .B1(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _14631_ (.A(_04558_),
    .B(_05198_),
    .Y(_05582_));
 sky130_fd_sc_hd__o21ai_1 _14632_ (.A1(_04576_),
    .A2(_05581_),
    .B1(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__a21oi_1 _14633_ (.A1(_05449_),
    .A2(_05583_),
    .B1(_05202_),
    .Y(_05584_));
 sky130_fd_sc_hd__nand2_1 _14634_ (.A(\samples_real[4][1] ),
    .B(_04646_),
    .Y(_05585_));
 sky130_fd_sc_hd__o21ai_1 _14635_ (.A1(_05548_),
    .A2(_05584_),
    .B1(_05585_),
    .Y(_00491_));
 sky130_fd_sc_hd__nor2_4 _14636_ (.A(_04655_),
    .B(_05207_),
    .Y(_05586_));
 sky130_fd_sc_hd__a211oi_2 _14637_ (.A1(\samples_real[4][2] ),
    .A2(_04560_),
    .B1(_05555_),
    .C1(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__a21oi_1 _14638_ (.A1(_05549_),
    .A2(_05206_),
    .B1(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__a21oi_1 _14639_ (.A1(_05449_),
    .A2(_05588_),
    .B1(_05213_),
    .Y(_05589_));
 sky130_fd_sc_hd__nand2_1 _14640_ (.A(\samples_real[4][2] ),
    .B(_04569_),
    .Y(_05590_));
 sky130_fd_sc_hd__o21ai_1 _14641_ (.A1(_05548_),
    .A2(_05589_),
    .B1(_05590_),
    .Y(_00492_));
 sky130_fd_sc_hd__nor2_4 _14642_ (.A(_04655_),
    .B(net619),
    .Y(_05591_));
 sky130_fd_sc_hd__a211oi_2 _14643_ (.A1(\samples_real[4][3] ),
    .A2(_04560_),
    .B1(_05555_),
    .C1(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__a21oi_2 _14644_ (.A1(_05549_),
    .A2(_05218_),
    .B1(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__a21oi_2 _14645_ (.A1(_05593_),
    .A2(_05449_),
    .B1(_05226_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _14646_ (.A(\samples_real[4][3] ),
    .B(_04569_),
    .Y(_05595_));
 sky130_fd_sc_hd__o21ai_1 _14647_ (.A1(_05548_),
    .A2(_05594_),
    .B1(_05595_),
    .Y(_00493_));
 sky130_fd_sc_hd__clkbuf_4 _14648_ (.A(_04236_),
    .X(_05596_));
 sky130_fd_sc_hd__nor2_4 _14649_ (.A(_04561_),
    .B(_05231_),
    .Y(_05597_));
 sky130_fd_sc_hd__a211oi_2 _14650_ (.A1(\samples_real[4][4] ),
    .A2(_04560_),
    .B1(_05555_),
    .C1(_05597_),
    .Y(_05598_));
 sky130_fd_sc_hd__a21oi_1 _14651_ (.A1(_05549_),
    .A2(_05230_),
    .B1(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__a21oi_1 _14652_ (.A1(_05599_),
    .A2(_05596_),
    .B1(_05237_),
    .Y(_05600_));
 sky130_fd_sc_hd__nand2_1 _14653_ (.A(\samples_real[4][4] ),
    .B(_04569_),
    .Y(_05601_));
 sky130_fd_sc_hd__o21ai_1 _14654_ (.A1(_05548_),
    .A2(_05600_),
    .B1(_05601_),
    .Y(_00494_));
 sky130_fd_sc_hd__nor2_1 _14655_ (.A(_04561_),
    .B(_05242_),
    .Y(_05602_));
 sky130_fd_sc_hd__a211oi_1 _14656_ (.A1(\samples_real[4][5] ),
    .A2(_04560_),
    .B1(_05555_),
    .C1(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__a21oi_2 _14657_ (.A1(_05549_),
    .A2(_05241_),
    .B1(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__a21oi_2 _14658_ (.A1(_05604_),
    .A2(_05596_),
    .B1(_05249_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _14659_ (.A(\samples_real[4][5] ),
    .B(_04569_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_1 _14660_ (.A1(_05605_),
    .A2(_05548_),
    .B1(_05606_),
    .Y(_00495_));
 sky130_fd_sc_hd__nor2_4 _14661_ (.A(_04561_),
    .B(_05254_),
    .Y(_05607_));
 sky130_fd_sc_hd__a211oi_2 _14662_ (.A1(\samples_real[4][6] ),
    .A2(_04560_),
    .B1(_05555_),
    .C1(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21oi_1 _14663_ (.A1(_05549_),
    .A2(_05253_),
    .B1(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__a21oi_1 _14664_ (.A1(_05596_),
    .A2(_05609_),
    .B1(_05261_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand2_1 _14665_ (.A(\samples_real[4][6] ),
    .B(_04569_),
    .Y(_05611_));
 sky130_fd_sc_hd__o21ai_1 _14666_ (.A1(_04593_),
    .A2(_05610_),
    .B1(_05611_),
    .Y(_00496_));
 sky130_fd_sc_hd__nor2_2 _14667_ (.A(_04561_),
    .B(_05266_),
    .Y(_05612_));
 sky130_fd_sc_hd__a211oi_1 _14668_ (.A1(\samples_real[4][7] ),
    .A2(_04560_),
    .B1(_05612_),
    .C1(_05555_),
    .Y(_05613_));
 sky130_fd_sc_hd__a21oi_1 _14669_ (.A1(_04571_),
    .A2(_05265_),
    .B1(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__a21oi_1 _14670_ (.A1(_05614_),
    .A2(_05596_),
    .B1(_05272_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(\samples_real[4][7] ),
    .B(_04569_),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_1 _14672_ (.A1(_04593_),
    .A2(_05615_),
    .B1(_05616_),
    .Y(_00497_));
 sky130_fd_sc_hd__nor2_4 _14673_ (.A(_04561_),
    .B(_05277_),
    .Y(_05617_));
 sky130_fd_sc_hd__a211oi_2 _14674_ (.A1(\samples_real[4][8] ),
    .A2(_04560_),
    .B1(_05617_),
    .C1(_03467_),
    .Y(_05618_));
 sky130_fd_sc_hd__a21oi_1 _14675_ (.A1(_04571_),
    .A2(_05276_),
    .B1(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__a21oi_1 _14676_ (.A1(_05619_),
    .A2(_05596_),
    .B1(_05283_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _14677_ (.A(\samples_real[4][8] ),
    .B(_04569_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_1 _14678_ (.A1(_05620_),
    .A2(_04593_),
    .B1(_05621_),
    .Y(_00498_));
 sky130_fd_sc_hd__nor2_4 _14679_ (.A(_05288_),
    .B(_04561_),
    .Y(_05622_));
 sky130_fd_sc_hd__a211oi_2 _14680_ (.A1(\samples_real[4][9] ),
    .A2(_04560_),
    .B1(_03467_),
    .C1(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__a21oi_2 _14681_ (.A1(_04571_),
    .A2(_05287_),
    .B1(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__a21oi_1 _14682_ (.A1(_05624_),
    .A2(_05596_),
    .B1(_05294_),
    .Y(_05625_));
 sky130_fd_sc_hd__nand2_1 _14683_ (.A(\samples_real[4][9] ),
    .B(_04569_),
    .Y(_05626_));
 sky130_fd_sc_hd__o21ai_1 _14684_ (.A1(_05625_),
    .A2(_04593_),
    .B1(_05626_),
    .Y(_00499_));
 sky130_fd_sc_hd__a22oi_1 _14685_ (.A1(\samples_real[5][0] ),
    .A2(_04673_),
    .B1(_04675_),
    .B2(_05107_),
    .Y(_05627_));
 sky130_fd_sc_hd__nor2_1 _14686_ (.A(_04672_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__nor3_1 _14687_ (.A(_04680_),
    .B(_04670_),
    .C(_05041_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_0 _14688_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_04004_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _14689_ (.A(\samples_real[5][0] ),
    .B(_04685_),
    .Y(_05631_));
 sky130_fd_sc_hd__o211ai_1 _14690_ (.A1(_04719_),
    .A2(_05113_),
    .B1(_05630_),
    .C1(_05631_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _14691_ (.A(_04672_),
    .B(_05125_),
    .Y(_05632_));
 sky130_fd_sc_hd__buf_2 _14692_ (.A(_03773_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_4 _14693_ (.A(_03773_),
    .X(_05634_));
 sky130_fd_sc_hd__nand2_1 _14694_ (.A(\samples_real[5][10] ),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__o211ai_2 _14695_ (.A1(_05633_),
    .A2(_05127_),
    .B1(_05635_),
    .C1(_04680_),
    .Y(_05636_));
 sky130_fd_sc_hd__a31oi_1 _14696_ (.A1(_05527_),
    .A2(_05636_),
    .A3(_05632_),
    .B1(_05133_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(\samples_real[5][10] ),
    .B(_04755_),
    .Y(_05638_));
 sky130_fd_sc_hd__o21ai_1 _14698_ (.A1(_04757_),
    .A2(_05637_),
    .B1(_05638_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _14699_ (.A(_04672_),
    .B(_05138_),
    .Y(_05639_));
 sky130_fd_sc_hd__nand2_1 _14700_ (.A(\samples_real[5][11] ),
    .B(_05634_),
    .Y(_05640_));
 sky130_fd_sc_hd__o211ai_2 _14701_ (.A1(_05633_),
    .A2(_05139_),
    .B1(_05640_),
    .C1(_04680_),
    .Y(_05641_));
 sky130_fd_sc_hd__a31oi_1 _14702_ (.A1(_05527_),
    .A2(_05639_),
    .A3(_05641_),
    .B1(_05145_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_1 _14703_ (.A(\samples_real[5][11] ),
    .B(_04755_),
    .Y(_05643_));
 sky130_fd_sc_hd__o21ai_1 _14704_ (.A1(_04757_),
    .A2(_05642_),
    .B1(_05643_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _14705_ (.A(_04672_),
    .B(_05151_),
    .Y(_05644_));
 sky130_fd_sc_hd__nand2_1 _14706_ (.A(\samples_real[5][12] ),
    .B(_05634_),
    .Y(_05645_));
 sky130_fd_sc_hd__o211ai_2 _14707_ (.A1(_05633_),
    .A2(_05152_),
    .B1(_05645_),
    .C1(_04680_),
    .Y(_05646_));
 sky130_fd_sc_hd__a31oi_1 _14708_ (.A1(_05527_),
    .A2(_05646_),
    .A3(_05644_),
    .B1(_05159_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _14709_ (.A(\samples_real[5][12] ),
    .B(_04755_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_1 _14710_ (.A1(_05647_),
    .A2(_04757_),
    .B1(_05648_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _14711_ (.A(_04672_),
    .B(_05163_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_1 _14712_ (.A(\samples_real[5][13] ),
    .B(_05634_),
    .Y(_05650_));
 sky130_fd_sc_hd__o211ai_2 _14713_ (.A1(_05633_),
    .A2(_05164_),
    .B1(_05650_),
    .C1(_04680_),
    .Y(_05651_));
 sky130_fd_sc_hd__a31oi_1 _14714_ (.A1(_05527_),
    .A2(_05651_),
    .A3(_05649_),
    .B1(_05171_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _14715_ (.A(\samples_real[5][13] ),
    .B(_04755_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_1 _14716_ (.A1(_04757_),
    .A2(_05652_),
    .B1(_05653_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _14717_ (.A(_04672_),
    .B(_05177_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _14718_ (.A(\samples_real[5][14] ),
    .B(_05634_),
    .Y(_05655_));
 sky130_fd_sc_hd__o211ai_2 _14719_ (.A1(_05633_),
    .A2(_05178_),
    .B1(_05655_),
    .C1(_04680_),
    .Y(_05656_));
 sky130_fd_sc_hd__a31oi_1 _14720_ (.A1(_05527_),
    .A2(_05654_),
    .A3(_05656_),
    .B1(_05185_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_1 _14721_ (.A(\samples_real[5][14] ),
    .B(_04755_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_1 _14722_ (.A1(_04757_),
    .A2(_05657_),
    .B1(_05658_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _14723_ (.A(\samples_real[5][15] ),
    .B(_03773_),
    .Y(_05659_));
 sky130_fd_sc_hd__o211ai_1 _14724_ (.A1(_04720_),
    .A2(_05188_),
    .B1(_05659_),
    .C1(_04679_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21ai_0 _14725_ (.A1(_04679_),
    .A2(net593),
    .B1(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__a211oi_1 _14726_ (.A1(_04029_),
    .A2(_05661_),
    .B1(_05192_),
    .C1(_04670_),
    .Y(_05662_));
 sky130_fd_sc_hd__a21o_1 _14727_ (.A1(\samples_real[5][15] ),
    .A2(_04670_),
    .B1(_05662_),
    .X(_00506_));
 sky130_fd_sc_hd__nor2_2 _14728_ (.A(_04720_),
    .B(_05194_),
    .Y(_05663_));
 sky130_fd_sc_hd__a21oi_1 _14729_ (.A1(\samples_real[5][1] ),
    .A2(_04674_),
    .B1(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_03346_),
    .B(_05198_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_1 _14731_ (.A1(_05664_),
    .A2(_04689_),
    .B1(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__a21oi_1 _14732_ (.A1(_05666_),
    .A2(_05596_),
    .B1(_05202_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _14733_ (.A(\samples_real[5][1] ),
    .B(_04683_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_1 _14734_ (.A1(_04757_),
    .A2(_05667_),
    .B1(_05668_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _14735_ (.A(_04672_),
    .B(_05206_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_1 _14736_ (.A(\samples_real[5][2] ),
    .B(_05634_),
    .Y(_05670_));
 sky130_fd_sc_hd__o211ai_2 _14737_ (.A1(_05633_),
    .A2(_05207_),
    .B1(_05670_),
    .C1(_04680_),
    .Y(_05671_));
 sky130_fd_sc_hd__a31oi_1 _14738_ (.A1(_05527_),
    .A2(_05671_),
    .A3(_05669_),
    .B1(_05213_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand2_1 _14739_ (.A(\samples_real[5][2] ),
    .B(_04683_),
    .Y(_05673_));
 sky130_fd_sc_hd__o21ai_1 _14740_ (.A1(_04719_),
    .A2(_05672_),
    .B1(_05673_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_2 _14741_ (.A(_04672_),
    .B(_05218_),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _14742_ (.A(\samples_real[5][3] ),
    .B(_05634_),
    .Y(_05675_));
 sky130_fd_sc_hd__o211ai_2 _14743_ (.A1(_05633_),
    .A2(net619),
    .B1(_05675_),
    .C1(_04680_),
    .Y(_05676_));
 sky130_fd_sc_hd__a31oi_1 _14744_ (.A1(_05527_),
    .A2(_05674_),
    .A3(_05676_),
    .B1(_05226_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _14745_ (.A(\samples_real[5][3] ),
    .B(_04683_),
    .Y(_05678_));
 sky130_fd_sc_hd__o21ai_1 _14746_ (.A1(_04719_),
    .A2(_05677_),
    .B1(_05678_),
    .Y(_00509_));
 sky130_fd_sc_hd__clkbuf_4 _14747_ (.A(_04236_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _14748_ (.A(_04672_),
    .B(_05230_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand2_1 _14749_ (.A(\samples_real[5][4] ),
    .B(_04673_),
    .Y(_05681_));
 sky130_fd_sc_hd__o211ai_1 _14750_ (.A1(_05633_),
    .A2(_05231_),
    .B1(_05681_),
    .C1(_04680_),
    .Y(_05682_));
 sky130_fd_sc_hd__a31oi_1 _14751_ (.A1(_05679_),
    .A2(_05682_),
    .A3(_05680_),
    .B1(_05237_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(\samples_real[5][4] ),
    .B(_04683_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_0 _14753_ (.A1(_04719_),
    .A2(_05683_),
    .B1(_05684_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _14754_ (.A(_04686_),
    .B(_05241_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_1 _14755_ (.A(\samples_real[5][5] ),
    .B(_04673_),
    .Y(_05686_));
 sky130_fd_sc_hd__o211ai_1 _14756_ (.A1(_05633_),
    .A2(_05242_),
    .B1(_05686_),
    .C1(_04679_),
    .Y(_05687_));
 sky130_fd_sc_hd__a31oi_1 _14757_ (.A1(_05679_),
    .A2(_05685_),
    .A3(_05687_),
    .B1(_05249_),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _14758_ (.A(\samples_real[5][5] ),
    .B(_04683_),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ai_0 _14759_ (.A1(_04719_),
    .A2(_05688_),
    .B1(_05689_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _14760_ (.A(_04686_),
    .B(_05253_),
    .Y(_05690_));
 sky130_fd_sc_hd__nand2_1 _14761_ (.A(\samples_real[5][6] ),
    .B(_04673_),
    .Y(_05691_));
 sky130_fd_sc_hd__o211ai_1 _14762_ (.A1(_05633_),
    .A2(_05254_),
    .B1(_05691_),
    .C1(_04679_),
    .Y(_05692_));
 sky130_fd_sc_hd__a31oi_1 _14763_ (.A1(_05679_),
    .A2(_05690_),
    .A3(_05692_),
    .B1(_05261_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_1 _14764_ (.A(\samples_real[5][6] ),
    .B(_04683_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_0 _14765_ (.A1(_04719_),
    .A2(_05693_),
    .B1(_05694_),
    .Y(_00512_));
 sky130_fd_sc_hd__nand2_1 _14766_ (.A(_04686_),
    .B(_05265_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _14767_ (.A(\samples_real[5][7] ),
    .B(_04673_),
    .Y(_05696_));
 sky130_fd_sc_hd__o211ai_2 _14768_ (.A1(_05634_),
    .A2(_05266_),
    .B1(_05696_),
    .C1(_04679_),
    .Y(_05697_));
 sky130_fd_sc_hd__a31oi_1 _14769_ (.A1(_05695_),
    .A2(_05697_),
    .A3(_05679_),
    .B1(_05272_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(\samples_real[5][7] ),
    .B(_04683_),
    .Y(_05699_));
 sky130_fd_sc_hd__o21ai_1 _14771_ (.A1(_04719_),
    .A2(_05698_),
    .B1(_05699_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _14772_ (.A(_04686_),
    .B(_05276_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _14773_ (.A(\samples_real[5][8] ),
    .B(_04673_),
    .Y(_05701_));
 sky130_fd_sc_hd__o211ai_2 _14774_ (.A1(_05277_),
    .A2(_05634_),
    .B1(_05701_),
    .C1(_04679_),
    .Y(_05702_));
 sky130_fd_sc_hd__a31oi_1 _14775_ (.A1(_05679_),
    .A2(_05700_),
    .A3(_05702_),
    .B1(_05283_),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_1 _14776_ (.A(\samples_real[5][8] ),
    .B(_04683_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_1 _14777_ (.A1(_04719_),
    .A2(_05703_),
    .B1(_05704_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_04686_),
    .B(_05287_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _14779_ (.A(\samples_real[5][9] ),
    .B(_04673_),
    .Y(_05706_));
 sky130_fd_sc_hd__o211ai_2 _14780_ (.A1(_05634_),
    .A2(_05288_),
    .B1(_05706_),
    .C1(_04679_),
    .Y(_05707_));
 sky130_fd_sc_hd__a31oi_1 _14781_ (.A1(_05679_),
    .A2(_05707_),
    .A3(_05705_),
    .B1(_05294_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _14782_ (.A(\samples_real[5][9] ),
    .B(_04683_),
    .Y(_05709_));
 sky130_fd_sc_hd__o21ai_1 _14783_ (.A1(_04719_),
    .A2(_05708_),
    .B1(_05709_),
    .Y(_00515_));
 sky130_fd_sc_hd__a22oi_2 _14784_ (.A1(\samples_real[6][0] ),
    .A2(_04797_),
    .B1(_05107_),
    .B2(_04787_),
    .Y(_05710_));
 sky130_fd_sc_hd__o22ai_1 _14785_ (.A1(_04791_),
    .A2(_05041_),
    .B1(_04795_),
    .B2(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__nor2_1 _14786_ (.A(_04784_),
    .B(_05113_),
    .Y(_05712_));
 sky130_fd_sc_hd__a221o_1 _14787_ (.A1(\samples_real[6][0] ),
    .A2(_04784_),
    .B1(_05711_),
    .B2(_04088_),
    .C1(_05712_),
    .X(_00516_));
 sky130_fd_sc_hd__clkbuf_4 _14788_ (.A(_03676_),
    .X(_05713_));
 sky130_fd_sc_hd__nand2_2 _14789_ (.A(_05713_),
    .B(_05125_),
    .Y(_05714_));
 sky130_fd_sc_hd__buf_2 _14790_ (.A(_04785_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_4 _14791_ (.A(_04785_),
    .X(_05716_));
 sky130_fd_sc_hd__nand2_1 _14792_ (.A(\samples_real[6][10] ),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__clkbuf_4 _14793_ (.A(_04790_),
    .X(_05718_));
 sky130_fd_sc_hd__o211ai_2 _14794_ (.A1(_05715_),
    .A2(_05127_),
    .B1(_05717_),
    .C1(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__a31oi_1 _14795_ (.A1(_05714_),
    .A2(_05719_),
    .A3(_05679_),
    .B1(_05133_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand2_1 _14796_ (.A(\samples_real[6][10] ),
    .B(_04874_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21ai_1 _14797_ (.A1(_04882_),
    .A2(_05720_),
    .B1(_05721_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _14798_ (.A(_05713_),
    .B(_05138_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _14799_ (.A(\samples_real[6][11] ),
    .B(_05716_),
    .Y(_05723_));
 sky130_fd_sc_hd__o211ai_2 _14800_ (.A1(_05715_),
    .A2(_05139_),
    .B1(_05723_),
    .C1(_05718_),
    .Y(_05724_));
 sky130_fd_sc_hd__a31oi_1 _14801_ (.A1(_05679_),
    .A2(_05724_),
    .A3(_05722_),
    .B1(_05145_),
    .Y(_05725_));
 sky130_fd_sc_hd__nand2_1 _14802_ (.A(\samples_real[6][11] ),
    .B(_04874_),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_1 _14803_ (.A1(_04882_),
    .A2(_05725_),
    .B1(_05726_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _14804_ (.A(_05713_),
    .B(_05151_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _14805_ (.A(\samples_real[6][12] ),
    .B(_05716_),
    .Y(_05728_));
 sky130_fd_sc_hd__o211ai_2 _14806_ (.A1(_05715_),
    .A2(_05152_),
    .B1(_05728_),
    .C1(_05718_),
    .Y(_05729_));
 sky130_fd_sc_hd__a31oi_1 _14807_ (.A1(_05679_),
    .A2(_05729_),
    .A3(_05727_),
    .B1(_05159_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_1 _14808_ (.A(\samples_real[6][12] ),
    .B(_04874_),
    .Y(_05731_));
 sky130_fd_sc_hd__o21ai_1 _14809_ (.A1(_04882_),
    .A2(_05730_),
    .B1(_05731_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _14810_ (.A(_05713_),
    .B(_05163_),
    .Y(_05732_));
 sky130_fd_sc_hd__nand2_1 _14811_ (.A(\samples_real[6][13] ),
    .B(_05716_),
    .Y(_05733_));
 sky130_fd_sc_hd__o211ai_2 _14812_ (.A1(_05715_),
    .A2(_05164_),
    .B1(_05733_),
    .C1(_05718_),
    .Y(_05734_));
 sky130_fd_sc_hd__a31oi_1 _14813_ (.A1(_05679_),
    .A2(_05734_),
    .A3(_05732_),
    .B1(_05171_),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _14814_ (.A(\samples_real[6][13] ),
    .B(_04874_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_1 _14815_ (.A1(_04882_),
    .A2(_05735_),
    .B1(_05736_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _14816_ (.A(_05713_),
    .B(_05177_),
    .Y(_05737_));
 sky130_fd_sc_hd__nand2_1 _14817_ (.A(\samples_real[6][14] ),
    .B(_05716_),
    .Y(_05738_));
 sky130_fd_sc_hd__o211ai_1 _14818_ (.A1(_05715_),
    .A2(_05178_),
    .B1(_05738_),
    .C1(_05718_),
    .Y(_05739_));
 sky130_fd_sc_hd__a31oi_1 _14819_ (.A1(_05324_),
    .A2(_05737_),
    .A3(_05739_),
    .B1(_05185_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_1 _14820_ (.A(\samples_real[6][14] ),
    .B(_04874_),
    .Y(_05741_));
 sky130_fd_sc_hd__o21ai_0 _14821_ (.A1(_04882_),
    .A2(_05740_),
    .B1(_05741_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand2_1 _14822_ (.A(\samples_real[6][15] ),
    .B(_04785_),
    .Y(_05742_));
 sky130_fd_sc_hd__o211ai_1 _14823_ (.A1(_04786_),
    .A2(_05188_),
    .B1(_05742_),
    .C1(_04790_),
    .Y(_05743_));
 sky130_fd_sc_hd__o21ai_0 _14824_ (.A1(_04790_),
    .A2(net593),
    .B1(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__a211oi_1 _14825_ (.A1(_04029_),
    .A2(_05744_),
    .B1(_05192_),
    .C1(_04833_),
    .Y(_05745_));
 sky130_fd_sc_hd__a21o_1 _14826_ (.A1(\samples_real[6][15] ),
    .A2(_04833_),
    .B1(_05745_),
    .X(_00522_));
 sky130_fd_sc_hd__nor2_4 _14827_ (.A(_05194_),
    .B(_04786_),
    .Y(_05746_));
 sky130_fd_sc_hd__a21oi_2 _14828_ (.A1(\samples_real[6][1] ),
    .A2(_04797_),
    .B1(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(_03676_),
    .B(_05198_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_2 _14830_ (.A1(_04800_),
    .A2(_05747_),
    .B1(_05748_),
    .Y(_05749_));
 sky130_fd_sc_hd__a21oi_1 _14831_ (.A1(_05596_),
    .A2(_05749_),
    .B1(_05202_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_1 _14832_ (.A(\samples_real[6][1] ),
    .B(_04874_),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_1 _14833_ (.A1(_04882_),
    .A2(_05750_),
    .B1(_05751_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _14834_ (.A(_05713_),
    .B(_05206_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_1 _14835_ (.A(\samples_real[6][2] ),
    .B(_05716_),
    .Y(_05753_));
 sky130_fd_sc_hd__o211ai_2 _14836_ (.A1(_05715_),
    .A2(_05207_),
    .B1(_05753_),
    .C1(_05718_),
    .Y(_05754_));
 sky130_fd_sc_hd__a31oi_1 _14837_ (.A1(_05324_),
    .A2(_05754_),
    .A3(_05752_),
    .B1(_05213_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _14838_ (.A(\samples_real[6][2] ),
    .B(_04794_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_1 _14839_ (.A1(_05755_),
    .A2(_04882_),
    .B1(_05756_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _14840_ (.A(_05713_),
    .B(_05218_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_1 _14841_ (.A(\samples_real[6][3] ),
    .B(_05716_),
    .Y(_05758_));
 sky130_fd_sc_hd__o211ai_2 _14842_ (.A1(_05715_),
    .A2(net619),
    .B1(_05758_),
    .C1(_05718_),
    .Y(_05759_));
 sky130_fd_sc_hd__a31oi_1 _14843_ (.A1(_05324_),
    .A2(_05759_),
    .A3(_05757_),
    .B1(_05226_),
    .Y(_05760_));
 sky130_fd_sc_hd__nand2_1 _14844_ (.A(\samples_real[6][3] ),
    .B(_04794_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_1 _14845_ (.A1(_05760_),
    .A2(_04882_),
    .B1(_05761_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _14846_ (.A(_05713_),
    .B(_05230_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _14847_ (.A(\samples_real[6][4] ),
    .B(_04796_),
    .Y(_05763_));
 sky130_fd_sc_hd__o211ai_1 _14848_ (.A1(_05715_),
    .A2(_05231_),
    .B1(_05763_),
    .C1(_05718_),
    .Y(_05764_));
 sky130_fd_sc_hd__a31oi_1 _14849_ (.A1(_05324_),
    .A2(_05764_),
    .A3(_05762_),
    .B1(_05237_),
    .Y(_05765_));
 sky130_fd_sc_hd__nand2_1 _14850_ (.A(\samples_real[6][4] ),
    .B(_04794_),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_0 _14851_ (.A1(_05765_),
    .A2(_04833_),
    .B1(_05766_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _14852_ (.A(_05713_),
    .B(_05241_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_1 _14853_ (.A(\samples_real[6][5] ),
    .B(_04796_),
    .Y(_05768_));
 sky130_fd_sc_hd__o211ai_1 _14854_ (.A1(_05715_),
    .A2(_05242_),
    .B1(_05768_),
    .C1(_05718_),
    .Y(_05769_));
 sky130_fd_sc_hd__a31oi_1 _14855_ (.A1(_05324_),
    .A2(_05767_),
    .A3(_05769_),
    .B1(_05249_),
    .Y(_05770_));
 sky130_fd_sc_hd__nand2_1 _14856_ (.A(\samples_real[6][5] ),
    .B(_04794_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_0 _14857_ (.A1(_04833_),
    .A2(_05770_),
    .B1(_05771_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _14858_ (.A(_05713_),
    .B(_05253_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2_1 _14859_ (.A(\samples_real[6][6] ),
    .B(_04796_),
    .Y(_05773_));
 sky130_fd_sc_hd__o211ai_1 _14860_ (.A1(_05715_),
    .A2(_05254_),
    .B1(_05773_),
    .C1(_05718_),
    .Y(_05774_));
 sky130_fd_sc_hd__a31oi_1 _14861_ (.A1(_05324_),
    .A2(_05772_),
    .A3(_05774_),
    .B1(_05261_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_1 _14862_ (.A(\samples_real[6][6] ),
    .B(_04794_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_0 _14863_ (.A1(_04833_),
    .A2(_05775_),
    .B1(_05776_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_2 _14864_ (.A(_05265_),
    .B(_04795_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _14865_ (.A(\samples_real[6][7] ),
    .B(_04796_),
    .Y(_05778_));
 sky130_fd_sc_hd__o211ai_2 _14866_ (.A1(_05716_),
    .A2(_05266_),
    .B1(_05778_),
    .C1(_04790_),
    .Y(_05779_));
 sky130_fd_sc_hd__a31oi_1 _14867_ (.A1(_05777_),
    .A2(_05779_),
    .A3(_05324_),
    .B1(_05272_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(\samples_real[6][7] ),
    .B(_04794_),
    .Y(_05781_));
 sky130_fd_sc_hd__o21ai_2 _14869_ (.A1(_04833_),
    .A2(_05780_),
    .B1(_05781_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _14870_ (.A(_04795_),
    .B(_05276_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _14871_ (.A(\samples_real[6][8] ),
    .B(_04796_),
    .Y(_05783_));
 sky130_fd_sc_hd__o211ai_2 _14872_ (.A1(_05277_),
    .A2(_05716_),
    .B1(_05783_),
    .C1(_04790_),
    .Y(_05784_));
 sky130_fd_sc_hd__a31oi_1 _14873_ (.A1(_05324_),
    .A2(_05782_),
    .A3(_05784_),
    .B1(_05283_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _14874_ (.A(\samples_real[6][8] ),
    .B(_04794_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_1 _14875_ (.A1(_04833_),
    .A2(_05785_),
    .B1(_05786_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _14876_ (.A(_04795_),
    .B(_05287_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_1 _14877_ (.A(\samples_real[6][9] ),
    .B(_04796_),
    .Y(_05788_));
 sky130_fd_sc_hd__o211ai_2 _14878_ (.A1(_05716_),
    .A2(_05288_),
    .B1(_05788_),
    .C1(_04790_),
    .Y(_05789_));
 sky130_fd_sc_hd__a31oi_1 _14879_ (.A1(_05324_),
    .A2(_05789_),
    .A3(_05787_),
    .B1(_05294_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _14880_ (.A(\samples_real[6][9] ),
    .B(_04794_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_1 _14881_ (.A1(_04833_),
    .A2(_05790_),
    .B1(_05791_),
    .Y(_00531_));
 sky130_fd_sc_hd__a22oi_1 _14882_ (.A1(\samples_real[7][0] ),
    .A2(_04901_),
    .B1(_05107_),
    .B2(_04902_),
    .Y(_05792_));
 sky130_fd_sc_hd__buf_2 _14883_ (.A(_04909_),
    .X(_05793_));
 sky130_fd_sc_hd__o22ai_1 _14884_ (.A1(_04905_),
    .A2(_05041_),
    .B1(_05793_),
    .B2(_05792_),
    .Y(_05794_));
 sky130_fd_sc_hd__nor2_1 _14885_ (.A(_04898_),
    .B(_05113_),
    .Y(_05795_));
 sky130_fd_sc_hd__a221o_1 _14886_ (.A1(\samples_real[7][0] ),
    .A2(_04898_),
    .B1(_05794_),
    .B2(_04088_),
    .C1(_05795_),
    .X(_00532_));
 sky130_fd_sc_hd__nor2_4 _14887_ (.A(_04949_),
    .B(_05127_),
    .Y(_05796_));
 sky130_fd_sc_hd__a211oi_1 _14888_ (.A1(\samples_real[7][10] ),
    .A2(_04984_),
    .B1(_04899_),
    .C1(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__a21oi_1 _14889_ (.A1(_05793_),
    .A2(_05125_),
    .B1(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__a21oi_1 _14890_ (.A1(_05798_),
    .A2(_05596_),
    .B1(_05133_),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_1 _14891_ (.A(\samples_real[7][10] ),
    .B(_04990_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_1 _14892_ (.A1(_04999_),
    .A2(_05799_),
    .B1(_05800_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_4 _14893_ (.A(_04949_),
    .B(_05139_),
    .Y(_05801_));
 sky130_fd_sc_hd__a211oi_2 _14894_ (.A1(\samples_real[7][11] ),
    .A2(_04984_),
    .B1(_04899_),
    .C1(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__a21oi_1 _14895_ (.A1(_05793_),
    .A2(_05138_),
    .B1(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__a21oi_1 _14896_ (.A1(_05803_),
    .A2(_05596_),
    .B1(_05145_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _14897_ (.A(\samples_real[7][11] ),
    .B(_04990_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_1 _14898_ (.A1(_04999_),
    .A2(_05804_),
    .B1(_05805_),
    .Y(_00534_));
 sky130_fd_sc_hd__clkbuf_4 _14899_ (.A(_04236_),
    .X(_05806_));
 sky130_fd_sc_hd__nor2_2 _14900_ (.A(_04949_),
    .B(_05152_),
    .Y(_05807_));
 sky130_fd_sc_hd__a211oi_1 _14901_ (.A1(\samples_real[7][12] ),
    .A2(_04984_),
    .B1(_04899_),
    .C1(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__a21oi_1 _14902_ (.A1(_05793_),
    .A2(_05151_),
    .B1(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__a21oi_1 _14903_ (.A1(_05806_),
    .A2(_05809_),
    .B1(_05159_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_1 _14904_ (.A(\samples_real[7][12] ),
    .B(_04990_),
    .Y(_05811_));
 sky130_fd_sc_hd__o21ai_1 _14905_ (.A1(_04999_),
    .A2(_05810_),
    .B1(_05811_),
    .Y(_00535_));
 sky130_fd_sc_hd__clkbuf_4 _14906_ (.A(_04900_),
    .X(_05812_));
 sky130_fd_sc_hd__nor2_4 _14907_ (.A(_05164_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__a211oi_2 _14908_ (.A1(\samples_real[7][13] ),
    .A2(_04984_),
    .B1(_04899_),
    .C1(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__a21oi_2 _14909_ (.A1(_05793_),
    .A2(_05163_),
    .B1(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__a21oi_1 _14910_ (.A1(_05815_),
    .A2(_05806_),
    .B1(_05171_),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2_1 _14911_ (.A(\samples_real[7][13] ),
    .B(_04990_),
    .Y(_05817_));
 sky130_fd_sc_hd__o21ai_1 _14912_ (.A1(_04999_),
    .A2(_05816_),
    .B1(_05817_),
    .Y(_00536_));
 sky130_fd_sc_hd__nor2_4 _14913_ (.A(_05812_),
    .B(_05178_),
    .Y(_05818_));
 sky130_fd_sc_hd__a211oi_2 _14914_ (.A1(\samples_real[7][14] ),
    .A2(_04984_),
    .B1(_04899_),
    .C1(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__a21oi_1 _14915_ (.A1(_05793_),
    .A2(_05177_),
    .B1(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__a21oi_1 _14916_ (.A1(_05806_),
    .A2(_05820_),
    .B1(_05185_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2_1 _14917_ (.A(\samples_real[7][14] ),
    .B(_04990_),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_1 _14918_ (.A1(_04999_),
    .A2(_05821_),
    .B1(_05822_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _14919_ (.A(\samples_real[7][15] ),
    .B(_04900_),
    .Y(_05823_));
 sky130_fd_sc_hd__o211ai_1 _14920_ (.A1(_04949_),
    .A2(_05188_),
    .B1(_05823_),
    .C1(_04904_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_0 _14921_ (.A1(_04904_),
    .A2(net52),
    .B1(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__a211oi_1 _14922_ (.A1(_04029_),
    .A2(_05825_),
    .B1(_05192_),
    .C1(_04948_),
    .Y(_05826_));
 sky130_fd_sc_hd__a21o_1 _14923_ (.A1(\samples_real[7][15] ),
    .A2(_04948_),
    .B1(_05826_),
    .X(_00538_));
 sky130_fd_sc_hd__nor2_4 _14924_ (.A(_05194_),
    .B(_04949_),
    .Y(_05827_));
 sky130_fd_sc_hd__a21oi_1 _14925_ (.A1(\samples_real[7][1] ),
    .A2(_04984_),
    .B1(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__nand2_1 _14926_ (.A(_04899_),
    .B(_05198_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_1 _14927_ (.A1(_04915_),
    .A2(_05828_),
    .B1(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21oi_1 _14928_ (.A1(_05830_),
    .A2(_05806_),
    .B1(_05202_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_1 _14929_ (.A(\samples_real[7][1] ),
    .B(_04990_),
    .Y(_05832_));
 sky130_fd_sc_hd__o21ai_1 _14930_ (.A1(_04999_),
    .A2(_05831_),
    .B1(_05832_),
    .Y(_00539_));
 sky130_fd_sc_hd__nor2_2 _14931_ (.A(_05812_),
    .B(_05207_),
    .Y(_05833_));
 sky130_fd_sc_hd__a211oi_1 _14932_ (.A1(\samples_real[7][2] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21oi_1 _14933_ (.A1(_05793_),
    .A2(_05206_),
    .B1(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__a21oi_1 _14934_ (.A1(_05806_),
    .A2(_05835_),
    .B1(_05213_),
    .Y(_05836_));
 sky130_fd_sc_hd__nand2_1 _14935_ (.A(\samples_real[7][2] ),
    .B(_04908_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_1 _14936_ (.A1(_04999_),
    .A2(_05836_),
    .B1(_05837_),
    .Y(_00540_));
 sky130_fd_sc_hd__nor2_4 _14937_ (.A(_05812_),
    .B(net619),
    .Y(_05838_));
 sky130_fd_sc_hd__a211oi_2 _14938_ (.A1(\samples_real[7][3] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__a21oi_1 _14939_ (.A1(_05793_),
    .A2(_05218_),
    .B1(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__a21oi_1 _14940_ (.A1(_05806_),
    .A2(_05840_),
    .B1(_05226_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_1 _14941_ (.A(\samples_real[7][3] ),
    .B(_04908_),
    .Y(_05842_));
 sky130_fd_sc_hd__o21ai_1 _14942_ (.A1(_04999_),
    .A2(_05841_),
    .B1(_05842_),
    .Y(_00541_));
 sky130_fd_sc_hd__nor2_2 _14943_ (.A(_05812_),
    .B(_05231_),
    .Y(_05843_));
 sky130_fd_sc_hd__a211oi_1 _14944_ (.A1(\samples_real[7][4] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__a21oi_1 _14945_ (.A1(_05793_),
    .A2(_05230_),
    .B1(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__a21oi_1 _14946_ (.A1(_05806_),
    .A2(_05845_),
    .B1(_05237_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _14947_ (.A(\samples_real[7][4] ),
    .B(_04908_),
    .Y(_05847_));
 sky130_fd_sc_hd__o21ai_1 _14948_ (.A1(_04948_),
    .A2(_05846_),
    .B1(_05847_),
    .Y(_00542_));
 sky130_fd_sc_hd__nor2_4 _14949_ (.A(_05812_),
    .B(_05242_),
    .Y(_05848_));
 sky130_fd_sc_hd__a211oi_2 _14950_ (.A1(\samples_real[7][5] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__a21oi_1 _14951_ (.A1(_05793_),
    .A2(_05241_),
    .B1(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__a21oi_1 _14952_ (.A1(_05806_),
    .A2(_05850_),
    .B1(_05249_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_1 _14953_ (.A(\samples_real[7][5] ),
    .B(_04908_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_1 _14954_ (.A1(_04948_),
    .A2(_05851_),
    .B1(_05852_),
    .Y(_00543_));
 sky130_fd_sc_hd__nor2_2 _14955_ (.A(_05812_),
    .B(_05254_),
    .Y(_05853_));
 sky130_fd_sc_hd__a211oi_1 _14956_ (.A1(\samples_real[7][6] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__a21oi_1 _14957_ (.A1(_04910_),
    .A2(_05253_),
    .B1(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__a21oi_1 _14958_ (.A1(_05806_),
    .A2(_05855_),
    .B1(_05261_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _14959_ (.A(\samples_real[7][6] ),
    .B(_04908_),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_1 _14960_ (.A1(_04948_),
    .A2(_05856_),
    .B1(_05857_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_4 _14961_ (.A(_05266_),
    .B(_05812_),
    .Y(_05858_));
 sky130_fd_sc_hd__a211oi_1 _14962_ (.A1(\samples_real[7][7] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__a21oi_1 _14963_ (.A1(_04910_),
    .A2(_05265_),
    .B1(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__a21oi_1 _14964_ (.A1(_05860_),
    .A2(_05806_),
    .B1(_05272_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _14965_ (.A(\samples_real[7][7] ),
    .B(_04908_),
    .Y(_05862_));
 sky130_fd_sc_hd__o21ai_1 _14966_ (.A1(_04948_),
    .A2(_05861_),
    .B1(_05862_),
    .Y(_00545_));
 sky130_fd_sc_hd__nor2_4 _14967_ (.A(_05812_),
    .B(_05277_),
    .Y(_05863_));
 sky130_fd_sc_hd__a211oi_2 _14968_ (.A1(\samples_real[7][8] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__a21oi_1 _14969_ (.A1(_04910_),
    .A2(_05276_),
    .B1(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21oi_1 _14970_ (.A1(_04237_),
    .A2(_05865_),
    .B1(_05283_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _14971_ (.A(\samples_real[7][8] ),
    .B(_04908_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_1 _14972_ (.A1(_04948_),
    .A2(_05866_),
    .B1(_05867_),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_4 _14973_ (.A(_05812_),
    .B(_05288_),
    .Y(_05868_));
 sky130_fd_sc_hd__a211oi_2 _14974_ (.A1(\samples_real[7][9] ),
    .A2(_04901_),
    .B1(_04909_),
    .C1(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__a21oi_1 _14975_ (.A1(_04910_),
    .A2(_05287_),
    .B1(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__a21oi_1 _14976_ (.A1(_04237_),
    .A2(_05870_),
    .B1(_05294_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _14977_ (.A(\samples_real[7][9] ),
    .B(_04908_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_1 _14978_ (.A1(_04948_),
    .A2(_05871_),
    .B1(_05872_),
    .Y(_00547_));
 sky130_fd_sc_hd__a21boi_2 _14979_ (.A1(_07819_),
    .A2(_03144_),
    .B1_N(_03846_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand3_1 _14980_ (.A(_04004_),
    .B(_07803_),
    .C(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__o21ai_0 _14981_ (.A1(_07803_),
    .A2(_05873_),
    .B1(_05874_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand3_1 _14982_ (.A(_04004_),
    .B(_07806_),
    .C(_05873_),
    .Y(_05875_));
 sky130_fd_sc_hd__o21ai_0 _14983_ (.A1(_07804_),
    .A2(_05873_),
    .B1(_05875_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand3_1 _14984_ (.A(_04004_),
    .B(_07820_),
    .C(_05873_),
    .Y(_05876_));
 sky130_fd_sc_hd__o21ai_0 _14985_ (.A1(_07817_),
    .A2(_05873_),
    .B1(_05876_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2b_1 _14986_ (.A_N(_00002_),
    .B(_03192_),
    .Y(_00021_));
 sky130_fd_sc_hd__fa_2 _14987_ (.A(_05882_),
    .B(_05883_),
    .CIN(_05884_),
    .COUT(_05885_),
    .SUM(_05886_));
 sky130_fd_sc_hd__fa_2 _14988_ (.A(_05882_),
    .B(net588),
    .CIN(_05888_),
    .COUT(_05889_),
    .SUM(_05890_));
 sky130_fd_sc_hd__fa_1 _14989_ (.A(_05892_),
    .B(_05893_),
    .CIN(_05894_),
    .COUT(_05895_),
    .SUM(_05896_));
 sky130_fd_sc_hd__fa_2 _14990_ (.A(_05897_),
    .B(_05898_),
    .CIN(_05899_),
    .COUT(_05900_),
    .SUM(_05901_));
 sky130_fd_sc_hd__fa_2 _14991_ (.A(_05897_),
    .B(_05902_),
    .CIN(_05903_),
    .COUT(_05904_),
    .SUM(_05905_));
 sky130_fd_sc_hd__fa_1 _14992_ (.A(_05907_),
    .B(_05880_),
    .CIN(_05908_),
    .COUT(_05909_),
    .SUM(_05910_));
 sky130_fd_sc_hd__fa_1 _14993_ (.A(_05911_),
    .B(_05912_),
    .CIN(_05913_),
    .COUT(_05914_),
    .SUM(_05915_));
 sky130_fd_sc_hd__fa_1 _14994_ (.A(_05916_),
    .B(_05917_),
    .CIN(_05918_),
    .COUT(_05919_),
    .SUM(_05920_));
 sky130_fd_sc_hd__fa_1 _14995_ (.A(_05921_),
    .B(_05922_),
    .CIN(_05923_),
    .COUT(_05917_),
    .SUM(_05924_));
 sky130_fd_sc_hd__fa_1 _14996_ (.A(_05925_),
    .B(_05926_),
    .CIN(_05927_),
    .COUT(_05928_),
    .SUM(_05929_));
 sky130_fd_sc_hd__fa_1 _14997_ (.A(_05920_),
    .B(_05930_),
    .CIN(_05931_),
    .COUT(_05932_),
    .SUM(_05933_));
 sky130_fd_sc_hd__fa_1 _14998_ (.A(_05924_),
    .B(_05934_),
    .CIN(_05935_),
    .COUT(_05930_),
    .SUM(_05936_));
 sky130_fd_sc_hd__fa_1 _14999_ (.A(_05937_),
    .B(_05938_),
    .CIN(_05939_),
    .COUT(_05940_),
    .SUM(_05941_));
 sky130_fd_sc_hd__fa_1 _15000_ (.A(_05942_),
    .B(_05943_),
    .CIN(_05944_),
    .COUT(_05945_),
    .SUM(_05946_));
 sky130_fd_sc_hd__fa_1 _15001_ (.A(_05947_),
    .B(_05948_),
    .CIN(_05949_),
    .COUT(_05950_),
    .SUM(_05951_));
 sky130_fd_sc_hd__fa_1 _15002_ (.A(_05952_),
    .B(_05953_),
    .CIN(_05954_),
    .COUT(_05955_),
    .SUM(_05956_));
 sky130_fd_sc_hd__fa_1 _15003_ (.A(_05923_),
    .B(_05957_),
    .CIN(_05958_),
    .COUT(_05959_),
    .SUM(_05960_));
 sky130_fd_sc_hd__fa_1 _15004_ (.A(_05961_),
    .B(net454),
    .CIN(_05963_),
    .COUT(_05964_),
    .SUM(_05965_));
 sky130_fd_sc_hd__fa_1 _15005_ (.A(_05960_),
    .B(_05966_),
    .CIN(_05965_),
    .COUT(_05967_),
    .SUM(_05968_));
 sky130_fd_sc_hd__fa_1 _15006_ (.A(_05970_),
    .B(_05969_),
    .CIN(_05933_),
    .COUT(_05971_),
    .SUM(_05972_));
 sky130_fd_sc_hd__fa_1 _15007_ (.A(_05936_),
    .B(_05973_),
    .CIN(_05974_),
    .COUT(_05969_),
    .SUM(_05975_));
 sky130_fd_sc_hd__fa_1 _15008_ (.A(_05976_),
    .B(_05977_),
    .CIN(_05978_),
    .COUT(_05973_),
    .SUM(_05979_));
 sky130_fd_sc_hd__fa_1 _15009_ (.A(_05938_),
    .B(_05980_),
    .CIN(_05981_),
    .COUT(_05982_),
    .SUM(_05983_));
 sky130_fd_sc_hd__fa_1 _15010_ (.A(_05984_),
    .B(_05985_),
    .CIN(_05986_),
    .COUT(_05987_),
    .SUM(_05988_));
 sky130_fd_sc_hd__fa_1 _15011_ (.A(_05989_),
    .B(_05990_),
    .CIN(_05991_),
    .COUT(_05992_),
    .SUM(_05993_));
 sky130_fd_sc_hd__fa_1 _15012_ (.A(_05994_),
    .B(_05995_),
    .CIN(_05996_),
    .COUT(_05997_),
    .SUM(_05998_));
 sky130_fd_sc_hd__fa_1 _15013_ (.A(_05939_),
    .B(_05981_),
    .CIN(_05999_),
    .COUT(_06000_),
    .SUM(_06001_));
 sky130_fd_sc_hd__fa_1 _15014_ (.A(_06003_),
    .B(_06004_),
    .CIN(_06005_),
    .COUT(_06006_),
    .SUM(_06007_));
 sky130_fd_sc_hd__fa_1 _15015_ (.A(_06001_),
    .B(_06008_),
    .CIN(_06007_),
    .COUT(_06009_),
    .SUM(_06010_));
 sky130_fd_sc_hd__fa_1 _15016_ (.A(_06012_),
    .B(_06013_),
    .CIN(_06014_),
    .COUT(_06015_),
    .SUM(_06016_));
 sky130_fd_sc_hd__fa_1 _15017_ (.A(_06018_),
    .B(_06017_),
    .CIN(_06019_),
    .COUT(_06020_),
    .SUM(_06021_));
 sky130_fd_sc_hd__fa_1 _15018_ (.A(_06022_),
    .B(_06024_),
    .CIN(_06023_),
    .COUT(_06025_),
    .SUM(_06026_));
 sky130_fd_sc_hd__fa_1 _15019_ (.A(_06019_),
    .B(_06027_),
    .CIN(_06028_),
    .COUT(_06029_),
    .SUM(_06030_));
 sky130_fd_sc_hd__fa_2 _15020_ (.A(_06031_),
    .B(_06032_),
    .CIN(_06033_),
    .COUT(_06034_),
    .SUM(_06035_));
 sky130_fd_sc_hd__fa_1 _15021_ (.A(_06036_),
    .B(_06037_),
    .CIN(_06026_),
    .COUT(_06038_),
    .SUM(_06039_));
 sky130_fd_sc_hd__fa_1 _15022_ (.A(_05958_),
    .B(_06002_),
    .CIN(net454),
    .COUT(_06011_),
    .SUM(_06040_));
 sky130_fd_sc_hd__fa_1 _15023_ (.A(_05963_),
    .B(net449),
    .CIN(_06031_),
    .COUT(_06042_),
    .SUM(_06043_));
 sky130_fd_sc_hd__fa_1 _15024_ (.A(_06042_),
    .B(_06030_),
    .CIN(_06044_),
    .COUT(_06037_),
    .SUM(_06045_));
 sky130_fd_sc_hd__fa_1 _15025_ (.A(_06028_),
    .B(_06046_),
    .CIN(_06047_),
    .COUT(_06048_),
    .SUM(_06049_));
 sky130_fd_sc_hd__fa_1 _15026_ (.A(_06050_),
    .B(_06051_),
    .CIN(_06052_),
    .COUT(_06053_),
    .SUM(_06054_));
 sky130_fd_sc_hd__fa_1 _15027_ (.A(_06056_),
    .B(_06055_),
    .CIN(_05972_),
    .COUT(_06057_),
    .SUM(_06058_));
 sky130_fd_sc_hd__fa_1 _15028_ (.A(_05975_),
    .B(_06059_),
    .CIN(_06060_),
    .COUT(_06055_),
    .SUM(_06061_));
 sky130_fd_sc_hd__fa_1 _15029_ (.A(_05979_),
    .B(_06062_),
    .CIN(_06063_),
    .COUT(_06059_),
    .SUM(_06064_));
 sky130_fd_sc_hd__fa_1 _15030_ (.A(_06065_),
    .B(_06066_),
    .CIN(_06067_),
    .COUT(_06062_),
    .SUM(_06068_));
 sky130_fd_sc_hd__fa_1 _15031_ (.A(_06069_),
    .B(_06070_),
    .CIN(_06002_),
    .COUT(_06066_),
    .SUM(_06071_));
 sky130_fd_sc_hd__fa_1 _15032_ (.A(_06072_),
    .B(_06073_),
    .CIN(_06074_),
    .COUT(_06075_),
    .SUM(_06076_));
 sky130_fd_sc_hd__fa_1 _15033_ (.A(_06077_),
    .B(_06078_),
    .CIN(_06010_),
    .COUT(_06014_),
    .SUM(_06079_));
 sky130_fd_sc_hd__fa_1 _15034_ (.A(_05957_),
    .B(_06080_),
    .CIN(_06081_),
    .COUT(_06082_),
    .SUM(_06083_));
 sky130_fd_sc_hd__fa_1 _15035_ (.A(_06040_),
    .B(_06084_),
    .CIN(_06085_),
    .COUT(_06086_),
    .SUM(_06087_));
 sky130_fd_sc_hd__fa_1 _15036_ (.A(_06054_),
    .B(_06088_),
    .CIN(_06039_),
    .COUT(_06089_),
    .SUM(_06090_));
 sky130_fd_sc_hd__fa_1 _15037_ (.A(_06086_),
    .B(_06092_),
    .CIN(_06091_),
    .COUT(_06088_),
    .SUM(_06093_));
 sky130_fd_sc_hd__fa_1 _15038_ (.A(_06002_),
    .B(net454),
    .CIN(_06095_),
    .COUT(_06084_),
    .SUM(_06096_));
 sky130_fd_sc_hd__fa_1 _15039_ (.A(_06005_),
    .B(_06019_),
    .CIN(_06027_),
    .COUT(_06097_),
    .SUM(_06098_));
 sky130_fd_sc_hd__fa_1 _15040_ (.A(_06099_),
    .B(_06097_),
    .CIN(_06100_),
    .COUT(_06094_),
    .SUM(_06101_));
 sky130_fd_sc_hd__fa_1 _15041_ (.A(_06102_),
    .B(_06103_),
    .CIN(_06090_),
    .COUT(_06104_),
    .SUM(_06105_));
 sky130_fd_sc_hd__fa_1 _15042_ (.A(_06058_),
    .B(_06107_),
    .CIN(_06108_),
    .COUT(_06109_),
    .SUM(_06110_));
 sky130_fd_sc_hd__fa_1 _15043_ (.A(_06061_),
    .B(_06111_),
    .CIN(_06112_),
    .COUT(_06107_),
    .SUM(_06113_));
 sky130_fd_sc_hd__fa_1 _15044_ (.A(_06064_),
    .B(_06115_),
    .CIN(_06075_),
    .COUT(_06111_),
    .SUM(_06116_));
 sky130_fd_sc_hd__fa_1 _15045_ (.A(_06068_),
    .B(_06117_),
    .CIN(_06118_),
    .COUT(_06115_),
    .SUM(_06119_));
 sky130_fd_sc_hd__fa_1 _15046_ (.A(_06071_),
    .B(_06120_),
    .CIN(_06121_),
    .COUT(_06117_),
    .SUM(_06122_));
 sky130_fd_sc_hd__fa_1 _15047_ (.A(_06123_),
    .B(_06124_),
    .CIN(_06125_),
    .COUT(_06126_),
    .SUM(_06127_));
 sky130_fd_sc_hd__fa_1 _15048_ (.A(_06128_),
    .B(_06129_),
    .CIN(_06130_),
    .COUT(_06131_),
    .SUM(_06132_));
 sky130_fd_sc_hd__fa_1 _15049_ (.A(_05958_),
    .B(_06133_),
    .CIN(_06134_),
    .COUT(_06135_),
    .SUM(_06136_));
 sky130_fd_sc_hd__fa_1 _15050_ (.A(_06096_),
    .B(_06137_),
    .CIN(_06098_),
    .COUT(_06138_),
    .SUM(_06139_));
 sky130_fd_sc_hd__fa_1 _15051_ (.A(_06142_),
    .B(_06141_),
    .CIN(_06093_),
    .COUT(_06103_),
    .SUM(_06143_));
 sky130_fd_sc_hd__fa_1 _15052_ (.A(_06138_),
    .B(_06144_),
    .CIN(_06145_),
    .COUT(_06141_),
    .SUM(_06146_));
 sky130_fd_sc_hd__fa_1 _15053_ (.A(_06125_),
    .B(_06004_),
    .CIN(_06017_),
    .COUT(_06140_),
    .SUM(_06147_));
 sky130_fd_sc_hd__fa_1 _15054_ (.A(_06148_),
    .B(_06143_),
    .CIN(_06149_),
    .COUT(_06150_),
    .SUM(_06151_));
 sky130_fd_sc_hd__fa_1 _15055_ (.A(_06154_),
    .B(_06153_),
    .CIN(_06110_),
    .COUT(_06155_),
    .SUM(_06156_));
 sky130_fd_sc_hd__fa_1 _15056_ (.A(_06113_),
    .B(_06157_),
    .CIN(_06158_),
    .COUT(_06153_),
    .SUM(_06159_));
 sky130_fd_sc_hd__fa_1 _15057_ (.A(_06116_),
    .B(_06160_),
    .CIN(_06161_),
    .COUT(_06157_),
    .SUM(_06162_));
 sky130_fd_sc_hd__fa_1 _15058_ (.A(_06119_),
    .B(_06164_),
    .CIN(_06165_),
    .COUT(_06160_),
    .SUM(_06166_));
 sky130_fd_sc_hd__fa_1 _15059_ (.A(_06122_),
    .B(_06168_),
    .CIN(_06169_),
    .COUT(_06164_),
    .SUM(_06170_));
 sky130_fd_sc_hd__fa_1 _15060_ (.A(_06171_),
    .B(_06172_),
    .CIN(_06173_),
    .COUT(_06168_),
    .SUM(_06174_));
 sky130_fd_sc_hd__fa_1 _15061_ (.A(_06175_),
    .B(_06124_),
    .CIN(_06004_),
    .COUT(_06176_),
    .SUM(_06177_));
 sky130_fd_sc_hd__fa_1 _15062_ (.A(_06178_),
    .B(_06179_),
    .CIN(_06180_),
    .COUT(_06181_),
    .SUM(_06182_));
 sky130_fd_sc_hd__fa_1 _15063_ (.A(_05999_),
    .B(_06183_),
    .CIN(_06184_),
    .COUT(_06185_),
    .SUM(_06186_));
 sky130_fd_sc_hd__fa_1 _15064_ (.A(_06187_),
    .B(_06188_),
    .CIN(_06035_),
    .COUT(_06189_),
    .SUM(_06190_));
 sky130_fd_sc_hd__fa_1 _15065_ (.A(_06146_),
    .B(_06192_),
    .CIN(_06193_),
    .COUT(_06149_),
    .SUM(_06194_));
 sky130_fd_sc_hd__fa_1 _15066_ (.A(_06189_),
    .B(_06195_),
    .CIN(_06196_),
    .COUT(_06192_),
    .SUM(_06197_));
 sky130_fd_sc_hd__fa_1 _15067_ (.A(_06004_),
    .B(_06017_),
    .CIN(_06027_),
    .COUT(_06191_),
    .SUM(_06198_));
 sky130_fd_sc_hd__fa_1 _15068_ (.A(_06200_),
    .B(_06201_),
    .CIN(_06202_),
    .COUT(_06203_),
    .SUM(_06204_));
 sky130_fd_sc_hd__fa_1 _15069_ (.A(_06205_),
    .B(_06206_),
    .CIN(_06207_),
    .COUT(_06208_),
    .SUM(_06209_));
 sky130_fd_sc_hd__fa_2 _15070_ (.A(_06211_),
    .B(_06210_),
    .CIN(_06156_),
    .COUT(_06212_),
    .SUM(_06213_));
 sky130_fd_sc_hd__fa_2 _15071_ (.A(_06159_),
    .B(_06214_),
    .CIN(_06215_),
    .COUT(_06210_),
    .SUM(_06216_));
 sky130_fd_sc_hd__fa_1 _15072_ (.A(_06162_),
    .B(_06217_),
    .CIN(_06218_),
    .COUT(_06214_),
    .SUM(_06219_));
 sky130_fd_sc_hd__fa_1 _15073_ (.A(_06166_),
    .B(_06220_),
    .CIN(_06221_),
    .COUT(_06217_),
    .SUM(_06222_));
 sky130_fd_sc_hd__fa_1 _15074_ (.A(_06170_),
    .B(_06224_),
    .CIN(_06225_),
    .COUT(_06220_),
    .SUM(_06226_));
 sky130_fd_sc_hd__fa_1 _15075_ (.A(_06174_),
    .B(_06228_),
    .CIN(_06229_),
    .COUT(_06224_),
    .SUM(_06230_));
 sky130_fd_sc_hd__fa_1 _15076_ (.A(_06231_),
    .B(_06232_),
    .CIN(_06233_),
    .COUT(_06228_),
    .SUM(_06234_));
 sky130_fd_sc_hd__fa_1 _15077_ (.A(_06017_),
    .B(_06235_),
    .CIN(_06175_),
    .COUT(_06236_),
    .SUM(_06237_));
 sky130_fd_sc_hd__fa_1 _15078_ (.A(_06238_),
    .B(_06239_),
    .CIN(_06240_),
    .COUT(_06241_),
    .SUM(_06242_));
 sky130_fd_sc_hd__fa_1 _15079_ (.A(net453),
    .B(_06243_),
    .CIN(_06244_),
    .COUT(_06245_),
    .SUM(_06246_));
 sky130_fd_sc_hd__fa_1 _15080_ (.A(_06247_),
    .B(_06248_),
    .CIN(_06204_),
    .COUT(_06249_),
    .SUM(_06250_));
 sky130_fd_sc_hd__fa_1 _15081_ (.A(_06251_),
    .B(_06252_),
    .CIN(_06253_),
    .COUT(_06207_),
    .SUM(_06254_));
 sky130_fd_sc_hd__fa_1 _15082_ (.A(_06199_),
    .B(net450),
    .CIN(_06033_),
    .COUT(_06248_),
    .SUM(_06255_));
 sky130_fd_sc_hd__fa_1 _15083_ (.A(_06256_),
    .B(_06254_),
    .CIN(_06257_),
    .COUT(_06258_),
    .SUM(_06259_));
 sky130_fd_sc_hd__fa_1 _15084_ (.A(_06216_),
    .B(_06260_),
    .CIN(_06261_),
    .COUT(_06262_),
    .SUM(_06263_));
 sky130_fd_sc_hd__fa_1 _15085_ (.A(_06219_),
    .B(_06264_),
    .CIN(_06265_),
    .COUT(_06260_),
    .SUM(_06266_));
 sky130_fd_sc_hd__fa_1 _15086_ (.A(_06222_),
    .B(_06267_),
    .CIN(_06268_),
    .COUT(_06264_),
    .SUM(_06269_));
 sky130_fd_sc_hd__fa_1 _15087_ (.A(_06226_),
    .B(_06270_),
    .CIN(_06271_),
    .COUT(_06267_),
    .SUM(_06272_));
 sky130_fd_sc_hd__fa_1 _15088_ (.A(_06230_),
    .B(_06274_),
    .CIN(_06275_),
    .COUT(_06270_),
    .SUM(_06276_));
 sky130_fd_sc_hd__fa_1 _15089_ (.A(_06234_),
    .B(_06278_),
    .CIN(_06279_),
    .COUT(_06274_),
    .SUM(_06280_));
 sky130_fd_sc_hd__fa_1 _15090_ (.A(_06283_),
    .B(_06282_),
    .CIN(_06281_),
    .COUT(_06278_),
    .SUM(_06284_));
 sky130_fd_sc_hd__fa_1 _15091_ (.A(_06285_),
    .B(_06286_),
    .CIN(_06199_),
    .COUT(_06282_),
    .SUM(_06287_));
 sky130_fd_sc_hd__fa_1 _15092_ (.A(_06288_),
    .B(_06289_),
    .CIN(_06290_),
    .COUT(_06291_),
    .SUM(_06292_));
 sky130_fd_sc_hd__fa_1 _15093_ (.A(_06095_),
    .B(_06293_),
    .CIN(_06294_),
    .COUT(_06295_),
    .SUM(_06296_));
 sky130_fd_sc_hd__fa_1 _15094_ (.A(_06255_),
    .B(_06297_),
    .CIN(_06298_),
    .COUT(_06299_),
    .SUM(_06300_));
 sky130_fd_sc_hd__fa_1 _15095_ (.A(_06301_),
    .B(_06302_),
    .CIN(_06303_),
    .COUT(_06257_),
    .SUM(_06304_));
 sky130_fd_sc_hd__fa_1 _15096_ (.A(_06305_),
    .B(_06306_),
    .CIN(_06307_),
    .COUT(_06308_),
    .SUM(_06309_));
 sky130_fd_sc_hd__fa_1 _15097_ (.A(_06266_),
    .B(_06311_),
    .CIN(_06312_),
    .COUT(_06313_),
    .SUM(_06314_));
 sky130_fd_sc_hd__fa_1 _15098_ (.A(_06269_),
    .B(_06315_),
    .CIN(_06316_),
    .COUT(_06311_),
    .SUM(_06317_));
 sky130_fd_sc_hd__fa_1 _15099_ (.A(_06272_),
    .B(_06318_),
    .CIN(_06309_),
    .COUT(_06315_),
    .SUM(_06319_));
 sky130_fd_sc_hd__fa_1 _15100_ (.A(_06276_),
    .B(_06320_),
    .CIN(_06321_),
    .COUT(_06318_),
    .SUM(_06322_));
 sky130_fd_sc_hd__fa_1 _15101_ (.A(_06326_),
    .B(_06325_),
    .CIN(_06284_),
    .COUT(_06327_),
    .SUM(_06328_));
 sky130_fd_sc_hd__fa_1 _15102_ (.A(_06287_),
    .B(_06330_),
    .CIN(_06331_),
    .COUT(_06325_),
    .SUM(_06332_));
 sky130_fd_sc_hd__fa_1 _15103_ (.A(_06286_),
    .B(_06333_),
    .CIN(_06033_),
    .COUT(_06330_),
    .SUM(_06334_));
 sky130_fd_sc_hd__fa_1 _15104_ (.A(_06335_),
    .B(_06337_),
    .CIN(_06336_),
    .COUT(_06338_),
    .SUM(_06339_));
 sky130_fd_sc_hd__fa_1 _15105_ (.A(_06341_),
    .B(_06340_),
    .CIN(net448),
    .COUT(_06342_),
    .SUM(_06343_));
 sky130_fd_sc_hd__fa_1 _15106_ (.A(_06199_),
    .B(_06033_),
    .CIN(_06202_),
    .COUT(_06297_),
    .SUM(_06344_));
 sky130_fd_sc_hd__fa_1 _15107_ (.A(_06201_),
    .B(_06344_),
    .CIN(_06345_),
    .COUT(_06346_),
    .SUM(_06347_));
 sky130_fd_sc_hd__fa_1 _15108_ (.A(_06348_),
    .B(_06349_),
    .CIN(_06350_),
    .COUT(_06351_),
    .SUM(_06352_));
 sky130_fd_sc_hd__fa_1 _15109_ (.A(_06317_),
    .B(_06353_),
    .CIN(_06354_),
    .COUT(_06355_),
    .SUM(_06356_));
 sky130_fd_sc_hd__fa_1 _15110_ (.A(_06319_),
    .B(_06357_),
    .CIN(_06358_),
    .COUT(_06353_),
    .SUM(_06359_));
 sky130_fd_sc_hd__fa_1 _15111_ (.A(_06322_),
    .B(_06360_),
    .CIN(_06352_),
    .COUT(_06357_),
    .SUM(_06361_));
 sky130_fd_sc_hd__fa_1 _15112_ (.A(_06363_),
    .B(_06364_),
    .CIN(_06365_),
    .COUT(_06362_),
    .SUM(_06366_));
 sky130_fd_sc_hd__fa_1 _15113_ (.A(_06367_),
    .B(_06334_),
    .CIN(_06368_),
    .COUT(_06369_),
    .SUM(_06370_));
 sky130_fd_sc_hd__fa_1 _15114_ (.A(_06373_),
    .B(_06374_),
    .CIN(_06375_),
    .COUT(_06376_),
    .SUM(_06377_));
 sky130_fd_sc_hd__fa_1 _15115_ (.A(_06027_),
    .B(_06378_),
    .CIN(_06379_),
    .COUT(_06380_),
    .SUM(_06381_));
 sky130_fd_sc_hd__fa_1 _15116_ (.A(_06033_),
    .B(_06202_),
    .CIN(_06382_),
    .COUT(_06345_),
    .SUM(_06383_));
 sky130_fd_sc_hd__fa_1 _15117_ (.A(_06384_),
    .B(_06385_),
    .CIN(_06386_),
    .COUT(_06387_),
    .SUM(_06388_));
 sky130_fd_sc_hd__fa_1 _15118_ (.A(_06359_),
    .B(_06389_),
    .CIN(_06390_),
    .COUT(_06391_),
    .SUM(_06392_));
 sky130_fd_sc_hd__fa_1 _15119_ (.A(_06361_),
    .B(_06393_),
    .CIN(_06394_),
    .COUT(_06389_),
    .SUM(_06395_));
 sky130_fd_sc_hd__fa_1 _15120_ (.A(_06388_),
    .B(_06397_),
    .CIN(_06396_),
    .COUT(_06393_),
    .SUM(_06398_));
 sky130_fd_sc_hd__fa_1 _15121_ (.A(_06400_),
    .B(_06401_),
    .CIN(_06402_),
    .COUT(_06399_),
    .SUM(_06403_));
 sky130_fd_sc_hd__fa_1 _15122_ (.A(_06404_),
    .B(_06405_),
    .CIN(_06406_),
    .COUT(_06407_),
    .SUM(_06408_));
 sky130_fd_sc_hd__fa_1 _15123_ (.A(_06411_),
    .B(_06412_),
    .CIN(_06413_),
    .COUT(_06414_),
    .SUM(_06415_));
 sky130_fd_sc_hd__fa_1 _15124_ (.A(_06395_),
    .B(_06416_),
    .CIN(_06417_),
    .COUT(_06418_),
    .SUM(_06419_));
 sky130_fd_sc_hd__fa_1 _15125_ (.A(_06421_),
    .B(_06398_),
    .CIN(_06420_),
    .COUT(_06416_),
    .SUM(_06422_));
 sky130_fd_sc_hd__fa_1 _15126_ (.A(_06424_),
    .B(_06423_),
    .CIN(_06415_),
    .COUT(_06420_),
    .SUM(_06425_));
 sky130_fd_sc_hd__fa_1 _15127_ (.A(_06427_),
    .B(_06428_),
    .CIN(_06429_),
    .COUT(_06430_),
    .SUM(_06431_));
 sky130_fd_sc_hd__fa_1 _15128_ (.A(_06434_),
    .B(_06435_),
    .CIN(_06436_),
    .COUT(_06437_),
    .SUM(_06438_));
 sky130_fd_sc_hd__fa_1 _15129_ (.A(_06440_),
    .B(_06439_),
    .CIN(_06422_),
    .COUT(_06441_),
    .SUM(_06442_));
 sky130_fd_sc_hd__fa_1 _15130_ (.A(_06444_),
    .B(_06443_),
    .CIN(_06425_),
    .COUT(_06439_),
    .SUM(_06445_));
 sky130_fd_sc_hd__fa_1 _15131_ (.A(_06446_),
    .B(_06447_),
    .CIN(_06448_),
    .COUT(_06443_),
    .SUM(_06449_));
 sky130_fd_sc_hd__fa_1 _15132_ (.A(_06367_),
    .B(_06452_),
    .CIN(_06453_),
    .COUT(_06454_),
    .SUM(_06455_));
 sky130_fd_sc_hd__fa_1 _15133_ (.A(_06458_),
    .B(_06459_),
    .CIN(_06460_),
    .COUT(_06461_),
    .SUM(_06462_));
 sky130_fd_sc_hd__fa_1 _15134_ (.A(_06465_),
    .B(_06466_),
    .CIN(_06467_),
    .COUT(_06468_),
    .SUM(_06469_));
 sky130_fd_sc_hd__fa_1 _15135_ (.A(_06471_),
    .B(_06470_),
    .CIN(_06445_),
    .COUT(_06472_),
    .SUM(_06473_));
 sky130_fd_sc_hd__fa_1 _15136_ (.A(_06449_),
    .B(_06474_),
    .CIN(_06475_),
    .COUT(_06470_),
    .SUM(_06476_));
 sky130_fd_sc_hd__fa_1 _15137_ (.A(_06477_),
    .B(_06478_),
    .CIN(_06479_),
    .COUT(_06474_),
    .SUM(_06480_));
 sky130_fd_sc_hd__fa_1 _15138_ (.A(_06235_),
    .B(_06481_),
    .CIN(_06482_),
    .COUT(_06483_),
    .SUM(_06484_));
 sky130_fd_sc_hd__fa_1 _15139_ (.A(_06486_),
    .B(_06476_),
    .CIN(_06485_),
    .COUT(_06487_),
    .SUM(_06488_));
 sky130_fd_sc_hd__fa_1 _15140_ (.A(_06489_),
    .B(_06483_),
    .CIN(_06480_),
    .COUT(_06485_),
    .SUM(_06490_));
 sky130_fd_sc_hd__fa_1 _15141_ (.A(_06492_),
    .B(_06493_),
    .CIN(_06494_),
    .COUT(_06491_),
    .SUM(_06495_));
 sky130_fd_sc_hd__fa_1 _15142_ (.A(_06329_),
    .B(_06497_),
    .CIN(_06498_),
    .COUT(_06499_),
    .SUM(_06500_));
 sky130_fd_sc_hd__fa_1 _15143_ (.A(_06501_),
    .B(_06502_),
    .CIN(_06503_),
    .COUT(_06504_),
    .SUM(_06505_));
 sky130_fd_sc_hd__fa_1 _15144_ (.A(_06509_),
    .B(_06508_),
    .CIN(_06490_),
    .COUT(_06510_),
    .SUM(_06511_));
 sky130_fd_sc_hd__fa_1 _15145_ (.A(_06512_),
    .B(_06513_),
    .CIN(_06514_),
    .COUT(_06508_),
    .SUM(_06515_));
 sky130_fd_sc_hd__fa_1 _15146_ (.A(_06515_),
    .B(_06517_),
    .CIN(_06518_),
    .COUT(_06519_),
    .SUM(_06520_));
 sky130_fd_sc_hd__fa_1 _15147_ (.A(_06521_),
    .B(_06522_),
    .CIN(_06523_),
    .COUT(_06524_),
    .SUM(_06525_));
 sky130_fd_sc_hd__fa_1 _15148_ (.A(_06526_),
    .B(_06527_),
    .CIN(_06528_),
    .COUT(_06529_),
    .SUM(_06530_));
 sky130_fd_sc_hd__fa_1 _15149_ (.A(_06531_),
    .B(_06527_),
    .CIN(_06532_),
    .COUT(_06533_),
    .SUM(_06534_));
 sky130_fd_sc_hd__fa_2 _15150_ (.A(_06535_),
    .B(_06537_),
    .CIN(_06536_),
    .COUT(_06538_),
    .SUM(_06539_));
 sky130_fd_sc_hd__fa_1 _15151_ (.A(_06540_),
    .B(_06542_),
    .CIN(_06541_),
    .COUT(_06543_),
    .SUM(_06544_));
 sky130_fd_sc_hd__fa_2 _15152_ (.A(_06545_),
    .B(_06546_),
    .CIN(_06547_),
    .COUT(_06548_),
    .SUM(_06549_));
 sky130_fd_sc_hd__fa_1 _15153_ (.A(_06550_),
    .B(_06551_),
    .CIN(_06552_),
    .COUT(_06553_),
    .SUM(_06554_));
 sky130_fd_sc_hd__fa_1 _15154_ (.A(_06555_),
    .B(_06546_),
    .CIN(_06547_),
    .COUT(_06556_),
    .SUM(_06557_));
 sky130_fd_sc_hd__fa_1 _15155_ (.A(_06558_),
    .B(_06560_),
    .CIN(_06559_),
    .COUT(_06561_),
    .SUM(_06562_));
 sky130_fd_sc_hd__fa_1 _15156_ (.A(_06563_),
    .B(_06564_),
    .CIN(_06565_),
    .COUT(_06542_),
    .SUM(_06566_));
 sky130_fd_sc_hd__fa_1 _15157_ (.A(_06567_),
    .B(_06568_),
    .CIN(_06569_),
    .COUT(_06570_),
    .SUM(_06571_));
 sky130_fd_sc_hd__fa_1 _15158_ (.A(_06572_),
    .B(_06573_),
    .CIN(_06557_),
    .COUT(_06574_),
    .SUM(_06575_));
 sky130_fd_sc_hd__fa_1 _15159_ (.A(_06576_),
    .B(_06577_),
    .CIN(_06551_),
    .COUT(_06578_),
    .SUM(_06579_));
 sky130_fd_sc_hd__fa_1 _15160_ (.A(_06580_),
    .B(_06582_),
    .CIN(_06581_),
    .COUT(_06583_),
    .SUM(_06584_));
 sky130_fd_sc_hd__fa_1 _15161_ (.A(_06586_),
    .B(_06585_),
    .CIN(_06548_),
    .COUT(_06587_),
    .SUM(_06588_));
 sky130_fd_sc_hd__fa_1 _15162_ (.A(_06589_),
    .B(_06584_),
    .CIN(_06590_),
    .COUT(_06591_),
    .SUM(_06592_));
 sky130_fd_sc_hd__fa_1 _15163_ (.A(_06593_),
    .B(_06594_),
    .CIN(_06571_),
    .COUT(_06595_),
    .SUM(_06596_));
 sky130_fd_sc_hd__fa_1 _15164_ (.A(_06597_),
    .B(_06598_),
    .CIN(_06599_),
    .COUT(_06600_),
    .SUM(_06601_));
 sky130_fd_sc_hd__fa_1 _15165_ (.A(_06602_),
    .B(_06549_),
    .CIN(_06603_),
    .COUT(_06604_),
    .SUM(_06605_));
 sky130_fd_sc_hd__fa_1 _15166_ (.A(_06607_),
    .B(_06608_),
    .CIN(_06577_),
    .COUT(_06606_),
    .SUM(_06609_));
 sky130_fd_sc_hd__fa_1 _15167_ (.A(_06551_),
    .B(_06552_),
    .CIN(_06610_),
    .COUT(_06611_),
    .SUM(_06612_));
 sky130_fd_sc_hd__fa_1 _15168_ (.A(_06613_),
    .B(_06614_),
    .CIN(_06605_),
    .COUT(_06615_),
    .SUM(_06616_));
 sky130_fd_sc_hd__fa_1 _15169_ (.A(_06588_),
    .B(_06617_),
    .CIN(_06618_),
    .COUT(_06619_),
    .SUM(_06620_));
 sky130_fd_sc_hd__fa_1 _15170_ (.A(_06621_),
    .B(_06622_),
    .CIN(_06623_),
    .COUT(_06617_),
    .SUM(_06624_));
 sky130_fd_sc_hd__fa_1 _15171_ (.A(_06625_),
    .B(_06627_),
    .CIN(_06626_),
    .COUT(_06628_),
    .SUM(_06629_));
 sky130_fd_sc_hd__fa_1 _15172_ (.A(_06630_),
    .B(net466),
    .CIN(_06632_),
    .COUT(_06633_),
    .SUM(_06634_));
 sky130_fd_sc_hd__fa_1 _15173_ (.A(_06636_),
    .B(_06637_),
    .CIN(_06638_),
    .COUT(_06639_),
    .SUM(_06640_));
 sky130_fd_sc_hd__fa_1 _15174_ (.A(_06641_),
    .B(_06642_),
    .CIN(_06643_),
    .COUT(_06644_),
    .SUM(_06645_));
 sky130_fd_sc_hd__fa_1 _15175_ (.A(net466),
    .B(_06648_),
    .CIN(_06632_),
    .COUT(_06647_),
    .SUM(_06649_));
 sky130_fd_sc_hd__fa_1 _15176_ (.A(_06629_),
    .B(_06650_),
    .CIN(_06592_),
    .COUT(_06651_),
    .SUM(_06652_));
 sky130_fd_sc_hd__fa_1 _15177_ (.A(_06653_),
    .B(_06654_),
    .CIN(_06655_),
    .COUT(_06650_),
    .SUM(_06656_));
 sky130_fd_sc_hd__fa_1 _15178_ (.A(_06657_),
    .B(_06658_),
    .CIN(_06659_),
    .COUT(_06654_),
    .SUM(_06660_));
 sky130_fd_sc_hd__fa_1 _15179_ (.A(_06661_),
    .B(_06662_),
    .CIN(_06565_),
    .COUT(_06663_),
    .SUM(_06664_));
 sky130_fd_sc_hd__fa_1 _15180_ (.A(_06665_),
    .B(_06666_),
    .CIN(_06612_),
    .COUT(_06614_),
    .SUM(_06667_));
 sky130_fd_sc_hd__fa_1 _15181_ (.A(_06563_),
    .B(_06564_),
    .CIN(_06608_),
    .COUT(_06668_),
    .SUM(_06669_));
 sky130_fd_sc_hd__fa_1 _15182_ (.A(_06577_),
    .B(_06551_),
    .CIN(_06552_),
    .COUT(_06670_),
    .SUM(_06671_));
 sky130_fd_sc_hd__fa_1 _15183_ (.A(_06672_),
    .B(_06667_),
    .CIN(_06673_),
    .COUT(_06674_),
    .SUM(_06675_));
 sky130_fd_sc_hd__fa_1 _15184_ (.A(_06624_),
    .B(_06676_),
    .CIN(_06677_),
    .COUT(_06678_),
    .SUM(_06679_));
 sky130_fd_sc_hd__fa_2 _15185_ (.A(_06680_),
    .B(_06681_),
    .CIN(_06682_),
    .COUT(_06676_),
    .SUM(_06683_));
 sky130_fd_sc_hd__fa_1 _15186_ (.A(_06684_),
    .B(_06685_),
    .CIN(_06686_),
    .COUT(_06687_),
    .SUM(_06688_));
 sky130_fd_sc_hd__fa_1 _15187_ (.A(_06640_),
    .B(_06689_),
    .CIN(_06690_),
    .COUT(_06691_),
    .SUM(_06692_));
 sky130_fd_sc_hd__fa_1 _15188_ (.A(_06693_),
    .B(_06649_),
    .CIN(_06694_),
    .COUT(_06695_),
    .SUM(_06696_));
 sky130_fd_sc_hd__fa_1 _15189_ (.A(_06697_),
    .B(_06698_),
    .CIN(_06635_),
    .COUT(_06699_),
    .SUM(_06700_));
 sky130_fd_sc_hd__fa_1 _15190_ (.A(_06687_),
    .B(_06692_),
    .CIN(_06701_),
    .COUT(_06702_),
    .SUM(_06703_));
 sky130_fd_sc_hd__fa_1 _15191_ (.A(_06703_),
    .B(_06704_),
    .CIN(_06652_),
    .COUT(_06705_),
    .SUM(_06706_));
 sky130_fd_sc_hd__fa_2 _15192_ (.A(_06707_),
    .B(_06656_),
    .CIN(_06688_),
    .COUT(_06704_),
    .SUM(_06708_));
 sky130_fd_sc_hd__fa_1 _15193_ (.A(_06709_),
    .B(_06710_),
    .CIN(_06675_),
    .COUT(_06711_),
    .SUM(_06712_));
 sky130_fd_sc_hd__fa_1 _15194_ (.A(_06531_),
    .B(net460),
    .CIN(_06532_),
    .COUT(_06714_),
    .SUM(_06715_));
 sky130_fd_sc_hd__fa_1 _15195_ (.A(_06716_),
    .B(_06717_),
    .CIN(_06671_),
    .COUT(_06673_),
    .SUM(_06718_));
 sky130_fd_sc_hd__fa_1 _15196_ (.A(_06598_),
    .B(_06564_),
    .CIN(_06599_),
    .COUT(_06719_),
    .SUM(_06720_));
 sky130_fd_sc_hd__fa_1 _15197_ (.A(_06537_),
    .B(_06721_),
    .CIN(_06722_),
    .COUT(_06723_),
    .SUM(_06724_));
 sky130_fd_sc_hd__fa_1 _15198_ (.A(_06725_),
    .B(_06718_),
    .CIN(_06726_),
    .COUT(_06727_),
    .SUM(_06728_));
 sky130_fd_sc_hd__fa_1 _15199_ (.A(net491),
    .B(_06683_),
    .CIN(_06730_),
    .COUT(_06731_),
    .SUM(_06732_));
 sky130_fd_sc_hd__fa_1 _15200_ (.A(_06723_),
    .B(_06733_),
    .CIN(_06734_),
    .COUT(_06730_),
    .SUM(_06735_));
 sky130_fd_sc_hd__fa_1 _15201_ (.A(_06736_),
    .B(_06737_),
    .CIN(_06738_),
    .COUT(_06739_),
    .SUM(_06740_));
 sky130_fd_sc_hd__fa_1 _15202_ (.A(_06741_),
    .B(_06742_),
    .CIN(_06743_),
    .COUT(_06701_),
    .SUM(_06744_));
 sky130_fd_sc_hd__fa_1 _15203_ (.A(net466),
    .B(_06745_),
    .CIN(_06746_),
    .COUT(_06747_),
    .SUM(_06748_));
 sky130_fd_sc_hd__fa_1 _15204_ (.A(_06697_),
    .B(_06698_),
    .CIN(_06749_),
    .COUT(_06750_),
    .SUM(_06751_));
 sky130_fd_sc_hd__fa_1 _15205_ (.A(_06739_),
    .B(_06744_),
    .CIN(_06752_),
    .COUT(_06753_),
    .SUM(_06754_));
 sky130_fd_sc_hd__fa_1 _15206_ (.A(_06757_),
    .B(_06755_),
    .CIN(_06756_),
    .COUT(_06758_),
    .SUM(_06759_));
 sky130_fd_sc_hd__fa_1 _15207_ (.A(_06754_),
    .B(_06761_),
    .CIN(_06708_),
    .COUT(_06760_),
    .SUM(_06762_));
 sky130_fd_sc_hd__fa_1 _15208_ (.A(_06763_),
    .B(_06764_),
    .CIN(_06740_),
    .COUT(_06761_),
    .SUM(_06765_));
 sky130_fd_sc_hd__fa_1 _15209_ (.A(_06766_),
    .B(_06767_),
    .CIN(_06728_),
    .COUT(_06768_),
    .SUM(_06769_));
 sky130_fd_sc_hd__fa_1 _15210_ (.A(_06770_),
    .B(_06771_),
    .CIN(_06724_),
    .COUT(_06726_),
    .SUM(_06772_));
 sky130_fd_sc_hd__fa_1 _15211_ (.A(_06662_),
    .B(_06599_),
    .CIN(_06565_),
    .COUT(_06773_),
    .SUM(_06774_));
 sky130_fd_sc_hd__fa_1 _15212_ (.A(_06775_),
    .B(_06537_),
    .CIN(_06721_),
    .COUT(_06776_),
    .SUM(_06777_));
 sky130_fd_sc_hd__fa_1 _15213_ (.A(_06778_),
    .B(_06735_),
    .CIN(_06779_),
    .COUT(_06780_),
    .SUM(_06781_));
 sky130_fd_sc_hd__fa_1 _15214_ (.A(_06776_),
    .B(_06782_),
    .CIN(_06783_),
    .COUT(_06779_),
    .SUM(_06784_));
 sky130_fd_sc_hd__fa_1 _15215_ (.A(_06785_),
    .B(_06781_),
    .CIN(_06786_),
    .COUT(_06787_),
    .SUM(_06788_));
 sky130_fd_sc_hd__fa_1 _15216_ (.A(_06789_),
    .B(_06790_),
    .CIN(_06791_),
    .COUT(_06752_),
    .SUM(_06792_));
 sky130_fd_sc_hd__fa_1 _15217_ (.A(_06632_),
    .B(_06793_),
    .CIN(_06794_),
    .COUT(_06795_),
    .SUM(_06796_));
 sky130_fd_sc_hd__fa_1 _15218_ (.A(_06797_),
    .B(_06697_),
    .CIN(_06749_),
    .COUT(_06798_),
    .SUM(_06799_));
 sky130_fd_sc_hd__fa_1 _15219_ (.A(_06800_),
    .B(_06792_),
    .CIN(_06801_),
    .COUT(_06802_),
    .SUM(_06803_));
 sky130_fd_sc_hd__fa_2 _15220_ (.A(_06805_),
    .B(_06759_),
    .CIN(_06804_),
    .COUT(_06806_),
    .SUM(_06807_));
 sky130_fd_sc_hd__fa_1 _15221_ (.A(_06810_),
    .B(_06809_),
    .CIN(_06808_),
    .COUT(_06804_),
    .SUM(_06811_));
 sky130_fd_sc_hd__fa_1 _15222_ (.A(_06765_),
    .B(_06813_),
    .CIN(_06803_),
    .COUT(_06812_),
    .SUM(_06814_));
 sky130_fd_sc_hd__fa_1 _15223_ (.A(_06815_),
    .B(_06816_),
    .CIN(_06817_),
    .COUT(_06813_),
    .SUM(_06818_));
 sky130_fd_sc_hd__fa_1 _15224_ (.A(_06819_),
    .B(_06820_),
    .CIN(_06821_),
    .COUT(_06822_),
    .SUM(_06823_));
 sky130_fd_sc_hd__fa_1 _15225_ (.A(_06824_),
    .B(_06825_),
    .CIN(_06777_),
    .COUT(_06826_),
    .SUM(_06827_));
 sky130_fd_sc_hd__fa_1 _15226_ (.A(_06829_),
    .B(_06597_),
    .CIN(_06565_),
    .COUT(_06828_),
    .SUM(_06830_));
 sky130_fd_sc_hd__fa_1 _15227_ (.A(_06564_),
    .B(_06599_),
    .CIN(_06608_),
    .COUT(_06831_),
    .SUM(_06832_));
 sky130_fd_sc_hd__fa_1 _15228_ (.A(_06833_),
    .B(_06784_),
    .CIN(_06834_),
    .COUT(_06786_),
    .SUM(_06835_));
 sky130_fd_sc_hd__fa_1 _15229_ (.A(_06836_),
    .B(_06837_),
    .CIN(_06838_),
    .COUT(_06834_),
    .SUM(_06839_));
 sky130_fd_sc_hd__fa_1 _15230_ (.A(_06840_),
    .B(_06841_),
    .CIN(_06842_),
    .COUT(_06843_),
    .SUM(_06844_));
 sky130_fd_sc_hd__fa_1 _15231_ (.A(_06845_),
    .B(_06846_),
    .CIN(_06847_),
    .COUT(_06801_),
    .SUM(_06848_));
 sky130_fd_sc_hd__fa_1 _15232_ (.A(_06648_),
    .B(_06849_),
    .CIN(_06850_),
    .COUT(_06851_),
    .SUM(_06852_));
 sky130_fd_sc_hd__fa_1 _15233_ (.A(_06853_),
    .B(_06797_),
    .CIN(_06749_),
    .COUT(_06854_),
    .SUM(_06855_));
 sky130_fd_sc_hd__fa_1 _15234_ (.A(_06856_),
    .B(_06857_),
    .CIN(_06858_),
    .COUT(_06859_),
    .SUM(_06860_));
 sky130_fd_sc_hd__fa_1 _15235_ (.A(_06811_),
    .B(_06861_),
    .CIN(_06862_),
    .COUT(_06863_),
    .SUM(_06864_));
 sky130_fd_sc_hd__fa_1 _15236_ (.A(_06865_),
    .B(_06866_),
    .CIN(_06867_),
    .COUT(_06861_),
    .SUM(_06868_));
 sky130_fd_sc_hd__fa_1 _15237_ (.A(_06818_),
    .B(_06870_),
    .CIN(_06871_),
    .COUT(_06869_),
    .SUM(_06872_));
 sky130_fd_sc_hd__fa_1 _15238_ (.A(_06873_),
    .B(_06874_),
    .CIN(_06844_),
    .COUT(_06870_),
    .SUM(_06875_));
 sky130_fd_sc_hd__fa_1 _15239_ (.A(_06876_),
    .B(_06877_),
    .CIN(_06878_),
    .COUT(_06874_),
    .SUM(_06879_));
 sky130_fd_sc_hd__fa_1 _15240_ (.A(_06880_),
    .B(_06881_),
    .CIN(_06882_),
    .COUT(_06883_),
    .SUM(_06884_));
 sky130_fd_sc_hd__fa_1 _15241_ (.A(_06661_),
    .B(_06597_),
    .CIN(_06886_),
    .COUT(_06885_),
    .SUM(_06887_));
 sky130_fd_sc_hd__fa_1 _15242_ (.A(_06564_),
    .B(_06599_),
    .CIN(_06565_),
    .COUT(_06888_),
    .SUM(_06889_));
 sky130_fd_sc_hd__fa_1 _15243_ (.A(_06890_),
    .B(_06891_),
    .CIN(_06892_),
    .COUT(_06893_),
    .SUM(_06894_));
 sky130_fd_sc_hd__fa_1 _15244_ (.A(_06895_),
    .B(_06896_),
    .CIN(_06897_),
    .COUT(_06898_),
    .SUM(_06899_));
 sky130_fd_sc_hd__fa_1 _15245_ (.A(_06697_),
    .B(_06855_),
    .CIN(_06900_),
    .COUT(_06901_),
    .SUM(_06902_));
 sky130_fd_sc_hd__fa_1 _15246_ (.A(_06853_),
    .B(_06903_),
    .CIN(_06797_),
    .COUT(_06900_),
    .SUM(_06904_));
 sky130_fd_sc_hd__fa_1 _15247_ (.A(_06905_),
    .B(_06906_),
    .CIN(_06907_),
    .COUT(_06908_),
    .SUM(_06909_));
 sky130_fd_sc_hd__fa_1 _15248_ (.A(_06868_),
    .B(_06910_),
    .CIN(_06911_),
    .COUT(_06912_),
    .SUM(_06913_));
 sky130_fd_sc_hd__fa_1 _15249_ (.A(_06914_),
    .B(_06915_),
    .CIN(_06916_),
    .COUT(_06910_),
    .SUM(_06917_));
 sky130_fd_sc_hd__fa_1 _15250_ (.A(_06875_),
    .B(_06919_),
    .CIN(_06920_),
    .COUT(_06918_),
    .SUM(_06921_));
 sky130_fd_sc_hd__fa_1 _15251_ (.A(_06922_),
    .B(_06923_),
    .CIN(_06924_),
    .COUT(_06925_),
    .SUM(_06926_));
 sky130_fd_sc_hd__fa_1 _15252_ (.A(_06887_),
    .B(_06927_),
    .CIN(_06889_),
    .COUT(_06928_),
    .SUM(_06929_));
 sky130_fd_sc_hd__fa_1 _15253_ (.A(_06597_),
    .B(_06599_),
    .CIN(_06565_),
    .COUT(_06931_),
    .SUM(_06932_));
 sky130_fd_sc_hd__fa_1 _15254_ (.A(_06933_),
    .B(_06934_),
    .CIN(_06935_),
    .COUT(_06936_),
    .SUM(_06937_));
 sky130_fd_sc_hd__fa_1 _15255_ (.A(_06938_),
    .B(_06939_),
    .CIN(_06940_),
    .COUT(_06941_),
    .SUM(_06942_));
 sky130_fd_sc_hd__fa_1 _15256_ (.A(_06943_),
    .B(_06944_),
    .CIN(_06945_),
    .COUT(_06946_),
    .SUM(_06947_));
 sky130_fd_sc_hd__fa_1 _15257_ (.A(_06948_),
    .B(_06853_),
    .CIN(_06903_),
    .COUT(_06949_),
    .SUM(_06950_));
 sky130_fd_sc_hd__fa_1 _15258_ (.A(_06951_),
    .B(_06952_),
    .CIN(_06953_),
    .COUT(_06954_),
    .SUM(_06955_));
 sky130_fd_sc_hd__fa_1 _15259_ (.A(_06917_),
    .B(_06956_),
    .CIN(_06957_),
    .COUT(_06958_),
    .SUM(_06959_));
 sky130_fd_sc_hd__fa_1 _15260_ (.A(_06960_),
    .B(_06961_),
    .CIN(_06962_),
    .COUT(_06956_),
    .SUM(_06963_));
 sky130_fd_sc_hd__fa_1 _15261_ (.A(_06965_),
    .B(_06966_),
    .CIN(_06967_),
    .COUT(_06964_),
    .SUM(_06968_));
 sky130_fd_sc_hd__fa_1 _15262_ (.A(_06969_),
    .B(_06970_),
    .CIN(_06971_),
    .COUT(_06972_),
    .SUM(_06973_));
 sky130_fd_sc_hd__fa_1 _15263_ (.A(_06597_),
    .B(_06661_),
    .CIN(_06565_),
    .COUT(_06974_),
    .SUM(_06975_));
 sky130_fd_sc_hd__fa_1 _15264_ (.A(_06976_),
    .B(_06977_),
    .CIN(_06978_),
    .COUT(_06979_),
    .SUM(_06980_));
 sky130_fd_sc_hd__fa_1 _15265_ (.A(_06981_),
    .B(_06982_),
    .CIN(_06983_),
    .COUT(_06984_),
    .SUM(_06985_));
 sky130_fd_sc_hd__fa_1 _15266_ (.A(_06986_),
    .B(_06987_),
    .CIN(_06988_),
    .COUT(_06989_),
    .SUM(_06990_));
 sky130_fd_sc_hd__fa_1 _15267_ (.A(net488),
    .B(_06778_),
    .CIN(_06991_),
    .COUT(_06988_),
    .SUM(_06992_));
 sky130_fd_sc_hd__fa_1 _15268_ (.A(_06993_),
    .B(_06994_),
    .CIN(_06995_),
    .COUT(_06996_),
    .SUM(_06997_));
 sky130_fd_sc_hd__fa_1 _15269_ (.A(_06963_),
    .B(_06998_),
    .CIN(_06999_),
    .COUT(_07000_),
    .SUM(_07001_));
 sky130_fd_sc_hd__fa_1 _15270_ (.A(_07004_),
    .B(_07003_),
    .CIN(_07002_),
    .COUT(_06998_),
    .SUM(_07005_));
 sky130_fd_sc_hd__fa_1 _15271_ (.A(_07007_),
    .B(_07008_),
    .CIN(_07009_),
    .COUT(_07006_),
    .SUM(_07010_));
 sky130_fd_sc_hd__fa_1 _15272_ (.A(_07011_),
    .B(_07012_),
    .CIN(_07013_),
    .COUT(_07014_),
    .SUM(_07015_));
 sky130_fd_sc_hd__fa_1 _15273_ (.A(_07016_),
    .B(_07017_),
    .CIN(_07018_),
    .COUT(_07019_),
    .SUM(_07020_));
 sky130_fd_sc_hd__fa_1 _15274_ (.A(_06853_),
    .B(_07021_),
    .CIN(_07022_),
    .COUT(_07023_),
    .SUM(_07024_));
 sky130_fd_sc_hd__fa_1 _15275_ (.A(net488),
    .B(_06778_),
    .CIN(_06833_),
    .COUT(_07025_),
    .SUM(_07026_));
 sky130_fd_sc_hd__fa_1 _15276_ (.A(_07027_),
    .B(_07028_),
    .CIN(_07029_),
    .COUT(_07030_),
    .SUM(_07031_));
 sky130_fd_sc_hd__fa_1 _15277_ (.A(_07005_),
    .B(_07032_),
    .CIN(_07033_),
    .COUT(_07034_),
    .SUM(_07035_));
 sky130_fd_sc_hd__fa_1 _15278_ (.A(_07038_),
    .B(_07037_),
    .CIN(_07036_),
    .COUT(_07032_),
    .SUM(_07039_));
 sky130_fd_sc_hd__fa_1 _15279_ (.A(_07015_),
    .B(_07040_),
    .CIN(_07041_),
    .COUT(_07037_),
    .SUM(_07042_));
 sky130_fd_sc_hd__fa_1 _15280_ (.A(_07043_),
    .B(_07044_),
    .CIN(_07045_),
    .COUT(_07040_),
    .SUM(_07046_));
 sky130_fd_sc_hd__fa_1 _15281_ (.A(net459),
    .B(_06526_),
    .CIN(_06532_),
    .COUT(_07016_),
    .SUM(_07047_));
 sky130_fd_sc_hd__fa_1 _15282_ (.A(_06927_),
    .B(_07048_),
    .CIN(_07049_),
    .COUT(_07050_),
    .SUM(_07051_));
 sky130_fd_sc_hd__fa_1 _15283_ (.A(_07039_),
    .B(_07052_),
    .CIN(_07053_),
    .COUT(_07054_),
    .SUM(_07055_));
 sky130_fd_sc_hd__fa_1 _15284_ (.A(_07042_),
    .B(_07056_),
    .CIN(_07057_),
    .COUT(_07052_),
    .SUM(_07058_));
 sky130_fd_sc_hd__fa_1 _15285_ (.A(_07046_),
    .B(_07059_),
    .CIN(_07060_),
    .COUT(_07056_),
    .SUM(_07061_));
 sky130_fd_sc_hd__fa_1 _15286_ (.A(_07062_),
    .B(_07063_),
    .CIN(_07064_),
    .COUT(_07059_),
    .SUM(_07065_));
 sky130_fd_sc_hd__fa_1 _15287_ (.A(_06991_),
    .B(_07066_),
    .CIN(_07026_),
    .COUT(_07067_),
    .SUM(_07068_));
 sky130_fd_sc_hd__fa_1 _15288_ (.A(_07069_),
    .B(_07070_),
    .CIN(_07071_),
    .COUT(_07072_),
    .SUM(_07073_));
 sky130_fd_sc_hd__fa_1 _15289_ (.A(_07058_),
    .B(_07074_),
    .CIN(_07075_),
    .COUT(_07076_),
    .SUM(_07077_));
 sky130_fd_sc_hd__fa_1 _15290_ (.A(_07061_),
    .B(_07078_),
    .CIN(_07079_),
    .COUT(_07074_),
    .SUM(_07080_));
 sky130_fd_sc_hd__fa_1 _15291_ (.A(_07065_),
    .B(_07081_),
    .CIN(_07082_),
    .COUT(_07078_),
    .SUM(_07083_));
 sky130_fd_sc_hd__fa_1 _15292_ (.A(_07084_),
    .B(_07085_),
    .CIN(_07086_),
    .COUT(_07081_),
    .SUM(_07087_));
 sky130_fd_sc_hd__fa_1 _15293_ (.A(_07088_),
    .B(_07083_),
    .CIN(_07089_),
    .COUT(_07090_),
    .SUM(_07091_));
 sky130_fd_sc_hd__fa_1 _15294_ (.A(_07087_),
    .B(_07092_),
    .CIN(_07093_),
    .COUT(_07089_),
    .SUM(_07094_));
 sky130_fd_sc_hd__fa_1 _15295_ (.A(_07096_),
    .B(_07097_),
    .CIN(_07098_),
    .COUT(_07095_),
    .SUM(_07099_));
 sky130_fd_sc_hd__fa_1 _15296_ (.A(_07099_),
    .B(_07100_),
    .CIN(_07101_),
    .COUT(_07102_),
    .SUM(_07103_));
 sky130_fd_sc_hd__ha_4 _15297_ (.A(net385),
    .B(_07106_),
    .COUT(_07107_),
    .SUM(_07108_));
 sky130_fd_sc_hd__ha_4 _15298_ (.A(_05892_),
    .B(_07109_),
    .COUT(_07110_),
    .SUM(_07111_));
 sky130_fd_sc_hd__ha_4 _15299_ (.A(_07113_),
    .B(_07112_),
    .COUT(_07114_),
    .SUM(_07115_));
 sky130_fd_sc_hd__ha_1 _15300_ (.A(_05892_),
    .B(_07116_),
    .COUT(_07117_),
    .SUM(_07118_));
 sky130_fd_sc_hd__ha_1 _15301_ (.A(_07106_),
    .B(net358),
    .COUT(_07119_),
    .SUM(_07120_));
 sky130_fd_sc_hd__ha_4 _15302_ (.A(_07121_),
    .B(_07122_),
    .COUT(_07123_),
    .SUM(_07124_));
 sky130_fd_sc_hd__ha_1 _15303_ (.A(_07112_),
    .B(_07125_),
    .COUT(_07126_),
    .SUM(_07127_));
 sky130_fd_sc_hd__ha_1 _15304_ (.A(_05892_),
    .B(_07128_),
    .COUT(_07129_),
    .SUM(_07130_));
 sky130_fd_sc_hd__ha_1 _15305_ (.A(_07106_),
    .B(net359),
    .COUT(_07131_),
    .SUM(_07132_));
 sky130_fd_sc_hd__ha_1 _15306_ (.A(_07133_),
    .B(_07134_),
    .COUT(_07135_),
    .SUM(_07136_));
 sky130_fd_sc_hd__ha_1 _15307_ (.A(_07121_),
    .B(_07137_),
    .COUT(_07138_),
    .SUM(_07139_));
 sky130_fd_sc_hd__ha_4 _15308_ (.A(_07112_),
    .B(_07140_),
    .COUT(_07141_),
    .SUM(_07142_));
 sky130_fd_sc_hd__ha_1 _15309_ (.A(_05892_),
    .B(_07143_),
    .COUT(_07144_),
    .SUM(_07145_));
 sky130_fd_sc_hd__ha_1 _15310_ (.A(_07106_),
    .B(net360),
    .COUT(_07146_),
    .SUM(_07147_));
 sky130_fd_sc_hd__ha_2 _15311_ (.A(_05892_),
    .B(_07148_),
    .COUT(_07149_),
    .SUM(_07150_));
 sky130_fd_sc_hd__ha_1 _15312_ (.A(_07106_),
    .B(net361),
    .COUT(_07151_),
    .SUM(_07152_));
 sky130_fd_sc_hd__ha_2 _15313_ (.A(_07154_),
    .B(_07153_),
    .COUT(_07155_),
    .SUM(_07156_));
 sky130_fd_sc_hd__ha_4 _15314_ (.A(_07133_),
    .B(_07157_),
    .COUT(_07158_),
    .SUM(_07159_));
 sky130_fd_sc_hd__ha_2 _15315_ (.A(_07121_),
    .B(_07160_),
    .COUT(_07161_),
    .SUM(_07162_));
 sky130_fd_sc_hd__ha_4 _15316_ (.A(_07163_),
    .B(_07112_),
    .COUT(_07164_),
    .SUM(_07165_));
 sky130_fd_sc_hd__ha_2 _15317_ (.A(_07167_),
    .B(_07166_),
    .COUT(_07168_),
    .SUM(_07169_));
 sky130_fd_sc_hd__ha_1 _15318_ (.A(_07153_),
    .B(_07170_),
    .COUT(_07171_),
    .SUM(_07172_));
 sky130_fd_sc_hd__ha_4 _15319_ (.A(_07173_),
    .B(_07133_),
    .COUT(_07174_),
    .SUM(_07175_));
 sky130_fd_sc_hd__ha_2 _15320_ (.A(_07121_),
    .B(_07176_),
    .COUT(_07177_),
    .SUM(_07178_));
 sky130_fd_sc_hd__ha_2 _15321_ (.A(_07112_),
    .B(_07179_),
    .COUT(_07180_),
    .SUM(_07181_));
 sky130_fd_sc_hd__ha_1 _15322_ (.A(_05892_),
    .B(_07182_),
    .COUT(_07183_),
    .SUM(_07184_));
 sky130_fd_sc_hd__ha_2 _15323_ (.A(_07106_),
    .B(net362),
    .COUT(_07185_),
    .SUM(_07186_));
 sky130_fd_sc_hd__ha_1 _15324_ (.A(_07166_),
    .B(_07187_),
    .COUT(_07188_),
    .SUM(_07189_));
 sky130_fd_sc_hd__ha_2 _15325_ (.A(_07153_),
    .B(_07190_),
    .COUT(_07191_),
    .SUM(_07192_));
 sky130_fd_sc_hd__ha_4 _15326_ (.A(_07193_),
    .B(_07133_),
    .COUT(_07194_),
    .SUM(_07195_));
 sky130_fd_sc_hd__ha_4 _15327_ (.A(_07196_),
    .B(_07121_),
    .COUT(_07197_),
    .SUM(_07198_));
 sky130_fd_sc_hd__ha_1 _15328_ (.A(_07112_),
    .B(_07199_),
    .COUT(_07200_),
    .SUM(_07201_));
 sky130_fd_sc_hd__ha_1 _15329_ (.A(_05892_),
    .B(_07202_),
    .COUT(_07203_),
    .SUM(_07204_));
 sky130_fd_sc_hd__ha_2 _15330_ (.A(_07106_),
    .B(net363),
    .COUT(_07205_),
    .SUM(_07206_));
 sky130_fd_sc_hd__ha_1 _15331_ (.A(_07207_),
    .B(_07208_),
    .COUT(_07209_),
    .SUM(_07210_));
 sky130_fd_sc_hd__ha_1 _15332_ (.A(_07166_),
    .B(_07211_),
    .COUT(_07212_),
    .SUM(_07213_));
 sky130_fd_sc_hd__ha_1 _15333_ (.A(_07153_),
    .B(_07214_),
    .COUT(_07215_),
    .SUM(_07216_));
 sky130_fd_sc_hd__ha_4 _15334_ (.A(_07217_),
    .B(_07133_),
    .COUT(_07218_),
    .SUM(_07219_));
 sky130_fd_sc_hd__ha_1 _15335_ (.A(_07121_),
    .B(_07220_),
    .COUT(_07221_),
    .SUM(_07222_));
 sky130_fd_sc_hd__ha_1 _15336_ (.A(_07112_),
    .B(_07223_),
    .COUT(_07224_),
    .SUM(_07225_));
 sky130_fd_sc_hd__ha_1 _15337_ (.A(_05892_),
    .B(_07226_),
    .COUT(_07227_),
    .SUM(_07228_));
 sky130_fd_sc_hd__ha_1 _15338_ (.A(net24),
    .B(net364),
    .COUT(_07229_),
    .SUM(_07230_));
 sky130_fd_sc_hd__ha_2 _15339_ (.A(_07166_),
    .B(_07231_),
    .COUT(_07232_),
    .SUM(_07233_));
 sky130_fd_sc_hd__ha_4 _15340_ (.A(_07153_),
    .B(_07234_),
    .COUT(_07235_),
    .SUM(_07236_));
 sky130_fd_sc_hd__ha_1 _15341_ (.A(_07133_),
    .B(_07237_),
    .COUT(_07238_),
    .SUM(_07239_));
 sky130_fd_sc_hd__ha_4 _15342_ (.A(_07121_),
    .B(_07240_),
    .COUT(_07241_),
    .SUM(_07242_));
 sky130_fd_sc_hd__ha_4 _15343_ (.A(_07112_),
    .B(_07243_),
    .COUT(_07244_),
    .SUM(_07245_));
 sky130_fd_sc_hd__ha_4 _15344_ (.A(_07246_),
    .B(_05892_),
    .COUT(_07247_),
    .SUM(_07248_));
 sky130_fd_sc_hd__ha_1 _15345_ (.A(net24),
    .B(net365),
    .COUT(_07249_),
    .SUM(_07250_));
 sky130_fd_sc_hd__ha_2 _15346_ (.A(_07166_),
    .B(_07251_),
    .COUT(_07252_),
    .SUM(_07253_));
 sky130_fd_sc_hd__ha_4 _15347_ (.A(_07254_),
    .B(_07153_),
    .COUT(_07255_),
    .SUM(_07256_));
 sky130_fd_sc_hd__ha_4 _15348_ (.A(_07257_),
    .B(_07133_),
    .COUT(_07258_),
    .SUM(_07259_));
 sky130_fd_sc_hd__ha_1 _15349_ (.A(_07112_),
    .B(_07260_),
    .COUT(_07261_),
    .SUM(_07262_));
 sky130_fd_sc_hd__ha_1 _15350_ (.A(_05892_),
    .B(_07263_),
    .COUT(_07264_),
    .SUM(_07265_));
 sky130_fd_sc_hd__ha_1 _15351_ (.A(net24),
    .B(net366),
    .COUT(_07266_),
    .SUM(_07267_));
 sky130_fd_sc_hd__ha_4 _15352_ (.A(_07121_),
    .B(_07268_),
    .COUT(_07269_),
    .SUM(_07270_));
 sky130_fd_sc_hd__ha_2 _15353_ (.A(_07166_),
    .B(_07271_),
    .COUT(_07272_),
    .SUM(_07273_));
 sky130_fd_sc_hd__ha_1 _15354_ (.A(_07153_),
    .B(_07274_),
    .COUT(_07275_),
    .SUM(_07276_));
 sky130_fd_sc_hd__ha_1 _15355_ (.A(_07133_),
    .B(_07277_),
    .COUT(_07278_),
    .SUM(_07279_));
 sky130_fd_sc_hd__ha_1 _15356_ (.A(_07121_),
    .B(_07280_),
    .COUT(_07281_),
    .SUM(_07282_));
 sky130_fd_sc_hd__ha_1 _15357_ (.A(_07283_),
    .B(_07112_),
    .COUT(_07284_),
    .SUM(_07285_));
 sky130_fd_sc_hd__ha_4 _15358_ (.A(_05892_),
    .B(_07286_),
    .COUT(_07287_),
    .SUM(_07288_));
 sky130_fd_sc_hd__ha_1 _15359_ (.A(net24),
    .B(net367),
    .COUT(_07289_),
    .SUM(_07290_));
 sky130_fd_sc_hd__ha_1 _15360_ (.A(_07112_),
    .B(_07291_),
    .COUT(_07292_),
    .SUM(_07293_));
 sky130_fd_sc_hd__ha_1 _15361_ (.A(_05892_),
    .B(_07294_),
    .COUT(_07295_),
    .SUM(_07296_));
 sky130_fd_sc_hd__ha_1 _15362_ (.A(_07133_),
    .B(_07297_),
    .COUT(_07298_),
    .SUM(_07299_));
 sky130_fd_sc_hd__ha_1 _15363_ (.A(_07121_),
    .B(_07300_),
    .COUT(_07301_),
    .SUM(_07302_));
 sky130_fd_sc_hd__ha_1 _15364_ (.A(net24),
    .B(net368),
    .COUT(_07303_),
    .SUM(_07304_));
 sky130_fd_sc_hd__ha_2 _15365_ (.A(_07166_),
    .B(_07305_),
    .COUT(_07306_),
    .SUM(_07307_));
 sky130_fd_sc_hd__ha_1 _15366_ (.A(_07153_),
    .B(_07308_),
    .COUT(_07309_),
    .SUM(_07310_));
 sky130_fd_sc_hd__ha_1 _15367_ (.A(_07166_),
    .B(_07311_),
    .COUT(_07312_),
    .SUM(_07313_));
 sky130_fd_sc_hd__ha_1 _15368_ (.A(_07153_),
    .B(_07314_),
    .COUT(_07315_),
    .SUM(_07316_));
 sky130_fd_sc_hd__ha_1 _15369_ (.A(_07133_),
    .B(_07317_),
    .COUT(_07318_),
    .SUM(_07319_));
 sky130_fd_sc_hd__ha_1 _15370_ (.A(_07121_),
    .B(_07320_),
    .COUT(_07321_),
    .SUM(_07322_));
 sky130_fd_sc_hd__ha_4 _15371_ (.A(_07112_),
    .B(_07323_),
    .COUT(_07324_),
    .SUM(_07325_));
 sky130_fd_sc_hd__ha_4 _15372_ (.A(_05892_),
    .B(_07326_),
    .COUT(_07327_),
    .SUM(_07328_));
 sky130_fd_sc_hd__ha_1 _15373_ (.A(net24),
    .B(net369),
    .COUT(_07329_),
    .SUM(_07330_));
 sky130_fd_sc_hd__ha_1 _15374_ (.A(_07166_),
    .B(_07331_),
    .COUT(_07332_),
    .SUM(_07333_));
 sky130_fd_sc_hd__ha_1 _15375_ (.A(_07153_),
    .B(_07334_),
    .COUT(_07335_),
    .SUM(_07336_));
 sky130_fd_sc_hd__ha_1 _15376_ (.A(_07133_),
    .B(_07337_),
    .COUT(_07338_),
    .SUM(_07339_));
 sky130_fd_sc_hd__ha_1 _15377_ (.A(_07121_),
    .B(_07340_),
    .COUT(_07341_),
    .SUM(_07342_));
 sky130_fd_sc_hd__ha_1 _15378_ (.A(_07112_),
    .B(_07343_),
    .COUT(_07344_),
    .SUM(_07345_));
 sky130_fd_sc_hd__ha_4 _15379_ (.A(_07346_),
    .B(_05892_),
    .COUT(_07347_),
    .SUM(_07348_));
 sky130_fd_sc_hd__ha_1 _15380_ (.A(net24),
    .B(net370),
    .COUT(_07349_),
    .SUM(_07350_));
 sky130_fd_sc_hd__ha_2 _15381_ (.A(_07166_),
    .B(_07351_),
    .COUT(_07352_),
    .SUM(_07353_));
 sky130_fd_sc_hd__ha_1 _15382_ (.A(_07153_),
    .B(_07354_),
    .COUT(_07355_),
    .SUM(_07356_));
 sky130_fd_sc_hd__ha_1 _15383_ (.A(_07133_),
    .B(_07357_),
    .COUT(_07358_),
    .SUM(_07359_));
 sky130_fd_sc_hd__ha_1 _15384_ (.A(_07121_),
    .B(_07360_),
    .COUT(_07361_),
    .SUM(_07362_));
 sky130_fd_sc_hd__ha_1 _15385_ (.A(_07363_),
    .B(_07112_),
    .COUT(_07364_),
    .SUM(_07365_));
 sky130_fd_sc_hd__ha_4 _15386_ (.A(_05892_),
    .B(_07366_),
    .COUT(_07367_),
    .SUM(_07368_));
 sky130_fd_sc_hd__ha_1 _15387_ (.A(net24),
    .B(net371),
    .COUT(_07369_),
    .SUM(_07370_));
 sky130_fd_sc_hd__ha_1 _15388_ (.A(net14),
    .B(net372),
    .COUT(_07371_),
    .SUM(_07372_));
 sky130_fd_sc_hd__ha_1 _15389_ (.A(_07166_),
    .B(_07373_),
    .COUT(_07374_),
    .SUM(_07375_));
 sky130_fd_sc_hd__ha_1 _15390_ (.A(_07153_),
    .B(_07376_),
    .COUT(_07377_),
    .SUM(_07378_));
 sky130_fd_sc_hd__ha_1 _15391_ (.A(_07133_),
    .B(_07379_),
    .COUT(_07380_),
    .SUM(_07381_));
 sky130_fd_sc_hd__ha_1 _15392_ (.A(_07121_),
    .B(_07382_),
    .COUT(_07383_),
    .SUM(_07384_));
 sky130_fd_sc_hd__ha_1 _15393_ (.A(_07385_),
    .B(_07112_),
    .COUT(_07386_),
    .SUM(_07387_));
 sky130_fd_sc_hd__ha_4 _15394_ (.A(_05892_),
    .B(_07388_),
    .COUT(_07389_),
    .SUM(_07390_));
 sky130_fd_sc_hd__ha_4 _15395_ (.A(_05892_),
    .B(_07391_),
    .COUT(_07392_),
    .SUM(_07393_));
 sky130_fd_sc_hd__ha_1 _15396_ (.A(net14),
    .B(net373),
    .COUT(_07394_),
    .SUM(_07395_));
 sky130_fd_sc_hd__ha_2 _15397_ (.A(_07166_),
    .B(_07396_),
    .COUT(_07397_),
    .SUM(_07398_));
 sky130_fd_sc_hd__ha_1 _15398_ (.A(_07153_),
    .B(_07399_),
    .COUT(_07400_),
    .SUM(_07401_));
 sky130_fd_sc_hd__ha_1 _15399_ (.A(_07133_),
    .B(_07402_),
    .COUT(_07403_),
    .SUM(_07404_));
 sky130_fd_sc_hd__ha_4 _15400_ (.A(_07121_),
    .B(_07405_),
    .COUT(_07406_),
    .SUM(_07407_));
 sky130_fd_sc_hd__ha_1 _15401_ (.A(_07112_),
    .B(_07408_),
    .COUT(_07409_),
    .SUM(_07410_));
 sky130_fd_sc_hd__ha_4 _15402_ (.A(_07112_),
    .B(_07411_),
    .COUT(_07412_),
    .SUM(_07413_));
 sky130_fd_sc_hd__ha_4 _15403_ (.A(_05892_),
    .B(_07414_),
    .COUT(_07415_),
    .SUM(_07416_));
 sky130_fd_sc_hd__ha_1 _15404_ (.A(net14),
    .B(net374),
    .COUT(_07417_),
    .SUM(_07418_));
 sky130_fd_sc_hd__ha_1 _15405_ (.A(_07166_),
    .B(_07419_),
    .COUT(_07420_),
    .SUM(_07421_));
 sky130_fd_sc_hd__ha_1 _15406_ (.A(_07153_),
    .B(_07422_),
    .COUT(_07423_),
    .SUM(_07424_));
 sky130_fd_sc_hd__ha_1 _15407_ (.A(_07133_),
    .B(_07425_),
    .COUT(_07426_),
    .SUM(_07427_));
 sky130_fd_sc_hd__ha_1 _15408_ (.A(_07121_),
    .B(_07428_),
    .COUT(_07429_),
    .SUM(_07430_));
 sky130_fd_sc_hd__ha_1 _15409_ (.A(_07121_),
    .B(_07431_),
    .COUT(_07432_),
    .SUM(_07433_));
 sky130_fd_sc_hd__ha_4 _15410_ (.A(_07112_),
    .B(_07434_),
    .COUT(_07435_),
    .SUM(_07436_));
 sky130_fd_sc_hd__ha_4 _15411_ (.A(_07437_),
    .B(_05892_),
    .COUT(_07438_),
    .SUM(_07439_));
 sky130_fd_sc_hd__ha_1 _15412_ (.A(net14),
    .B(net375),
    .COUT(_07440_),
    .SUM(_07441_));
 sky130_fd_sc_hd__ha_2 _15413_ (.A(_07166_),
    .B(_07442_),
    .COUT(_07443_),
    .SUM(_07444_));
 sky130_fd_sc_hd__ha_1 _15414_ (.A(_07153_),
    .B(_07445_),
    .COUT(_07446_),
    .SUM(_07447_));
 sky130_fd_sc_hd__ha_1 _15415_ (.A(_07133_),
    .B(_07448_),
    .COUT(_07449_),
    .SUM(_07450_));
 sky130_fd_sc_hd__ha_1 _15416_ (.A(_07133_),
    .B(_07451_),
    .COUT(_07452_),
    .SUM(_07453_));
 sky130_fd_sc_hd__ha_1 _15417_ (.A(_07121_),
    .B(_07454_),
    .COUT(_07455_),
    .SUM(_07456_));
 sky130_fd_sc_hd__ha_4 _15418_ (.A(_07112_),
    .B(_07457_),
    .COUT(_07458_),
    .SUM(_07459_));
 sky130_fd_sc_hd__ha_4 _15419_ (.A(_05892_),
    .B(_07460_),
    .COUT(_07461_),
    .SUM(_07462_));
 sky130_fd_sc_hd__ha_1 _15420_ (.A(net14),
    .B(net376),
    .COUT(_07463_),
    .SUM(_07464_));
 sky130_fd_sc_hd__ha_2 _15421_ (.A(_07166_),
    .B(_07465_),
    .COUT(_07466_),
    .SUM(_07467_));
 sky130_fd_sc_hd__ha_1 _15422_ (.A(_07153_),
    .B(_07468_),
    .COUT(_07469_),
    .SUM(_07470_));
 sky130_fd_sc_hd__ha_1 _15423_ (.A(_07153_),
    .B(_07471_),
    .COUT(_07472_),
    .SUM(_07473_));
 sky130_fd_sc_hd__ha_1 _15424_ (.A(_07133_),
    .B(_07474_),
    .COUT(_07475_),
    .SUM(_07476_));
 sky130_fd_sc_hd__ha_1 _15425_ (.A(_07121_),
    .B(_07477_),
    .COUT(_07478_),
    .SUM(_07479_));
 sky130_fd_sc_hd__ha_4 _15426_ (.A(_07112_),
    .B(_07480_),
    .COUT(_07481_),
    .SUM(_07482_));
 sky130_fd_sc_hd__ha_1 _15427_ (.A(_05892_),
    .B(_07483_),
    .COUT(_07484_),
    .SUM(_07485_));
 sky130_fd_sc_hd__ha_1 _15428_ (.A(net14),
    .B(net377),
    .COUT(_07486_),
    .SUM(_07487_));
 sky130_fd_sc_hd__ha_1 _15429_ (.A(_07166_),
    .B(_07488_),
    .COUT(_07489_),
    .SUM(_07490_));
 sky130_fd_sc_hd__ha_1 _15430_ (.A(_07166_),
    .B(_07491_),
    .COUT(_07492_),
    .SUM(_07493_));
 sky130_fd_sc_hd__ha_1 _15431_ (.A(_07153_),
    .B(_07494_),
    .COUT(_07495_),
    .SUM(_07496_));
 sky130_fd_sc_hd__ha_1 _15432_ (.A(_07133_),
    .B(_07497_),
    .COUT(_07498_),
    .SUM(_07499_));
 sky130_fd_sc_hd__ha_1 _15433_ (.A(_07121_),
    .B(_07500_),
    .COUT(_07501_),
    .SUM(_07502_));
 sky130_fd_sc_hd__ha_4 _15434_ (.A(_07112_),
    .B(_07503_),
    .COUT(_07504_),
    .SUM(_07505_));
 sky130_fd_sc_hd__ha_1 _15435_ (.A(_07506_),
    .B(_05892_),
    .COUT(_07507_),
    .SUM(_07508_));
 sky130_fd_sc_hd__ha_1 _15436_ (.A(net14),
    .B(net378),
    .COUT(_07509_),
    .SUM(_07510_));
 sky130_fd_sc_hd__ha_1 _15437_ (.A(_07166_),
    .B(_07511_),
    .COUT(_07512_),
    .SUM(_07513_));
 sky130_fd_sc_hd__ha_1 _15438_ (.A(_07153_),
    .B(_07514_),
    .COUT(_07515_),
    .SUM(_07516_));
 sky130_fd_sc_hd__ha_1 _15439_ (.A(_07133_),
    .B(_07517_),
    .COUT(_07518_),
    .SUM(_07519_));
 sky130_fd_sc_hd__ha_1 _15440_ (.A(_07121_),
    .B(_07520_),
    .COUT(_07521_),
    .SUM(_07522_));
 sky130_fd_sc_hd__ha_4 _15441_ (.A(_07112_),
    .B(_07523_),
    .COUT(_07524_),
    .SUM(_07525_));
 sky130_fd_sc_hd__ha_4 _15442_ (.A(_05892_),
    .B(_07526_),
    .COUT(_07527_),
    .SUM(_07528_));
 sky130_fd_sc_hd__ha_1 _15443_ (.A(net14),
    .B(net379),
    .COUT(_07529_),
    .SUM(_07530_));
 sky130_fd_sc_hd__ha_1 _15444_ (.A(net14),
    .B(net380),
    .COUT(_07531_),
    .SUM(_07532_));
 sky130_fd_sc_hd__ha_1 _15445_ (.A(_07166_),
    .B(_07533_),
    .COUT(_07534_),
    .SUM(_07535_));
 sky130_fd_sc_hd__ha_1 _15446_ (.A(_07153_),
    .B(_07536_),
    .COUT(_07537_),
    .SUM(_07538_));
 sky130_fd_sc_hd__ha_1 _15447_ (.A(_07133_),
    .B(_07539_),
    .COUT(_07540_),
    .SUM(_07541_));
 sky130_fd_sc_hd__ha_1 _15448_ (.A(_07121_),
    .B(_07542_),
    .COUT(_07543_),
    .SUM(_07544_));
 sky130_fd_sc_hd__ha_1 _15449_ (.A(_07545_),
    .B(_07112_),
    .COUT(_07546_),
    .SUM(_07547_));
 sky130_fd_sc_hd__ha_4 _15450_ (.A(_07548_),
    .B(_05892_),
    .COUT(_07549_),
    .SUM(_07550_));
 sky130_fd_sc_hd__ha_1 _15451_ (.A(_07551_),
    .B(_05892_),
    .COUT(_07552_),
    .SUM(_07553_));
 sky130_fd_sc_hd__ha_1 _15452_ (.A(net14),
    .B(net381),
    .COUT(_07554_),
    .SUM(_07555_));
 sky130_fd_sc_hd__ha_1 _15453_ (.A(_07207_),
    .B(_07556_),
    .COUT(_07557_),
    .SUM(_07558_));
 sky130_fd_sc_hd__ha_1 _15454_ (.A(_07166_),
    .B(_07559_),
    .COUT(_07560_),
    .SUM(_07561_));
 sky130_fd_sc_hd__ha_1 _15455_ (.A(_07153_),
    .B(_07562_),
    .COUT(_07563_),
    .SUM(_07564_));
 sky130_fd_sc_hd__ha_1 _15456_ (.A(_07133_),
    .B(_07565_),
    .COUT(_07566_),
    .SUM(_07567_));
 sky130_fd_sc_hd__ha_1 _15457_ (.A(_07121_),
    .B(_07568_),
    .COUT(_07569_),
    .SUM(_07570_));
 sky130_fd_sc_hd__ha_1 _15458_ (.A(_07112_),
    .B(_07571_),
    .COUT(_07572_),
    .SUM(_07573_));
 sky130_fd_sc_hd__ha_1 _15459_ (.A(net14),
    .B(net382),
    .COUT(_07574_),
    .SUM(_07575_));
 sky130_fd_sc_hd__ha_4 _15460_ (.A(_07112_),
    .B(_07576_),
    .COUT(_07577_),
    .SUM(_07578_));
 sky130_fd_sc_hd__ha_4 _15461_ (.A(_07579_),
    .B(_05892_),
    .COUT(_07580_),
    .SUM(_07581_));
 sky130_fd_sc_hd__ha_1 _15462_ (.A(_07207_),
    .B(_07582_),
    .COUT(_07583_),
    .SUM(_07584_));
 sky130_fd_sc_hd__ha_1 _15463_ (.A(_07166_),
    .B(_07585_),
    .COUT(_07586_),
    .SUM(_07587_));
 sky130_fd_sc_hd__ha_1 _15464_ (.A(_07153_),
    .B(_07588_),
    .COUT(_07589_),
    .SUM(_07590_));
 sky130_fd_sc_hd__ha_1 _15465_ (.A(_07133_),
    .B(_07591_),
    .COUT(_07592_),
    .SUM(_07593_));
 sky130_fd_sc_hd__ha_1 _15466_ (.A(_07121_),
    .B(_07594_),
    .COUT(_07595_),
    .SUM(_07596_));
 sky130_fd_sc_hd__ha_1 _15467_ (.A(_07121_),
    .B(_07597_),
    .COUT(_07598_),
    .SUM(_07599_));
 sky130_fd_sc_hd__ha_4 _15468_ (.A(_07112_),
    .B(_07600_),
    .COUT(_07601_),
    .SUM(_07602_));
 sky130_fd_sc_hd__ha_4 _15469_ (.A(_05892_),
    .B(_07603_),
    .COUT(_07604_),
    .SUM(_07605_));
 sky130_fd_sc_hd__ha_1 _15470_ (.A(net14),
    .B(net383),
    .COUT(_07606_),
    .SUM(_07607_));
 sky130_fd_sc_hd__ha_1 _15471_ (.A(_07207_),
    .B(_07608_),
    .COUT(_07609_),
    .SUM(_07610_));
 sky130_fd_sc_hd__ha_1 _15472_ (.A(_07166_),
    .B(_07611_),
    .COUT(_07612_),
    .SUM(_07613_));
 sky130_fd_sc_hd__ha_1 _15473_ (.A(_07153_),
    .B(_07614_),
    .COUT(_07615_),
    .SUM(_07616_));
 sky130_fd_sc_hd__ha_1 _15474_ (.A(_07133_),
    .B(_07617_),
    .COUT(_07618_),
    .SUM(_07619_));
 sky130_fd_sc_hd__ha_1 _15475_ (.A(net14),
    .B(net384),
    .COUT(_07620_),
    .SUM(_07621_));
 sky130_fd_sc_hd__ha_4 _15476_ (.A(_07112_),
    .B(_07622_),
    .COUT(_07623_),
    .SUM(_07624_));
 sky130_fd_sc_hd__ha_4 _15477_ (.A(_05892_),
    .B(_07625_),
    .COUT(_07626_),
    .SUM(_07627_));
 sky130_fd_sc_hd__ha_1 _15478_ (.A(_07133_),
    .B(_07628_),
    .COUT(_07629_),
    .SUM(_07630_));
 sky130_fd_sc_hd__ha_1 _15479_ (.A(_07121_),
    .B(_07631_),
    .COUT(_07632_),
    .SUM(_07633_));
 sky130_fd_sc_hd__ha_1 _15480_ (.A(_07166_),
    .B(_07634_),
    .COUT(_07635_),
    .SUM(_07636_));
 sky130_fd_sc_hd__ha_1 _15481_ (.A(_07153_),
    .B(_07637_),
    .COUT(_07638_),
    .SUM(_07639_));
 sky130_fd_sc_hd__ha_1 _15482_ (.A(_07207_),
    .B(_07640_),
    .COUT(_07641_),
    .SUM(_07642_));
 sky130_fd_sc_hd__ha_4 _15483_ (.A(_07643_),
    .B(_05892_),
    .COUT(_07644_),
    .SUM(_07645_));
 sky130_fd_sc_hd__ha_1 _15484_ (.A(\butterfly_count[2] ),
    .B(net14),
    .COUT(_07646_),
    .SUM(_07647_));
 sky130_fd_sc_hd__ha_1 _15485_ (.A(_07153_),
    .B(_07648_),
    .COUT(_07649_),
    .SUM(_07650_));
 sky130_fd_sc_hd__ha_1 _15486_ (.A(_07133_),
    .B(_07651_),
    .COUT(_07652_),
    .SUM(_07653_));
 sky130_fd_sc_hd__ha_1 _15487_ (.A(_07121_),
    .B(_07654_),
    .COUT(_07655_),
    .SUM(_07656_));
 sky130_fd_sc_hd__ha_1 _15488_ (.A(_07657_),
    .B(_07112_),
    .COUT(_07658_),
    .SUM(_07659_));
 sky130_fd_sc_hd__ha_1 _15489_ (.A(_07207_),
    .B(_07660_),
    .COUT(_07661_),
    .SUM(_07662_));
 sky130_fd_sc_hd__ha_1 _15490_ (.A(_07166_),
    .B(_07663_),
    .COUT(_07664_),
    .SUM(_07665_));
 sky130_fd_sc_hd__ha_1 _15491_ (.A(_07666_),
    .B(_07667_),
    .COUT(_07668_),
    .SUM(_07669_));
 sky130_fd_sc_hd__ha_1 _15492_ (.A(\butterfly_count[1] ),
    .B(net14),
    .COUT(_07670_),
    .SUM(_07671_));
 sky130_fd_sc_hd__ha_4 _15493_ (.A(_07112_),
    .B(_07672_),
    .COUT(_07673_),
    .SUM(_07674_));
 sky130_fd_sc_hd__ha_4 _15494_ (.A(_05892_),
    .B(_07675_),
    .COUT(_07676_),
    .SUM(_07677_));
 sky130_fd_sc_hd__ha_2 _15495_ (.A(_07166_),
    .B(_07678_),
    .COUT(_07679_),
    .SUM(_07680_));
 sky130_fd_sc_hd__ha_1 _15496_ (.A(_07153_),
    .B(_07681_),
    .COUT(_07682_),
    .SUM(_07683_));
 sky130_fd_sc_hd__ha_1 _15497_ (.A(_07133_),
    .B(_07684_),
    .COUT(_07685_),
    .SUM(_07686_));
 sky130_fd_sc_hd__ha_1 _15498_ (.A(_07121_),
    .B(_07687_),
    .COUT(_07688_),
    .SUM(_07689_));
 sky130_fd_sc_hd__ha_1 _15499_ (.A(_07690_),
    .B(_07691_),
    .COUT(_07692_),
    .SUM(_07693_));
 sky130_fd_sc_hd__ha_1 _15500_ (.A(_07695_),
    .B(_07694_),
    .COUT(_07696_),
    .SUM(_07697_));
 sky130_fd_sc_hd__ha_4 _15501_ (.A(_07698_),
    .B(_07699_),
    .COUT(_07700_),
    .SUM(_07701_));
 sky130_fd_sc_hd__ha_1 _15502_ (.A(_07702_),
    .B(_07703_),
    .COUT(_07704_),
    .SUM(_07705_));
 sky130_fd_sc_hd__ha_1 _15503_ (.A(_07706_),
    .B(_07707_),
    .COUT(_07708_),
    .SUM(_07709_));
 sky130_fd_sc_hd__ha_1 _15504_ (.A(_07710_),
    .B(_07711_),
    .COUT(_07712_),
    .SUM(_07713_));
 sky130_fd_sc_hd__ha_1 _15505_ (.A(_05892_),
    .B(_05893_),
    .COUT(_07714_),
    .SUM(_07715_));
 sky130_fd_sc_hd__ha_1 _15506_ (.A(_07716_),
    .B(net386),
    .COUT(_07717_),
    .SUM(_07718_));
 sky130_fd_sc_hd__ha_1 _15507_ (.A(\butterfly_count[0] ),
    .B(net14),
    .COUT(_07719_),
    .SUM(_07720_));
 sky130_fd_sc_hd__ha_2 _15508_ (.A(_05882_),
    .B(_07721_),
    .COUT(_07722_),
    .SUM(_07723_));
 sky130_fd_sc_hd__ha_1 _15509_ (.A(\temp_real[0] ),
    .B(_07721_),
    .COUT(_07724_),
    .SUM(_07725_));
 sky130_fd_sc_hd__ha_1 _15510_ (.A(_05882_),
    .B(_07726_),
    .COUT(_07727_),
    .SUM(_07728_));
 sky130_fd_sc_hd__ha_1 _15511_ (.A(net53),
    .B(_07726_),
    .COUT(_07729_),
    .SUM(_07730_));
 sky130_fd_sc_hd__ha_4 _15512_ (.A(net53),
    .B(net610),
    .COUT(_07731_),
    .SUM(_07733_));
 sky130_fd_sc_hd__ha_4 _15513_ (.A(net53),
    .B(_07734_),
    .COUT(_05891_),
    .SUM(_07735_));
 sky130_fd_sc_hd__ha_1 _15514_ (.A(_07736_),
    .B(_07737_),
    .COUT(_07738_),
    .SUM(_07739_));
 sky130_fd_sc_hd__ha_1 _15515_ (.A(_05882_),
    .B(_07740_),
    .COUT(_07741_),
    .SUM(_07742_));
 sky130_fd_sc_hd__ha_1 _15516_ (.A(net53),
    .B(_07740_),
    .COUT(_07743_),
    .SUM(_07744_));
 sky130_fd_sc_hd__ha_1 _15517_ (.A(_05882_),
    .B(_07745_),
    .COUT(_07746_),
    .SUM(_07747_));
 sky130_fd_sc_hd__ha_1 _15518_ (.A(net53),
    .B(_07745_),
    .COUT(_07748_),
    .SUM(_07749_));
 sky130_fd_sc_hd__ha_1 _15519_ (.A(_05882_),
    .B(_07750_),
    .COUT(_07751_),
    .SUM(_07752_));
 sky130_fd_sc_hd__ha_1 _15520_ (.A(net53),
    .B(_07750_),
    .COUT(_07753_),
    .SUM(_07754_));
 sky130_fd_sc_hd__ha_1 _15521_ (.A(_05882_),
    .B(_07755_),
    .COUT(_07756_),
    .SUM(_07757_));
 sky130_fd_sc_hd__ha_1 _15522_ (.A(net53),
    .B(_07755_),
    .COUT(_07758_),
    .SUM(_07759_));
 sky130_fd_sc_hd__ha_1 _15523_ (.A(_05882_),
    .B(_07760_),
    .COUT(_07761_),
    .SUM(_07762_));
 sky130_fd_sc_hd__ha_1 _15524_ (.A(net53),
    .B(_07760_),
    .COUT(_07763_),
    .SUM(_07764_));
 sky130_fd_sc_hd__ha_1 _15525_ (.A(_05882_),
    .B(_07765_),
    .COUT(_07766_),
    .SUM(_07767_));
 sky130_fd_sc_hd__ha_1 _15526_ (.A(net53),
    .B(_07765_),
    .COUT(_07768_),
    .SUM(_07769_));
 sky130_fd_sc_hd__ha_1 _15527_ (.A(_05882_),
    .B(_07770_),
    .COUT(_07771_),
    .SUM(_07772_));
 sky130_fd_sc_hd__ha_1 _15528_ (.A(net53),
    .B(_07770_),
    .COUT(_07773_),
    .SUM(_07774_));
 sky130_fd_sc_hd__ha_1 _15529_ (.A(_05882_),
    .B(_07775_),
    .COUT(_07776_),
    .SUM(_07777_));
 sky130_fd_sc_hd__ha_1 _15530_ (.A(net53),
    .B(_07775_),
    .COUT(_07778_),
    .SUM(_07779_));
 sky130_fd_sc_hd__ha_1 _15531_ (.A(_05882_),
    .B(_07780_),
    .COUT(_07781_),
    .SUM(_07782_));
 sky130_fd_sc_hd__ha_1 _15532_ (.A(net53),
    .B(_07780_),
    .COUT(_07783_),
    .SUM(_07784_));
 sky130_fd_sc_hd__ha_4 _15533_ (.A(_05882_),
    .B(_07785_),
    .COUT(_07786_),
    .SUM(_07787_));
 sky130_fd_sc_hd__ha_1 _15534_ (.A(net53),
    .B(_07785_),
    .COUT(_07788_),
    .SUM(_07789_));
 sky130_fd_sc_hd__ha_4 _15535_ (.A(_07790_),
    .B(_05882_),
    .COUT(_07791_),
    .SUM(_07792_));
 sky130_fd_sc_hd__ha_1 _15536_ (.A(net53),
    .B(_07790_),
    .COUT(_07793_),
    .SUM(_07794_));
 sky130_fd_sc_hd__ha_4 _15537_ (.A(_05887_),
    .B(_05882_),
    .COUT(_07795_),
    .SUM(_07796_));
 sky130_fd_sc_hd__ha_2 _15538_ (.A(net53),
    .B(net594),
    .COUT(_07797_),
    .SUM(_07798_));
 sky130_fd_sc_hd__ha_1 _15539_ (.A(_07716_),
    .B(_07666_),
    .COUT(_07799_),
    .SUM(_07800_));
 sky130_fd_sc_hd__ha_1 _15540_ (.A(\butterfly_count[0] ),
    .B(\butterfly_count[1] ),
    .COUT(_07801_),
    .SUM(_07802_));
 sky130_fd_sc_hd__ha_4 _15541_ (.A(_07804_),
    .B(_07803_),
    .COUT(_07805_),
    .SUM(_07806_));
 sky130_fd_sc_hd__ha_1 _15542_ (.A(_07803_),
    .B(_07804_),
    .COUT(_07807_),
    .SUM(_07808_));
 sky130_fd_sc_hd__ha_1 _15543_ (.A(_07803_),
    .B(\stage[1] ),
    .COUT(_07809_),
    .SUM(_07810_));
 sky130_fd_sc_hd__ha_4 _15544_ (.A(\stage[0] ),
    .B(_07804_),
    .COUT(_07811_),
    .SUM(_07812_));
 sky130_fd_sc_hd__ha_1 _15545_ (.A(\stage[0] ),
    .B(_07804_),
    .COUT(_07813_),
    .SUM(_07814_));
 sky130_fd_sc_hd__ha_2 _15546_ (.A(\stage[0] ),
    .B(\stage[1] ),
    .COUT(_07815_),
    .SUM(_07816_));
 sky130_fd_sc_hd__ha_2 _15547_ (.A(_07817_),
    .B(_07818_),
    .COUT(_07819_),
    .SUM(_07820_));
 sky130_fd_sc_hd__ha_4 _15548_ (.A(_07817_),
    .B(_07815_),
    .COUT(_07821_),
    .SUM(_07822_));
 sky130_fd_sc_hd__ha_4 _15549_ (.A(_07817_),
    .B(_07815_),
    .COUT(_07706_),
    .SUM(_07823_));
 sky130_fd_sc_hd__ha_1 _15550_ (.A(\stage[2] ),
    .B(_07815_),
    .COUT(_07824_),
    .SUM(_07825_));
 sky130_fd_sc_hd__ha_4 _15551_ (.A(\stage[2] ),
    .B(_07815_),
    .COUT(_07690_),
    .SUM(_07826_));
 sky130_fd_sc_hd__ha_1 _15552_ (.A(_07827_),
    .B(_07828_),
    .COUT(_07829_),
    .SUM(_07830_));
 sky130_fd_sc_hd__ha_1 _15553_ (.A(\sample_count[0] ),
    .B(\sample_count[1] ),
    .COUT(_07831_),
    .SUM(_07832_));
 sky130_fd_sc_hd__ha_1 _15554_ (.A(\sample_count[2] ),
    .B(_07831_),
    .COUT(_07833_),
    .SUM(_07834_));
 sky130_fd_sc_hd__ha_2 _15555_ (.A(_05897_),
    .B(_07835_),
    .COUT(_07836_),
    .SUM(_07837_));
 sky130_fd_sc_hd__ha_1 _15556_ (.A(\temp_imag[0] ),
    .B(_07835_),
    .COUT(_07838_),
    .SUM(_07839_));
 sky130_fd_sc_hd__ha_1 _15557_ (.A(_05897_),
    .B(_07840_),
    .COUT(_07841_),
    .SUM(_07842_));
 sky130_fd_sc_hd__ha_1 _15558_ (.A(\temp_imag[0] ),
    .B(_07840_),
    .COUT(_07843_),
    .SUM(_07844_));
 sky130_fd_sc_hd__ha_4 _15559_ (.A(\temp_imag[0] ),
    .B(net637),
    .COUT(_07845_),
    .SUM(_07847_));
 sky130_fd_sc_hd__ha_4 _15560_ (.A(\temp_imag[0] ),
    .B(_07848_),
    .COUT(_05906_),
    .SUM(_07849_));
 sky130_fd_sc_hd__ha_1 _15561_ (.A(_07850_),
    .B(_07851_),
    .COUT(_07852_),
    .SUM(_07853_));
 sky130_fd_sc_hd__ha_1 _15562_ (.A(_05897_),
    .B(_07854_),
    .COUT(_07855_),
    .SUM(_07856_));
 sky130_fd_sc_hd__ha_1 _15563_ (.A(\temp_imag[0] ),
    .B(_07854_),
    .COUT(_07857_),
    .SUM(_07858_));
 sky130_fd_sc_hd__ha_1 _15564_ (.A(_05897_),
    .B(_07859_),
    .COUT(_07860_),
    .SUM(_07861_));
 sky130_fd_sc_hd__ha_1 _15565_ (.A(\temp_imag[0] ),
    .B(_07859_),
    .COUT(_07862_),
    .SUM(_07863_));
 sky130_fd_sc_hd__ha_1 _15566_ (.A(_05897_),
    .B(_07864_),
    .COUT(_07865_),
    .SUM(_07866_));
 sky130_fd_sc_hd__ha_1 _15567_ (.A(\temp_imag[0] ),
    .B(_07864_),
    .COUT(_07867_),
    .SUM(_07868_));
 sky130_fd_sc_hd__ha_1 _15568_ (.A(_05897_),
    .B(_07869_),
    .COUT(_07870_),
    .SUM(_07871_));
 sky130_fd_sc_hd__ha_1 _15569_ (.A(\temp_imag[0] ),
    .B(_07869_),
    .COUT(_07872_),
    .SUM(_07873_));
 sky130_fd_sc_hd__ha_1 _15570_ (.A(_05897_),
    .B(_07874_),
    .COUT(_07875_),
    .SUM(_07876_));
 sky130_fd_sc_hd__ha_1 _15571_ (.A(\temp_imag[0] ),
    .B(_07874_),
    .COUT(_07877_),
    .SUM(_07878_));
 sky130_fd_sc_hd__ha_1 _15572_ (.A(_05897_),
    .B(_07879_),
    .COUT(_07880_),
    .SUM(_07881_));
 sky130_fd_sc_hd__ha_1 _15573_ (.A(\temp_imag[0] ),
    .B(_07879_),
    .COUT(_07882_),
    .SUM(_07883_));
 sky130_fd_sc_hd__ha_1 _15574_ (.A(_05897_),
    .B(_07884_),
    .COUT(_07885_),
    .SUM(_07886_));
 sky130_fd_sc_hd__ha_1 _15575_ (.A(\temp_imag[0] ),
    .B(_07884_),
    .COUT(_07887_),
    .SUM(_07888_));
 sky130_fd_sc_hd__ha_1 _15576_ (.A(_05897_),
    .B(_07889_),
    .COUT(_07890_),
    .SUM(_07891_));
 sky130_fd_sc_hd__ha_1 _15577_ (.A(\temp_imag[0] ),
    .B(_07889_),
    .COUT(_07892_),
    .SUM(_07893_));
 sky130_fd_sc_hd__ha_1 _15578_ (.A(_05897_),
    .B(_07894_),
    .COUT(_07895_),
    .SUM(_07896_));
 sky130_fd_sc_hd__ha_1 _15579_ (.A(\temp_imag[0] ),
    .B(_07894_),
    .COUT(_07897_),
    .SUM(_07898_));
 sky130_fd_sc_hd__ha_4 _15580_ (.A(_05897_),
    .B(_07899_),
    .COUT(_07900_),
    .SUM(_07901_));
 sky130_fd_sc_hd__ha_1 _15581_ (.A(\temp_imag[0] ),
    .B(_07899_),
    .COUT(_07902_),
    .SUM(_07903_));
 sky130_fd_sc_hd__ha_4 _15582_ (.A(_05897_),
    .B(_07904_),
    .COUT(_07905_),
    .SUM(_07906_));
 sky130_fd_sc_hd__ha_1 _15583_ (.A(\temp_imag[0] ),
    .B(_07904_),
    .COUT(_07907_),
    .SUM(_07908_));
 sky130_fd_sc_hd__ha_1 _15584_ (.A(_05902_),
    .B(_05897_),
    .COUT(_07909_),
    .SUM(_07910_));
 sky130_fd_sc_hd__ha_1 _15585_ (.A(\temp_imag[0] ),
    .B(_05902_),
    .COUT(_07911_),
    .SUM(_07912_));
 sky130_fd_sc_hd__ha_1 _15586_ (.A(\butterfly_in_group[0] ),
    .B(_07913_),
    .COUT(_07914_),
    .SUM(_05879_));
 sky130_fd_sc_hd__ha_1 _15587_ (.A(\butterfly_in_group[1] ),
    .B(_07915_),
    .COUT(_07916_),
    .SUM(_07917_));
 sky130_fd_sc_hd__ha_1 _15588_ (.A(_07917_),
    .B(_07918_),
    .COUT(_07919_),
    .SUM(_07920_));
 sky130_fd_sc_hd__ha_1 _15589_ (.A(_07920_),
    .B(_07914_),
    .COUT(_07921_),
    .SUM(_05880_));
 sky130_fd_sc_hd__ha_1 _15590_ (.A(net387),
    .B(_05879_),
    .COUT(_05908_),
    .SUM(_05881_));
 sky130_fd_sc_hd__ha_1 _15591_ (.A(_05912_),
    .B(_05913_),
    .COUT(_07922_),
    .SUM(_07923_));
 sky130_fd_sc_hd__ha_1 _15592_ (.A(_06123_),
    .B(_06175_),
    .COUT(_07924_),
    .SUM(_07925_));
 sky130_fd_sc_hd__ha_1 _15593_ (.A(_06124_),
    .B(_06235_),
    .COUT(_07926_),
    .SUM(_05943_));
 sky130_fd_sc_hd__ha_1 _15594_ (.A(_05945_),
    .B(_07928_),
    .COUT(_07929_),
    .SUM(_07930_));
 sky130_fd_sc_hd__ha_1 _15595_ (.A(_05951_),
    .B(_07931_),
    .COUT(_07932_),
    .SUM(_07933_));
 sky130_fd_sc_hd__ha_1 _15596_ (.A(_06175_),
    .B(_06501_),
    .COUT(_05944_),
    .SUM(_05985_));
 sky130_fd_sc_hd__ha_1 _15597_ (.A(_05987_),
    .B(_06371_),
    .COUT(_06012_),
    .SUM(_07935_));
 sky130_fd_sc_hd__ha_1 _15598_ (.A(_07936_),
    .B(_05997_),
    .COUT(_07937_),
    .SUM(_06077_));
 sky130_fd_sc_hd__ha_1 _15599_ (.A(_07938_),
    .B(_07939_),
    .COUT(_07940_),
    .SUM(_07941_));
 sky130_fd_sc_hd__ha_1 _15600_ (.A(_06201_),
    .B(_06202_),
    .COUT(_07942_),
    .SUM(_07943_));
 sky130_fd_sc_hd__ha_1 _15601_ (.A(_07944_),
    .B(_07943_),
    .COUT(_07945_),
    .SUM(_07946_));
 sky130_fd_sc_hd__ha_1 _15602_ (.A(_07938_),
    .B(_05912_),
    .COUT(_06052_),
    .SUM(_07947_));
 sky130_fd_sc_hd__ha_1 _15603_ (.A(_06235_),
    .B(_07928_),
    .COUT(_05986_),
    .SUM(_07949_));
 sky130_fd_sc_hd__ha_1 _15604_ (.A(_05998_),
    .B(_07950_),
    .COUT(_06078_),
    .SUM(_06128_));
 sky130_fd_sc_hd__ha_1 _15605_ (.A(_06079_),
    .B(_06131_),
    .COUT(_06106_),
    .SUM(_06114_));
 sky130_fd_sc_hd__ha_1 _15606_ (.A(_07951_),
    .B(_06382_),
    .COUT(_07948_),
    .SUM(_07952_));
 sky130_fd_sc_hd__ha_1 _15607_ (.A(_07952_),
    .B(_07953_),
    .COUT(_07954_),
    .SUM(_06142_));
 sky130_fd_sc_hd__ha_1 _15608_ (.A(_07955_),
    .B(_06285_),
    .COUT(_07956_),
    .SUM(_07957_));
 sky130_fd_sc_hd__ha_1 _15609_ (.A(_06175_),
    .B(_06235_),
    .COUT(_07958_),
    .SUM(_07959_));
 sky130_fd_sc_hd__ha_1 _15610_ (.A(_06501_),
    .B(_06371_),
    .COUT(_07960_),
    .SUM(_07961_));
 sky130_fd_sc_hd__ha_1 _15611_ (.A(_07958_),
    .B(_07961_),
    .COUT(_06167_),
    .SUM(_07962_));
 sky130_fd_sc_hd__ha_1 _15612_ (.A(_07963_),
    .B(_07964_),
    .COUT(_06129_),
    .SUM(_06178_));
 sky130_fd_sc_hd__ha_1 _15613_ (.A(_06132_),
    .B(_06181_),
    .COUT(_06152_),
    .SUM(_06163_));
 sky130_fd_sc_hd__ha_1 _15614_ (.A(_07943_),
    .B(_06034_),
    .COUT(_06145_),
    .SUM(_06195_));
 sky130_fd_sc_hd__ha_1 _15615_ (.A(_07965_),
    .B(_07966_),
    .COUT(_07967_),
    .SUM(_06193_));
 sky130_fd_sc_hd__ha_1 _15616_ (.A(_06150_),
    .B(_07954_),
    .COUT(_07968_),
    .SUM(_06154_));
 sky130_fd_sc_hd__ha_1 _15617_ (.A(_06235_),
    .B(_06501_),
    .COUT(_07969_),
    .SUM(_07970_));
 sky130_fd_sc_hd__ha_1 _15618_ (.A(_07928_),
    .B(_07969_),
    .COUT(_06227_),
    .SUM(_07971_));
 sky130_fd_sc_hd__ha_1 _15619_ (.A(_07972_),
    .B(_06185_),
    .COUT(_06179_),
    .SUM(_06238_));
 sky130_fd_sc_hd__ha_1 _15620_ (.A(_06182_),
    .B(_06241_),
    .COUT(_06205_),
    .SUM(_06223_));
 sky130_fd_sc_hd__ha_1 _15621_ (.A(_06382_),
    .B(_06203_),
    .COUT(_06196_),
    .SUM(_07973_));
 sky130_fd_sc_hd__ha_1 _15622_ (.A(_05913_),
    .B(_05937_),
    .COUT(_07974_),
    .SUM(_07975_));
 sky130_fd_sc_hd__ha_1 _15623_ (.A(_07976_),
    .B(_07977_),
    .COUT(_07978_),
    .SUM(_07979_));
 sky130_fd_sc_hd__ha_1 _15624_ (.A(_07981_),
    .B(_07967_),
    .COUT(_06211_),
    .SUM(_06215_));
 sky130_fd_sc_hd__ha_1 _15625_ (.A(_06371_),
    .B(_07982_),
    .COUT(_06277_),
    .SUM(_07983_));
 sky130_fd_sc_hd__ha_1 _15626_ (.A(_06186_),
    .B(_07984_),
    .COUT(_06239_),
    .SUM(_06288_));
 sky130_fd_sc_hd__ha_1 _15627_ (.A(_06242_),
    .B(_06291_),
    .COUT(_06256_),
    .SUM(_06273_));
 sky130_fd_sc_hd__ha_1 _15628_ (.A(_06249_),
    .B(_07973_),
    .COUT(_07980_),
    .SUM(_07985_));
 sky130_fd_sc_hd__ha_1 _15629_ (.A(_06032_),
    .B(_06382_),
    .COUT(_07986_),
    .SUM(_06298_));
 sky130_fd_sc_hd__ha_1 _15630_ (.A(_05937_),
    .B(_05938_),
    .COUT(_07987_),
    .SUM(_07988_));
 sky130_fd_sc_hd__ha_1 _15631_ (.A(_05925_),
    .B(_05918_),
    .COUT(_07989_),
    .SUM(_07990_));
 sky130_fd_sc_hd__ha_1 _15632_ (.A(_07992_),
    .B(_07978_),
    .COUT(_06261_),
    .SUM(_06265_));
 sky130_fd_sc_hd__ha_1 _15633_ (.A(_06213_),
    .B(_06262_),
    .COUT(_07993_),
    .SUM(_07994_));
 sky130_fd_sc_hd__ha_1 _15634_ (.A(_07995_),
    .B(_07996_),
    .COUT(_06289_),
    .SUM(_06335_));
 sky130_fd_sc_hd__ha_1 _15635_ (.A(_06292_),
    .B(_06338_),
    .COUT(_06310_),
    .SUM(_06324_));
 sky130_fd_sc_hd__ha_1 _15636_ (.A(_05938_),
    .B(_05980_),
    .COUT(_07997_),
    .SUM(_07998_));
 sky130_fd_sc_hd__ha_1 _15637_ (.A(_07927_),
    .B(_05935_),
    .COUT(_07999_),
    .SUM(_08000_));
 sky130_fd_sc_hd__ha_1 _15638_ (.A(_06299_),
    .B(_07986_),
    .COUT(_07991_),
    .SUM(_08001_));
 sky130_fd_sc_hd__ha_1 _15639_ (.A(_06308_),
    .B(_07989_),
    .COUT(_06312_),
    .SUM(_06316_));
 sky130_fd_sc_hd__ha_1 _15640_ (.A(_06263_),
    .B(_06313_),
    .COUT(_08002_),
    .SUM(_08003_));
 sky130_fd_sc_hd__ha_1 _15641_ (.A(_08004_),
    .B(_08005_),
    .COUT(_06323_),
    .SUM(_06363_));
 sky130_fd_sc_hd__ha_1 _15642_ (.A(_08006_),
    .B(_08007_),
    .COUT(_06336_),
    .SUM(_06373_));
 sky130_fd_sc_hd__ha_4 _15643_ (.A(_06376_),
    .B(_06339_),
    .COUT(_08008_),
    .SUM(_06365_));
 sky130_fd_sc_hd__ha_1 _15644_ (.A(_08000_),
    .B(_08001_),
    .COUT(_06307_),
    .SUM(_06349_));
 sky130_fd_sc_hd__ha_1 _15645_ (.A(_05980_),
    .B(_06123_),
    .COUT(_05942_),
    .SUM(_08009_));
 sky130_fd_sc_hd__ha_1 _15646_ (.A(_07934_),
    .B(_05978_),
    .COUT(_08010_),
    .SUM(_08011_));
 sky130_fd_sc_hd__ha_1 _15647_ (.A(_06351_),
    .B(_07999_),
    .COUT(_06354_),
    .SUM(_06358_));
 sky130_fd_sc_hd__ha_1 _15648_ (.A(_06314_),
    .B(_06355_),
    .COUT(_08012_),
    .SUM(_08013_));
 sky130_fd_sc_hd__ha_1 _15649_ (.A(_08015_),
    .B(_08014_),
    .COUT(_06364_),
    .SUM(_06400_));
 sky130_fd_sc_hd__ha_1 _15650_ (.A(_08016_),
    .B(_08017_),
    .COUT(_08015_),
    .SUM(_08018_));
 sky130_fd_sc_hd__ha_1 _15651_ (.A(_07928_),
    .B(_06434_),
    .COUT(_06372_),
    .SUM(_06456_));
 sky130_fd_sc_hd__ha_4 _15652_ (.A(_06380_),
    .B(_08019_),
    .COUT(_06374_),
    .SUM(_06409_));
 sky130_fd_sc_hd__ha_1 _15653_ (.A(_06383_),
    .B(_08020_),
    .COUT(_08021_),
    .SUM(_06406_));
 sky130_fd_sc_hd__ha_1 _15654_ (.A(_06377_),
    .B(_08022_),
    .COUT(_08023_),
    .SUM(_06402_));
 sky130_fd_sc_hd__ha_1 _15655_ (.A(_08011_),
    .B(_06346_),
    .COUT(_06350_),
    .SUM(_06385_));
 sky130_fd_sc_hd__ha_1 _15656_ (.A(_06123_),
    .B(_06124_),
    .COUT(_05984_),
    .SUM(_08024_));
 sky130_fd_sc_hd__ha_1 _15657_ (.A(_06072_),
    .B(_06067_),
    .COUT(_08025_),
    .SUM(_08026_));
 sky130_fd_sc_hd__ha_1 _15658_ (.A(_06387_),
    .B(_08010_),
    .COUT(_06390_),
    .SUM(_06394_));
 sky130_fd_sc_hd__ha_1 _15659_ (.A(_06356_),
    .B(_06391_),
    .COUT(_08027_),
    .SUM(_08028_));
 sky130_fd_sc_hd__ha_1 _15660_ (.A(_08018_),
    .B(_08029_),
    .COUT(_06401_),
    .SUM(_08030_));
 sky130_fd_sc_hd__ha_1 _15661_ (.A(_06381_),
    .B(_08031_),
    .COUT(_06410_),
    .SUM(_06432_));
 sky130_fd_sc_hd__ha_1 _15662_ (.A(_06046_),
    .B(_08032_),
    .COUT(_08031_),
    .SUM(_08033_));
 sky130_fd_sc_hd__ha_1 _15663_ (.A(_06202_),
    .B(_06382_),
    .COUT(_08020_),
    .SUM(_08034_));
 sky130_fd_sc_hd__ha_1 _15664_ (.A(_08034_),
    .B(_08035_),
    .COUT(_08036_),
    .SUM(_06429_));
 sky130_fd_sc_hd__ha_4 _15665_ (.A(_08038_),
    .B(_08037_),
    .COUT(_08039_),
    .SUM(_08040_));
 sky130_fd_sc_hd__ha_1 _15666_ (.A(_08026_),
    .B(_08021_),
    .COUT(_06386_),
    .SUM(_06412_));
 sky130_fd_sc_hd__ha_1 _15667_ (.A(_06175_),
    .B(_06124_),
    .COUT(_08041_),
    .SUM(_08042_));
 sky130_fd_sc_hd__ha_1 _15668_ (.A(_08043_),
    .B(_06121_),
    .COUT(_08044_),
    .SUM(_08045_));
 sky130_fd_sc_hd__ha_1 _15669_ (.A(_06414_),
    .B(_08025_),
    .COUT(_06417_),
    .SUM(_06421_));
 sky130_fd_sc_hd__ha_1 _15670_ (.A(_06392_),
    .B(_06418_),
    .COUT(_08046_),
    .SUM(_08047_));
 sky130_fd_sc_hd__ha_4 _15671_ (.A(_08040_),
    .B(_08030_),
    .COUT(_06426_),
    .SUM(_06450_));
 sky130_fd_sc_hd__ha_1 _15672_ (.A(_08048_),
    .B(_08049_),
    .COUT(_08029_),
    .SUM(_08050_));
 sky130_fd_sc_hd__ha_1 _15673_ (.A(_08033_),
    .B(_06437_),
    .COUT(_06433_),
    .SUM(_06463_));
 sky130_fd_sc_hd__ha_1 _15674_ (.A(_06382_),
    .B(_08051_),
    .COUT(_08035_),
    .SUM(_06460_));
 sky130_fd_sc_hd__ha_1 _15675_ (.A(_08052_),
    .B(_08053_),
    .COUT(_08054_),
    .SUM(_08055_));
 sky130_fd_sc_hd__ha_1 _15676_ (.A(_08045_),
    .B(_08036_),
    .COUT(_06413_),
    .SUM(_08056_));
 sky130_fd_sc_hd__ha_1 _15677_ (.A(_08057_),
    .B(_08056_),
    .COUT(_08058_),
    .SUM(_06446_));
 sky130_fd_sc_hd__ha_1 _15678_ (.A(_08058_),
    .B(_08044_),
    .COUT(_06440_),
    .SUM(_06444_));
 sky130_fd_sc_hd__ha_1 _15679_ (.A(_06419_),
    .B(_06441_),
    .COUT(_08059_),
    .SUM(_08060_));
 sky130_fd_sc_hd__ha_1 _15680_ (.A(_08050_),
    .B(_08055_),
    .COUT(_06451_),
    .SUM(_08061_));
 sky130_fd_sc_hd__ha_1 _15681_ (.A(_06438_),
    .B(_06468_),
    .COUT(_06464_),
    .SUM(_08062_));
 sky130_fd_sc_hd__ha_1 _15682_ (.A(_08063_),
    .B(_08064_),
    .COUT(_08065_),
    .SUM(_08066_));
 sky130_fd_sc_hd__ha_1 _15683_ (.A(_08067_),
    .B(_08068_),
    .COUT(_08069_),
    .SUM(_06479_));
 sky130_fd_sc_hd__ha_1 _15684_ (.A(_06442_),
    .B(_06472_),
    .COUT(_08070_),
    .SUM(_08071_));
 sky130_fd_sc_hd__ha_1 _15685_ (.A(_08072_),
    .B(_08066_),
    .COUT(_08073_),
    .SUM(_06492_));
 sky130_fd_sc_hd__ha_1 _15686_ (.A(_06371_),
    .B(_06465_),
    .COUT(_06457_),
    .SUM(_08074_));
 sky130_fd_sc_hd__ha_1 _15687_ (.A(_08075_),
    .B(_08076_),
    .COUT(_08077_),
    .SUM(_08078_));
 sky130_fd_sc_hd__ha_1 _15688_ (.A(_06469_),
    .B(_08079_),
    .COUT(_08080_),
    .SUM(_08081_));
 sky130_fd_sc_hd__ha_1 _15689_ (.A(_08082_),
    .B(_08083_),
    .COUT(_08084_),
    .SUM(_08085_));
 sky130_fd_sc_hd__ha_1 _15690_ (.A(_08086_),
    .B(_08087_),
    .COUT(_08088_),
    .SUM(_08089_));
 sky130_fd_sc_hd__ha_1 _15691_ (.A(_06235_),
    .B(_06481_),
    .COUT(_08090_),
    .SUM(_08091_));
 sky130_fd_sc_hd__ha_1 _15692_ (.A(_06482_),
    .B(_08091_),
    .COUT(_08092_),
    .SUM(_08093_));
 sky130_fd_sc_hd__ha_1 _15693_ (.A(_08092_),
    .B(_08090_),
    .COUT(_06486_),
    .SUM(_08094_));
 sky130_fd_sc_hd__ha_1 _15694_ (.A(_06487_),
    .B(_06473_),
    .COUT(_08095_),
    .SUM(_08096_));
 sky130_fd_sc_hd__ha_1 _15695_ (.A(_08097_),
    .B(_08098_),
    .COUT(_06496_),
    .SUM(_08099_));
 sky130_fd_sc_hd__ha_1 _15696_ (.A(_08100_),
    .B(_08085_),
    .COUT(_08101_),
    .SUM(_08102_));
 sky130_fd_sc_hd__ha_4 _15697_ (.A(_06501_),
    .B(_07928_),
    .COUT(_07982_),
    .SUM(_06498_));
 sky130_fd_sc_hd__ha_1 _15698_ (.A(_06326_),
    .B(_06283_),
    .COUT(_06507_),
    .SUM(_08103_));
 sky130_fd_sc_hd__ha_1 _15699_ (.A(_08102_),
    .B(_08103_),
    .COUT(_06506_),
    .SUM(_08104_));
 sky130_fd_sc_hd__ha_4 _15700_ (.A(_06488_),
    .B(_06510_),
    .COUT(_08105_),
    .SUM(_08106_));
 sky130_fd_sc_hd__ha_1 _15701_ (.A(_08107_),
    .B(_06500_),
    .COUT(_06516_),
    .SUM(_06521_));
 sky130_fd_sc_hd__ha_4 _15702_ (.A(_07928_),
    .B(_06371_),
    .COUT(_06329_),
    .SUM(_08108_));
 sky130_fd_sc_hd__ha_1 _15703_ (.A(_08109_),
    .B(_08108_),
    .COUT(_06523_),
    .SUM(_08110_));
 sky130_fd_sc_hd__ha_1 _15704_ (.A(_08111_),
    .B(_08108_),
    .COUT(_08112_),
    .SUM(_08113_));
 sky130_fd_sc_hd__ha_4 _15705_ (.A(_06519_),
    .B(_06511_),
    .COUT(_08115_),
    .SUM(_08116_));
 sky130_fd_sc_hd__ha_1 _15706_ (.A(_06497_),
    .B(_08117_),
    .COUT(_08114_),
    .SUM(_08118_));
 sky130_fd_sc_hd__ha_1 _15707_ (.A(_08119_),
    .B(_08120_),
    .COUT(_08111_),
    .SUM(_08121_));
 sky130_fd_sc_hd__ha_1 _15708_ (.A(_06520_),
    .B(_08122_),
    .COUT(_08123_),
    .SUM(_08124_));
 sky130_fd_sc_hd__ha_1 _15709_ (.A(_06525_),
    .B(_08125_),
    .COUT(_08122_),
    .SUM(_08126_));
 sky130_fd_sc_hd__ha_1 _15710_ (.A(_08118_),
    .B(_08127_),
    .COUT(_08128_),
    .SUM(_08129_));
 sky130_fd_sc_hd__ha_1 _15711_ (.A(_06371_),
    .B(_08121_),
    .COUT(_08127_),
    .SUM(_08130_));
 sky130_fd_sc_hd__ha_1 _15712_ (.A(_08131_),
    .B(_08132_),
    .COUT(_08133_),
    .SUM(_08134_));
 sky130_fd_sc_hd__ha_1 _15713_ (.A(_08135_),
    .B(_08134_),
    .COUT(_08136_),
    .SUM(_06558_));
 sky130_fd_sc_hd__ha_1 _15714_ (.A(_08137_),
    .B(_06721_),
    .COUT(_08138_),
    .SUM(_08139_));
 sky130_fd_sc_hd__ha_1 _15715_ (.A(_06534_),
    .B(_06646_),
    .COUT(_06559_),
    .SUM(_06593_));
 sky130_fd_sc_hd__ha_1 _15716_ (.A(_08131_),
    .B(_06531_),
    .COUT(_06567_),
    .SUM(_08140_));
 sky130_fd_sc_hd__ha_1 _15717_ (.A(_08141_),
    .B(_08142_),
    .COUT(_08143_),
    .SUM(_06585_));
 sky130_fd_sc_hd__ha_1 _15718_ (.A(_08144_),
    .B(_08145_),
    .COUT(_06586_),
    .SUM(_06622_));
 sky130_fd_sc_hd__ha_1 _15719_ (.A(_06778_),
    .B(net471),
    .COUT(_08147_),
    .SUM(_06618_));
 sky130_fd_sc_hd__ha_1 _15720_ (.A(_08140_),
    .B(_06693_),
    .COUT(_06594_),
    .SUM(_08148_));
 sky130_fd_sc_hd__ha_1 _15721_ (.A(_08149_),
    .B(_08150_),
    .COUT(_06613_),
    .SUM(_08151_));
 sky130_fd_sc_hd__ha_1 _15722_ (.A(_08153_),
    .B(_08154_),
    .COUT(_06623_),
    .SUM(_06681_));
 sky130_fd_sc_hd__ha_1 _15723_ (.A(_06833_),
    .B(_06991_),
    .COUT(_08155_),
    .SUM(_06677_));
 sky130_fd_sc_hd__ha_1 _15724_ (.A(_06986_),
    .B(_08156_),
    .COUT(_08157_),
    .SUM(_08158_));
 sky130_fd_sc_hd__ha_1 _15725_ (.A(_06648_),
    .B(_06943_),
    .COUT(_08159_),
    .SUM(_08160_));
 sky130_fd_sc_hd__ha_1 _15726_ (.A(_08157_),
    .B(_08160_),
    .COUT(_08161_),
    .SUM(_08162_));
 sky130_fd_sc_hd__ha_1 _15727_ (.A(net472),
    .B(_06943_),
    .COUT(_08164_),
    .SUM(_08165_));
 sky130_fd_sc_hd__ha_1 _15728_ (.A(_08158_),
    .B(_08164_),
    .COUT(_08163_),
    .SUM(_08166_));
 sky130_fd_sc_hd__ha_1 _15729_ (.A(_08167_),
    .B(_06695_),
    .COUT(_08168_),
    .SUM(_08169_));
 sky130_fd_sc_hd__ha_1 _15730_ (.A(_08171_),
    .B(_06714_),
    .COUT(_06672_),
    .SUM(_08172_));
 sky130_fd_sc_hd__ha_1 _15731_ (.A(_08131_),
    .B(net466),
    .COUT(_08152_),
    .SUM(_08173_));
 sky130_fd_sc_hd__ha_1 _15732_ (.A(_08174_),
    .B(_08175_),
    .COUT(_06682_),
    .SUM(_06733_));
 sky130_fd_sc_hd__ha_1 _15733_ (.A(_08176_),
    .B(_08166_),
    .COUT(_08170_),
    .SUM(_08177_));
 sky130_fd_sc_hd__ha_1 _15734_ (.A(_06991_),
    .B(_06986_),
    .COUT(_08178_),
    .SUM(_08179_));
 sky130_fd_sc_hd__ha_1 _15735_ (.A(_08178_),
    .B(_08165_),
    .COUT(_08176_),
    .SUM(_08180_));
 sky130_fd_sc_hd__ha_1 _15736_ (.A(_06696_),
    .B(_06747_),
    .COUT(_08181_),
    .SUM(_08182_));
 sky130_fd_sc_hd__ha_1 _15737_ (.A(_08172_),
    .B(_08173_),
    .COUT(_06710_),
    .SUM(_06766_));
 sky130_fd_sc_hd__ha_1 _15738_ (.A(_06715_),
    .B(_08184_),
    .COUT(_06725_),
    .SUM(_08185_));
 sky130_fd_sc_hd__ha_1 _15739_ (.A(_08186_),
    .B(_08187_),
    .COUT(_06734_),
    .SUM(_06782_));
 sky130_fd_sc_hd__ha_1 _15740_ (.A(_08188_),
    .B(_08180_),
    .COUT(_08183_),
    .SUM(_08189_));
 sky130_fd_sc_hd__ha_1 _15741_ (.A(net490),
    .B(net471),
    .COUT(_08190_),
    .SUM(_08191_));
 sky130_fd_sc_hd__ha_1 _15742_ (.A(_08190_),
    .B(_08179_),
    .COUT(_08188_),
    .SUM(_08192_));
 sky130_fd_sc_hd__ha_1 _15743_ (.A(_06748_),
    .B(_06795_),
    .COUT(_08193_),
    .SUM(_08194_));
 sky130_fd_sc_hd__ha_1 _15744_ (.A(_08196_),
    .B(_08181_),
    .COUT(_08197_),
    .SUM(_06757_));
 sky130_fd_sc_hd__ha_1 _15745_ (.A(_06632_),
    .B(_08185_),
    .COUT(_06767_),
    .SUM(_06819_));
 sky130_fd_sc_hd__ha_1 _15746_ (.A(_08131_),
    .B(_06526_),
    .COUT(_08184_),
    .SUM(_08198_));
 sky130_fd_sc_hd__ha_1 _15747_ (.A(_06772_),
    .B(_06826_),
    .COUT(_06785_),
    .SUM(_06821_));
 sky130_fd_sc_hd__ha_1 _15748_ (.A(_08199_),
    .B(_08200_),
    .COUT(_06783_),
    .SUM(_06837_));
 sky130_fd_sc_hd__ha_1 _15749_ (.A(_08201_),
    .B(_08192_),
    .COUT(_08195_),
    .SUM(_08202_));
 sky130_fd_sc_hd__ha_1 _15750_ (.A(_06778_),
    .B(_06991_),
    .COUT(_08203_),
    .SUM(_08204_));
 sky130_fd_sc_hd__ha_1 _15751_ (.A(_08203_),
    .B(_08191_),
    .COUT(_08201_),
    .SUM(_08205_));
 sky130_fd_sc_hd__ha_1 _15752_ (.A(_06796_),
    .B(_06851_),
    .COUT(_08206_),
    .SUM(_08207_));
 sky130_fd_sc_hd__ha_1 _15753_ (.A(_08209_),
    .B(_08193_),
    .COUT(_06805_),
    .SUM(_06810_));
 sky130_fd_sc_hd__ha_1 _15754_ (.A(_06648_),
    .B(_08198_),
    .COUT(_06820_),
    .SUM(_08210_));
 sky130_fd_sc_hd__ha_1 _15755_ (.A(_06827_),
    .B(_06883_),
    .COUT(_08211_),
    .SUM(_08212_));
 sky130_fd_sc_hd__ha_1 _15756_ (.A(_08214_),
    .B(_08215_),
    .COUT(_06838_),
    .SUM(_06891_));
 sky130_fd_sc_hd__ha_1 _15757_ (.A(_06852_),
    .B(_08217_),
    .COUT(_08218_),
    .SUM(_08219_));
 sky130_fd_sc_hd__ha_1 _15758_ (.A(_08220_),
    .B(_08205_),
    .COUT(_08208_),
    .SUM(_08221_));
 sky130_fd_sc_hd__ha_1 _15759_ (.A(_06859_),
    .B(_08206_),
    .COUT(_06862_),
    .SUM(_06867_));
 sky130_fd_sc_hd__ha_1 _15760_ (.A(_06807_),
    .B(_06863_),
    .COUT(_08222_),
    .SUM(_08223_));
 sky130_fd_sc_hd__ha_1 _15761_ (.A(_06884_),
    .B(_08224_),
    .COUT(_08225_),
    .SUM(_08226_));
 sky130_fd_sc_hd__ha_1 _15762_ (.A(_06532_),
    .B(_08156_),
    .COUT(_08213_),
    .SUM(_08227_));
 sky130_fd_sc_hd__ha_1 _15763_ (.A(_06839_),
    .B(_06893_),
    .COUT(_08216_),
    .SUM(_08228_));
 sky130_fd_sc_hd__ha_1 _15764_ (.A(_08229_),
    .B(_08230_),
    .COUT(_06892_),
    .SUM(_06934_));
 sky130_fd_sc_hd__ha_1 _15765_ (.A(_08219_),
    .B(_08221_),
    .COUT(_06858_),
    .SUM(_06906_));
 sky130_fd_sc_hd__ha_1 _15766_ (.A(_08232_),
    .B(_06946_),
    .COUT(_08233_),
    .SUM(_08234_));
 sky130_fd_sc_hd__ha_1 _15767_ (.A(_08235_),
    .B(_08204_),
    .COUT(_08220_),
    .SUM(_08236_));
 sky130_fd_sc_hd__ha_1 _15768_ (.A(_06908_),
    .B(_08218_),
    .COUT(_06911_),
    .SUM(_06916_));
 sky130_fd_sc_hd__ha_1 _15769_ (.A(_06864_),
    .B(_06912_),
    .COUT(_08237_),
    .SUM(_08238_));
 sky130_fd_sc_hd__ha_1 _15770_ (.A(_08226_),
    .B(_08227_),
    .COUT(_06923_),
    .SUM(_06969_));
 sky130_fd_sc_hd__ha_1 _15771_ (.A(_06526_),
    .B(_06532_),
    .COUT(_06930_),
    .SUM(_08239_));
 sky130_fd_sc_hd__ha_1 _15772_ (.A(_08240_),
    .B(_08241_),
    .COUT(_08242_),
    .SUM(_08243_));
 sky130_fd_sc_hd__ha_1 _15773_ (.A(_06894_),
    .B(_06936_),
    .COUT(_08231_),
    .SUM(_08244_));
 sky130_fd_sc_hd__ha_1 _15774_ (.A(_08245_),
    .B(_08246_),
    .COUT(_06935_),
    .SUM(_06977_));
 sky130_fd_sc_hd__ha_1 _15775_ (.A(_08234_),
    .B(_08236_),
    .COUT(_06907_),
    .SUM(_06952_));
 sky130_fd_sc_hd__ha_1 _15776_ (.A(_06947_),
    .B(_06989_),
    .COUT(_08248_),
    .SUM(_08249_));
 sky130_fd_sc_hd__ha_1 _15777_ (.A(net489),
    .B(_06833_),
    .COUT(_08235_),
    .SUM(_08250_));
 sky130_fd_sc_hd__ha_1 _15778_ (.A(_06954_),
    .B(_08233_),
    .COUT(_06957_),
    .SUM(_06962_));
 sky130_fd_sc_hd__ha_1 _15779_ (.A(_06913_),
    .B(_06958_),
    .COUT(_08251_),
    .SUM(_08252_));
 sky130_fd_sc_hd__ha_1 _15780_ (.A(_06943_),
    .B(_08243_),
    .COUT(_06970_),
    .SUM(_07011_));
 sky130_fd_sc_hd__ha_1 _15781_ (.A(_08253_),
    .B(_08239_),
    .COUT(_08241_),
    .SUM(_08254_));
 sky130_fd_sc_hd__ha_1 _15782_ (.A(_08254_),
    .B(_08255_),
    .COUT(_08256_),
    .SUM(_08257_));
 sky130_fd_sc_hd__ha_1 _15783_ (.A(_06937_),
    .B(_06979_),
    .COUT(_08247_),
    .SUM(_08258_));
 sky130_fd_sc_hd__ha_1 _15784_ (.A(_08259_),
    .B(_08260_),
    .COUT(_06978_),
    .SUM(_07017_));
 sky130_fd_sc_hd__ha_1 _15785_ (.A(_08249_),
    .B(_08250_),
    .COUT(_06953_),
    .SUM(_06994_));
 sky130_fd_sc_hd__ha_1 _15786_ (.A(_06778_),
    .B(_06833_),
    .COUT(_07066_),
    .SUM(_07104_));
 sky130_fd_sc_hd__ha_1 _15787_ (.A(_06990_),
    .B(_08262_),
    .COUT(_08263_),
    .SUM(_08264_));
 sky130_fd_sc_hd__ha_1 _15788_ (.A(_06996_),
    .B(_08248_),
    .COUT(_06999_),
    .SUM(_07004_));
 sky130_fd_sc_hd__ha_1 _15789_ (.A(_06959_),
    .B(_07000_),
    .COUT(_08265_),
    .SUM(_08266_));
 sky130_fd_sc_hd__ha_1 _15790_ (.A(_06986_),
    .B(_08257_),
    .COUT(_07012_),
    .SUM(_07043_));
 sky130_fd_sc_hd__ha_1 _15791_ (.A(_06532_),
    .B(_08267_),
    .COUT(_08255_),
    .SUM(_08268_));
 sky130_fd_sc_hd__ha_1 _15792_ (.A(_06980_),
    .B(_07019_),
    .COUT(_08261_),
    .SUM(_08269_));
 sky130_fd_sc_hd__ha_1 _15793_ (.A(_08270_),
    .B(_08271_),
    .COUT(_07018_),
    .SUM(_08272_));
 sky130_fd_sc_hd__ha_1 _15794_ (.A(_08269_),
    .B(_08273_),
    .COUT(_08274_),
    .SUM(_07045_));
 sky130_fd_sc_hd__ha_1 _15795_ (.A(_06778_),
    .B(_08264_),
    .COUT(_06995_),
    .SUM(_08275_));
 sky130_fd_sc_hd__ha_1 _15796_ (.A(net492),
    .B(_07104_),
    .COUT(_08276_),
    .SUM(_08277_));
 sky130_fd_sc_hd__ha_1 _15797_ (.A(_07066_),
    .B(_07026_),
    .COUT(_07088_),
    .SUM(_07093_));
 sky130_fd_sc_hd__ha_1 _15798_ (.A(_08278_),
    .B(_07067_),
    .COUT(_08279_),
    .SUM(_08280_));
 sky130_fd_sc_hd__ha_1 _15799_ (.A(_08282_),
    .B(_08263_),
    .COUT(_07033_),
    .SUM(_07038_));
 sky130_fd_sc_hd__ha_1 _15800_ (.A(_07001_),
    .B(_07034_),
    .COUT(_08283_),
    .SUM(_08284_));
 sky130_fd_sc_hd__ha_1 _15801_ (.A(net473),
    .B(_08268_),
    .COUT(_07044_),
    .SUM(_07062_));
 sky130_fd_sc_hd__ha_1 _15802_ (.A(_07020_),
    .B(_08285_),
    .COUT(_08273_),
    .SUM(_08286_));
 sky130_fd_sc_hd__ha_1 _15803_ (.A(_08288_),
    .B(_08289_),
    .COUT(_08287_),
    .SUM(_08290_));
 sky130_fd_sc_hd__ha_1 _15804_ (.A(_08286_),
    .B(_08291_),
    .COUT(_08292_),
    .SUM(_07064_));
 sky130_fd_sc_hd__ha_1 _15805_ (.A(_06833_),
    .B(_08280_),
    .COUT(_08281_),
    .SUM(_08293_));
 sky130_fd_sc_hd__ha_1 _15806_ (.A(_08292_),
    .B(_08293_),
    .COUT(_08294_),
    .SUM(_07060_));
 sky130_fd_sc_hd__ha_1 _15807_ (.A(_08294_),
    .B(_08279_),
    .COUT(_07053_),
    .SUM(_07057_));
 sky130_fd_sc_hd__ha_1 _15808_ (.A(_07035_),
    .B(_07054_),
    .COUT(_08295_),
    .SUM(_08296_));
 sky130_fd_sc_hd__ha_1 _15809_ (.A(_06991_),
    .B(_07047_),
    .COUT(_07063_),
    .SUM(_07084_));
 sky130_fd_sc_hd__ha_1 _15810_ (.A(_08297_),
    .B(_08298_),
    .COUT(_08291_),
    .SUM(_08299_));
 sky130_fd_sc_hd__ha_1 _15811_ (.A(_08300_),
    .B(_08290_),
    .COUT(_08298_),
    .SUM(_08301_));
 sky130_fd_sc_hd__ha_1 _15812_ (.A(_08302_),
    .B(_08303_),
    .COUT(_08300_),
    .SUM(_08304_));
 sky130_fd_sc_hd__ha_1 _15813_ (.A(_08299_),
    .B(_08305_),
    .COUT(_08306_),
    .SUM(_07086_));
 sky130_fd_sc_hd__ha_1 _15814_ (.A(_08276_),
    .B(_07068_),
    .COUT(_08307_),
    .SUM(_08308_));
 sky130_fd_sc_hd__ha_1 _15815_ (.A(_08306_),
    .B(_08308_),
    .COUT(_08309_),
    .SUM(_08310_));
 sky130_fd_sc_hd__ha_1 _15816_ (.A(_08309_),
    .B(_08307_),
    .COUT(_07075_),
    .SUM(_08311_));
 sky130_fd_sc_hd__ha_1 _15817_ (.A(_07055_),
    .B(_07076_),
    .COUT(_08312_),
    .SUM(_08313_));
 sky130_fd_sc_hd__ha_1 _15818_ (.A(net486),
    .B(_08239_),
    .COUT(_07085_),
    .SUM(_08314_));
 sky130_fd_sc_hd__ha_1 _15819_ (.A(_08301_),
    .B(_08315_),
    .COUT(_08305_),
    .SUM(_08316_));
 sky130_fd_sc_hd__ha_1 _15820_ (.A(_07077_),
    .B(_08318_),
    .COUT(_08319_),
    .SUM(_08320_));
 sky130_fd_sc_hd__ha_1 _15821_ (.A(_07080_),
    .B(_07090_),
    .COUT(_08318_),
    .SUM(_08321_));
 sky130_fd_sc_hd__ha_1 _15822_ (.A(_08322_),
    .B(_08304_),
    .COUT(_08315_),
    .SUM(_08323_));
 sky130_fd_sc_hd__ha_1 _15823_ (.A(_06532_),
    .B(_06778_),
    .COUT(_08317_),
    .SUM(_08324_));
 sky130_fd_sc_hd__ha_1 _15824_ (.A(_08321_),
    .B(_08325_),
    .COUT(_08326_),
    .SUM(_08327_));
 sky130_fd_sc_hd__ha_1 _15825_ (.A(_07091_),
    .B(_08328_),
    .COUT(_08325_),
    .SUM(_08329_));
 sky130_fd_sc_hd__ha_1 _15826_ (.A(_07094_),
    .B(_08330_),
    .COUT(_08328_),
    .SUM(_08331_));
 sky130_fd_sc_hd__ha_1 _15827_ (.A(_08323_),
    .B(_08324_),
    .COUT(_07105_),
    .SUM(_08332_));
 sky130_fd_sc_hd__ha_1 _15828_ (.A(_08333_),
    .B(_08334_),
    .COUT(_08322_),
    .SUM(_08335_));
 sky130_fd_sc_hd__ha_1 _15829_ (.A(_08332_),
    .B(_08336_),
    .COUT(_08337_),
    .SUM(_08338_));
 sky130_fd_sc_hd__dfxtp_1 _15830_ (.D(_00002_),
    .Q(_00011_),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 _15831_ (.D(_00001_),
    .Q(_00010_),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_4 _15832_ (.D(_00000_),
    .Q(_00008_),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 _15833_ (.D(_00020_),
    .Q(_00009_),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_2 _15834_ (.D(_00021_),
    .Q(_00012_),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _15835_ (.D(_00022_),
    .Q(_00016_),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _15836_ (.D(_00023_),
    .Q(_00017_),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__conb_1 _15297__327 (.HI(net385));
 sky130_fd_sc_hd__dfrtp_1 \bit_rev_idx[0]$_DFFE_PN0P_  (.D(_00024_),
    .Q(\bit_rev_idx[0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \bit_rev_idx[1]$_DFFE_PN0P_  (.D(_00025_),
    .Q(\bit_rev_idx[1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \bit_rev_idx[2]$_DFFE_PN0P_  (.D(_00026_),
    .Q(\bit_rev_idx[2] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \busy$_DFFE_PN0P_  (.D(_00027_),
    .Q(net94),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \butterfly_count[0]$_DFFE_PN0P_  (.D(_00028_),
    .Q(\butterfly_count[0] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \butterfly_count[1]$_DFFE_PN0P_  (.D(_00029_),
    .Q(\butterfly_count[1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \butterfly_count[2]$_DFFE_PN0P_  (.D(_00030_),
    .Q(\butterfly_count[2] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \butterfly_in_group[0]$_DFFE_PP_  (.D(_00554_),
    .DE(_00007_),
    .Q(\butterfly_in_group[0] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \butterfly_in_group[1]$_DFFE_PP_  (.D(_00555_),
    .DE(_00007_),
    .Q(\butterfly_in_group[1] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \butterfly_in_group[2]$_DFFE_PP_  (.D(_00556_),
    .DE(_00007_),
    .Q(\butterfly_in_group[2] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[0]$_DFFE_PN0P_  (.D(_00031_),
    .Q(net95),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[100]$_DFFE_PN0P_  (.D(_00032_),
    .Q(net96),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[101]$_DFFE_PN0P_  (.D(_00033_),
    .Q(net97),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[102]$_DFFE_PN0P_  (.D(_00034_),
    .Q(net98),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[103]$_DFFE_PN0P_  (.D(_00035_),
    .Q(net99),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[104]$_DFFE_PN0P_  (.D(_00036_),
    .Q(net100),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[105]$_DFFE_PN0P_  (.D(_00037_),
    .Q(net101),
    .RESET_B(net354),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[106]$_DFFE_PN0P_  (.D(_00038_),
    .Q(net102),
    .RESET_B(net354),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[107]$_DFFE_PN0P_  (.D(_00039_),
    .Q(net103),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[108]$_DFFE_PN0P_  (.D(_00040_),
    .Q(net104),
    .RESET_B(net354),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[109]$_DFFE_PN0P_  (.D(_00041_),
    .Q(net105),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[10]$_DFFE_PN0P_  (.D(_00042_),
    .Q(net106),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[110]$_DFFE_PN0P_  (.D(_00043_),
    .Q(net107),
    .RESET_B(net354),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[111]$_DFFE_PN0P_  (.D(_00044_),
    .Q(net108),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[112]$_DFFE_PN0P_  (.D(_00045_),
    .Q(net109),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[113]$_DFFE_PN0P_  (.D(_00046_),
    .Q(net110),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[114]$_DFFE_PN0P_  (.D(_00047_),
    .Q(net111),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[115]$_DFFE_PN0P_  (.D(_00048_),
    .Q(net112),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[116]$_DFFE_PN0P_  (.D(_00049_),
    .Q(net113),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[117]$_DFFE_PN0P_  (.D(_00050_),
    .Q(net114),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[118]$_DFFE_PN0P_  (.D(_00051_),
    .Q(net115),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[119]$_DFFE_PN0P_  (.D(_00052_),
    .Q(net116),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[11]$_DFFE_PN0P_  (.D(_00053_),
    .Q(net117),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[120]$_DFFE_PN0P_  (.D(_00054_),
    .Q(net118),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[121]$_DFFE_PN0P_  (.D(_00055_),
    .Q(net119),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[122]$_DFFE_PN0P_  (.D(_00056_),
    .Q(net120),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[123]$_DFFE_PN0P_  (.D(_00057_),
    .Q(net121),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[124]$_DFFE_PN0P_  (.D(_00058_),
    .Q(net122),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[125]$_DFFE_PN0P_  (.D(_00059_),
    .Q(net123),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[126]$_DFFE_PN0P_  (.D(_00060_),
    .Q(net124),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[127]$_DFFE_PN0P_  (.D(_00061_),
    .Q(net125),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[12]$_DFFE_PN0P_  (.D(_00062_),
    .Q(net126),
    .RESET_B(net353),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[13]$_DFFE_PN0P_  (.D(_00063_),
    .Q(net127),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[14]$_DFFE_PN0P_  (.D(_00064_),
    .Q(net128),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[15]$_DFFE_PN0P_  (.D(_00065_),
    .Q(net129),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[16]$_DFFE_PN0P_  (.D(_00066_),
    .Q(net130),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[17]$_DFFE_PN0P_  (.D(_00067_),
    .Q(net131),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[18]$_DFFE_PN0P_  (.D(_00068_),
    .Q(net132),
    .RESET_B(net354),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[19]$_DFFE_PN0P_  (.D(_00069_),
    .Q(net133),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[1]$_DFFE_PN0P_  (.D(_00070_),
    .Q(net134),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[20]$_DFFE_PN0P_  (.D(_00071_),
    .Q(net135),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[21]$_DFFE_PN0P_  (.D(_00072_),
    .Q(net136),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[22]$_DFFE_PN0P_  (.D(_00073_),
    .Q(net137),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[23]$_DFFE_PN0P_  (.D(_00074_),
    .Q(net138),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[24]$_DFFE_PN0P_  (.D(_00075_),
    .Q(net139),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[25]$_DFFE_PN0P_  (.D(_00076_),
    .Q(net140),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[26]$_DFFE_PN0P_  (.D(_00077_),
    .Q(net141),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[27]$_DFFE_PN0P_  (.D(_00078_),
    .Q(net142),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[28]$_DFFE_PN0P_  (.D(_00079_),
    .Q(net143),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[29]$_DFFE_PN0P_  (.D(_00080_),
    .Q(net144),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[2]$_DFFE_PN0P_  (.D(_00081_),
    .Q(net145),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[30]$_DFFE_PN0P_  (.D(_00082_),
    .Q(net146),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[31]$_DFFE_PN0P_  (.D(_00083_),
    .Q(net147),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[32]$_DFFE_PN0P_  (.D(_00084_),
    .Q(net148),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[33]$_DFFE_PN0P_  (.D(_00085_),
    .Q(net149),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[34]$_DFFE_PN0P_  (.D(_00086_),
    .Q(net150),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[35]$_DFFE_PN0P_  (.D(_00087_),
    .Q(net151),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[36]$_DFFE_PN0P_  (.D(_00088_),
    .Q(net152),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[37]$_DFFE_PN0P_  (.D(_00089_),
    .Q(net153),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[38]$_DFFE_PN0P_  (.D(_00090_),
    .Q(net154),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[39]$_DFFE_PN0P_  (.D(_00091_),
    .Q(net155),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[3]$_DFFE_PN0P_  (.D(_00092_),
    .Q(net156),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[40]$_DFFE_PN0P_  (.D(_00093_),
    .Q(net157),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[41]$_DFFE_PN0P_  (.D(_00094_),
    .Q(net158),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[42]$_DFFE_PN0P_  (.D(_00095_),
    .Q(net159),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[43]$_DFFE_PN0P_  (.D(_00096_),
    .Q(net160),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[44]$_DFFE_PN0P_  (.D(_00097_),
    .Q(net161),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[45]$_DFFE_PN0P_  (.D(_00098_),
    .Q(net162),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[46]$_DFFE_PN0P_  (.D(_00099_),
    .Q(net163),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[47]$_DFFE_PN0P_  (.D(_00100_),
    .Q(net164),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[48]$_DFFE_PN0P_  (.D(_00101_),
    .Q(net165),
    .RESET_B(net353),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[49]$_DFFE_PN0P_  (.D(_00102_),
    .Q(net166),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[4]$_DFFE_PN0P_  (.D(_00103_),
    .Q(net167),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[50]$_DFFE_PN0P_  (.D(_00104_),
    .Q(net168),
    .RESET_B(net353),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[51]$_DFFE_PN0P_  (.D(_00105_),
    .Q(net169),
    .RESET_B(net353),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[52]$_DFFE_PN0P_  (.D(_00106_),
    .Q(net170),
    .RESET_B(net353),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[53]$_DFFE_PN0P_  (.D(_00107_),
    .Q(net171),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[54]$_DFFE_PN0P_  (.D(_00108_),
    .Q(net172),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[55]$_DFFE_PN0P_  (.D(_00109_),
    .Q(net173),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[56]$_DFFE_PN0P_  (.D(_00110_),
    .Q(net174),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[57]$_DFFE_PN0P_  (.D(_00111_),
    .Q(net175),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[58]$_DFFE_PN0P_  (.D(_00112_),
    .Q(net176),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[59]$_DFFE_PN0P_  (.D(_00113_),
    .Q(net177),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[5]$_DFFE_PN0P_  (.D(_00114_),
    .Q(net178),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[60]$_DFFE_PN0P_  (.D(_00115_),
    .Q(net179),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[61]$_DFFE_PN0P_  (.D(_00116_),
    .Q(net180),
    .RESET_B(net353),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[62]$_DFFE_PN0P_  (.D(_00117_),
    .Q(net181),
    .RESET_B(net355),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[63]$_DFFE_PN0P_  (.D(_00118_),
    .Q(net182),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[64]$_DFFE_PN0P_  (.D(_00119_),
    .Q(net183),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[65]$_DFFE_PN0P_  (.D(_00120_),
    .Q(net184),
    .RESET_B(net356),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[66]$_DFFE_PN0P_  (.D(_00121_),
    .Q(net185),
    .RESET_B(net356),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[67]$_DFFE_PN0P_  (.D(_00122_),
    .Q(net186),
    .RESET_B(net356),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[68]$_DFFE_PN0P_  (.D(_00123_),
    .Q(net187),
    .RESET_B(net356),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[69]$_DFFE_PN0P_  (.D(_00124_),
    .Q(net188),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[6]$_DFFE_PN0P_  (.D(_00125_),
    .Q(net189),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[70]$_DFFE_PN0P_  (.D(_00126_),
    .Q(net190),
    .RESET_B(net356),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[71]$_DFFE_PN0P_  (.D(_00127_),
    .Q(net191),
    .RESET_B(net356),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[72]$_DFFE_PN0P_  (.D(_00128_),
    .Q(net192),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[73]$_DFFE_PN0P_  (.D(_00129_),
    .Q(net193),
    .RESET_B(net356),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[74]$_DFFE_PN0P_  (.D(_00130_),
    .Q(net194),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[75]$_DFFE_PN0P_  (.D(_00131_),
    .Q(net195),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[76]$_DFFE_PN0P_  (.D(_00132_),
    .Q(net196),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[77]$_DFFE_PN0P_  (.D(_00133_),
    .Q(net197),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[78]$_DFFE_PN0P_  (.D(_00134_),
    .Q(net198),
    .RESET_B(net356),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[79]$_DFFE_PN0P_  (.D(_00135_),
    .Q(net199),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[7]$_DFFE_PN0P_  (.D(_00136_),
    .Q(net200),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[80]$_DFFE_PN0P_  (.D(_00137_),
    .Q(net201),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[81]$_DFFE_PN0P_  (.D(_00138_),
    .Q(net202),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[82]$_DFFE_PN0P_  (.D(_00139_),
    .Q(net203),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[83]$_DFFE_PN0P_  (.D(_00140_),
    .Q(net204),
    .RESET_B(net355),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[84]$_DFFE_PN0P_  (.D(_00141_),
    .Q(net205),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[85]$_DFFE_PN0P_  (.D(_00142_),
    .Q(net206),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[86]$_DFFE_PN0P_  (.D(_00143_),
    .Q(net207),
    .RESET_B(net355),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[87]$_DFFE_PN0P_  (.D(_00144_),
    .Q(net208),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[88]$_DFFE_PN0P_  (.D(_00145_),
    .Q(net209),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[89]$_DFFE_PN0P_  (.D(_00146_),
    .Q(net210),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[8]$_DFFE_PN0P_  (.D(_00147_),
    .Q(net211),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[90]$_DFFE_PN0P_  (.D(_00148_),
    .Q(net212),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[91]$_DFFE_PN0P_  (.D(_00149_),
    .Q(net213),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[92]$_DFFE_PN0P_  (.D(_00150_),
    .Q(net214),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \data_out_imag[93]$_DFFE_PN0P_  (.D(_00151_),
    .Q(net215),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[94]$_DFFE_PN0P_  (.D(_00152_),
    .Q(net216),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[95]$_DFFE_PN0P_  (.D(_00153_),
    .Q(net217),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[96]$_DFFE_PN0P_  (.D(_00154_),
    .Q(net218),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[97]$_DFFE_PN0P_  (.D(_00155_),
    .Q(net219),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_imag[98]$_DFFE_PN0P_  (.D(_00156_),
    .Q(net220),
    .RESET_B(net353),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[99]$_DFFE_PN0P_  (.D(_00157_),
    .Q(net221),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_imag[9]$_DFFE_PN0P_  (.D(_00158_),
    .Q(net222),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[0]$_DFFE_PN0P_  (.D(_00159_),
    .Q(net223),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[100]$_DFFE_PN0P_  (.D(_00160_),
    .Q(net224),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[101]$_DFFE_PN0P_  (.D(_00161_),
    .Q(net225),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[102]$_DFFE_PN0P_  (.D(_00162_),
    .Q(net226),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[103]$_DFFE_PN0P_  (.D(_00163_),
    .Q(net227),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[104]$_DFFE_PN0P_  (.D(_00164_),
    .Q(net228),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[105]$_DFFE_PN0P_  (.D(_00165_),
    .Q(net229),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[106]$_DFFE_PN0P_  (.D(_00166_),
    .Q(net230),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[107]$_DFFE_PN0P_  (.D(_00167_),
    .Q(net231),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[108]$_DFFE_PN0P_  (.D(_00168_),
    .Q(net232),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[109]$_DFFE_PN0P_  (.D(_00169_),
    .Q(net233),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[10]$_DFFE_PN0P_  (.D(_00170_),
    .Q(net234),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[110]$_DFFE_PN0P_  (.D(_00171_),
    .Q(net235),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[111]$_DFFE_PN0P_  (.D(_00172_),
    .Q(net236),
    .RESET_B(net356),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[112]$_DFFE_PN0P_  (.D(_00173_),
    .Q(net237),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[113]$_DFFE_PN0P_  (.D(_00174_),
    .Q(net238),
    .RESET_B(net356),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[114]$_DFFE_PN0P_  (.D(_00175_),
    .Q(net239),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[115]$_DFFE_PN0P_  (.D(_00176_),
    .Q(net240),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[116]$_DFFE_PN0P_  (.D(_00177_),
    .Q(net241),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[117]$_DFFE_PN0P_  (.D(_00178_),
    .Q(net242),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[118]$_DFFE_PN0P_  (.D(_00179_),
    .Q(net243),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[119]$_DFFE_PN0P_  (.D(_00180_),
    .Q(net244),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[11]$_DFFE_PN0P_  (.D(_00181_),
    .Q(net245),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[120]$_DFFE_PN0P_  (.D(_00182_),
    .Q(net246),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[121]$_DFFE_PN0P_  (.D(_00183_),
    .Q(net247),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[122]$_DFFE_PN0P_  (.D(_00184_),
    .Q(net248),
    .RESET_B(net356),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[123]$_DFFE_PN0P_  (.D(_00185_),
    .Q(net249),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[124]$_DFFE_PN0P_  (.D(_00186_),
    .Q(net250),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[125]$_DFFE_PN0P_  (.D(_00187_),
    .Q(net251),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[126]$_DFFE_PN0P_  (.D(_00188_),
    .Q(net252),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[127]$_DFFE_PN0P_  (.D(_00189_),
    .Q(net253),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[12]$_DFFE_PN0P_  (.D(_00190_),
    .Q(net254),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[13]$_DFFE_PN0P_  (.D(_00191_),
    .Q(net255),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[14]$_DFFE_PN0P_  (.D(_00192_),
    .Q(net256),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[15]$_DFFE_PN0P_  (.D(_00193_),
    .Q(net257),
    .RESET_B(net353),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[16]$_DFFE_PN0P_  (.D(_00194_),
    .Q(net258),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[17]$_DFFE_PN0P_  (.D(_00195_),
    .Q(net259),
    .RESET_B(net353),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[18]$_DFFE_PN0P_  (.D(_00196_),
    .Q(net260),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[19]$_DFFE_PN0P_  (.D(_00197_),
    .Q(net261),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[1]$_DFFE_PN0P_  (.D(_00198_),
    .Q(net262),
    .RESET_B(net354),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[20]$_DFFE_PN0P_  (.D(_00199_),
    .Q(net263),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[21]$_DFFE_PN0P_  (.D(_00200_),
    .Q(net264),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[22]$_DFFE_PN0P_  (.D(_00201_),
    .Q(net265),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[23]$_DFFE_PN0P_  (.D(_00202_),
    .Q(net266),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[24]$_DFFE_PN0P_  (.D(_00203_),
    .Q(net267),
    .RESET_B(net354),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[25]$_DFFE_PN0P_  (.D(_00204_),
    .Q(net268),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[26]$_DFFE_PN0P_  (.D(_00205_),
    .Q(net269),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[27]$_DFFE_PN0P_  (.D(_00206_),
    .Q(net270),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[28]$_DFFE_PN0P_  (.D(_00207_),
    .Q(net271),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[29]$_DFFE_PN0P_  (.D(_00208_),
    .Q(net272),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[2]$_DFFE_PN0P_  (.D(_00209_),
    .Q(net273),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[30]$_DFFE_PN0P_  (.D(_00210_),
    .Q(net274),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[31]$_DFFE_PN0P_  (.D(_00211_),
    .Q(net275),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_2 \data_out_real[32]$_DFFE_PN0P_  (.D(_00212_),
    .Q(net276),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[33]$_DFFE_PN0P_  (.D(_00213_),
    .Q(net277),
    .RESET_B(net92),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[34]$_DFFE_PN0P_  (.D(_00214_),
    .Q(net278),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[35]$_DFFE_PN0P_  (.D(_00215_),
    .Q(net279),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[36]$_DFFE_PN0P_  (.D(_00216_),
    .Q(net280),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[37]$_DFFE_PN0P_  (.D(_00217_),
    .Q(net281),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[38]$_DFFE_PN0P_  (.D(_00218_),
    .Q(net282),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[39]$_DFFE_PN0P_  (.D(_00219_),
    .Q(net283),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[3]$_DFFE_PN0P_  (.D(_00220_),
    .Q(net284),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[40]$_DFFE_PN0P_  (.D(_00221_),
    .Q(net285),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[41]$_DFFE_PN0P_  (.D(_00222_),
    .Q(net286),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[42]$_DFFE_PN0P_  (.D(_00223_),
    .Q(net287),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[43]$_DFFE_PN0P_  (.D(_00224_),
    .Q(net288),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[44]$_DFFE_PN0P_  (.D(_00225_),
    .Q(net289),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[45]$_DFFE_PN0P_  (.D(_00226_),
    .Q(net290),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[46]$_DFFE_PN0P_  (.D(_00227_),
    .Q(net291),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[47]$_DFFE_PN0P_  (.D(_00228_),
    .Q(net292),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[48]$_DFFE_PN0P_  (.D(_00229_),
    .Q(net293),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[49]$_DFFE_PN0P_  (.D(_00230_),
    .Q(net294),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[4]$_DFFE_PN0P_  (.D(_00231_),
    .Q(net295),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[50]$_DFFE_PN0P_  (.D(_00232_),
    .Q(net296),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[51]$_DFFE_PN0P_  (.D(_00233_),
    .Q(net297),
    .RESET_B(net92),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[52]$_DFFE_PN0P_  (.D(_00234_),
    .Q(net298),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[53]$_DFFE_PN0P_  (.D(_00235_),
    .Q(net299),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[54]$_DFFE_PN0P_  (.D(_00236_),
    .Q(net300),
    .RESET_B(net92),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[55]$_DFFE_PN0P_  (.D(_00237_),
    .Q(net301),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[56]$_DFFE_PN0P_  (.D(_00238_),
    .Q(net302),
    .RESET_B(net354),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[57]$_DFFE_PN0P_  (.D(_00239_),
    .Q(net303),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[58]$_DFFE_PN0P_  (.D(_00240_),
    .Q(net304),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[59]$_DFFE_PN0P_  (.D(_00241_),
    .Q(net305),
    .RESET_B(net357),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[5]$_DFFE_PN0P_  (.D(_00242_),
    .Q(net306),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[60]$_DFFE_PN0P_  (.D(_00243_),
    .Q(net307),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[61]$_DFFE_PN0P_  (.D(_00244_),
    .Q(net308),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[62]$_DFFE_PN0P_  (.D(_00245_),
    .Q(net309),
    .RESET_B(net92),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[63]$_DFFE_PN0P_  (.D(_00246_),
    .Q(net310),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[64]$_DFFE_PN0P_  (.D(_00247_),
    .Q(net311),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[65]$_DFFE_PN0P_  (.D(_00248_),
    .Q(net312),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[66]$_DFFE_PN0P_  (.D(_00249_),
    .Q(net313),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[67]$_DFFE_PN0P_  (.D(_00250_),
    .Q(net314),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[68]$_DFFE_PN0P_  (.D(_00251_),
    .Q(net315),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[69]$_DFFE_PN0P_  (.D(_00252_),
    .Q(net316),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[6]$_DFFE_PN0P_  (.D(_00253_),
    .Q(net317),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[70]$_DFFE_PN0P_  (.D(_00254_),
    .Q(net318),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[71]$_DFFE_PN0P_  (.D(_00255_),
    .Q(net319),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[72]$_DFFE_PN0P_  (.D(_00256_),
    .Q(net320),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[73]$_DFFE_PN0P_  (.D(_00257_),
    .Q(net321),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[74]$_DFFE_PN0P_  (.D(_00258_),
    .Q(net322),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[75]$_DFFE_PN0P_  (.D(_00259_),
    .Q(net323),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[76]$_DFFE_PN0P_  (.D(_00260_),
    .Q(net324),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[77]$_DFFE_PN0P_  (.D(_00261_),
    .Q(net325),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[78]$_DFFE_PN0P_  (.D(_00262_),
    .Q(net326),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[79]$_DFFE_PN0P_  (.D(_00263_),
    .Q(net327),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[7]$_DFFE_PN0P_  (.D(_00264_),
    .Q(net328),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[80]$_DFFE_PN0P_  (.D(_00265_),
    .Q(net329),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[81]$_DFFE_PN0P_  (.D(_00266_),
    .Q(net330),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[82]$_DFFE_PN0P_  (.D(_00267_),
    .Q(net331),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[83]$_DFFE_PN0P_  (.D(_00268_),
    .Q(net332),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[84]$_DFFE_PN0P_  (.D(_00269_),
    .Q(net333),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[85]$_DFFE_PN0P_  (.D(_00270_),
    .Q(net334),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[86]$_DFFE_PN0P_  (.D(_00271_),
    .Q(net335),
    .RESET_B(net356),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[87]$_DFFE_PN0P_  (.D(_00272_),
    .Q(net336),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[88]$_DFFE_PN0P_  (.D(_00273_),
    .Q(net337),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[89]$_DFFE_PN0P_  (.D(_00274_),
    .Q(net338),
    .RESET_B(net356),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[8]$_DFFE_PN0P_  (.D(_00275_),
    .Q(net339),
    .RESET_B(net356),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[90]$_DFFE_PN0P_  (.D(_00276_),
    .Q(net340),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[91]$_DFFE_PN0P_  (.D(_00277_),
    .Q(net341),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[92]$_DFFE_PN0P_  (.D(_00278_),
    .Q(net342),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[93]$_DFFE_PN0P_  (.D(_00279_),
    .Q(net343),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[94]$_DFFE_PN0P_  (.D(_00280_),
    .Q(net344),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[95]$_DFFE_PN0P_  (.D(_00281_),
    .Q(net345),
    .RESET_B(net356),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[96]$_DFFE_PN0P_  (.D(_00282_),
    .Q(net346),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[97]$_DFFE_PN0P_  (.D(_00283_),
    .Q(net347),
    .RESET_B(net355),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[98]$_DFFE_PN0P_  (.D(_00284_),
    .Q(net348),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[99]$_DFFE_PN0P_  (.D(_00285_),
    .Q(net349),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out_real[9]$_DFFE_PN0P_  (.D(_00286_),
    .Q(net350),
    .RESET_B(net356),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfstp_1 \data_ready$_DFFE_PN1P_  (.D(_00287_),
    .Q(net351),
    .SET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_valid_out$_DFFE_PN0P_  (.D(_00288_),
    .Q(net352),
    .RESET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \group[0]$_DFFE_PP_  (.D(_00551_),
    .DE(_00007_),
    .Q(\group[0] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \group[1]$_DFFE_PP_  (.D(net35),
    .DE(_00007_),
    .Q(\group[1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \group[2]$_DFFE_PP_  (.D(net434),
    .DE(_00007_),
    .Q(\group[2] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx1[0]$_DFFE_PP_  (.D(_05879_),
    .DE(_00007_),
    .Q(\idx1[0] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx1[1]$_DFFE_PP_  (.D(_05880_),
    .DE(_00007_),
    .Q(\idx1[1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx1[2]$_DFFE_PP_  (.D(_00013_),
    .DE(_00007_),
    .Q(\idx1[2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx2[0]$_DFFE_PP_  (.D(_05881_),
    .DE(_00007_),
    .Q(\idx2[0] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx2[1]$_DFFE_PP_  (.D(_00014_),
    .DE(_00007_),
    .Q(\idx2[1] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \idx2[2]$_DFFE_PP_  (.D(_00015_),
    .DE(_00007_),
    .Q(\idx2[2] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \sample_count[0]$_DFFE_PN0P_  (.D(_00289_),
    .Q(\sample_count[0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \sample_count[1]$_DFFE_PN0P_  (.D(_00290_),
    .Q(\sample_count[1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \sample_count[2]$_DFFE_PN0P_  (.D(_00291_),
    .Q(\sample_count[2] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][0]$_DFFE_PN0P_  (.D(_00292_),
    .Q(\samples_imag[0][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][10]$_DFFE_PN0P_  (.D(_00293_),
    .Q(\samples_imag[0][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][11]$_DFFE_PN0P_  (.D(_00294_),
    .Q(\samples_imag[0][11] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][12]$_DFFE_PN0P_  (.D(_00295_),
    .Q(\samples_imag[0][12] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[0][13]$_DFFE_PN0P_  (.D(_00296_),
    .Q(\samples_imag[0][13] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[0][14]$_DFFE_PN0P_  (.D(_00297_),
    .Q(\samples_imag[0][14] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][15]$_DFFE_PN0P_  (.D(_00298_),
    .Q(\samples_imag[0][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][1]$_DFFE_PN0P_  (.D(_00299_),
    .Q(\samples_imag[0][1] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][2]$_DFFE_PN0P_  (.D(_00300_),
    .Q(\samples_imag[0][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][3]$_DFFE_PN0P_  (.D(_00301_),
    .Q(\samples_imag[0][3] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][4]$_DFFE_PN0P_  (.D(_00302_),
    .Q(\samples_imag[0][4] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][5]$_DFFE_PN0P_  (.D(_00303_),
    .Q(\samples_imag[0][5] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][6]$_DFFE_PN0P_  (.D(_00304_),
    .Q(\samples_imag[0][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][7]$_DFFE_PN0P_  (.D(_00305_),
    .Q(\samples_imag[0][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][8]$_DFFE_PN0P_  (.D(_00306_),
    .Q(\samples_imag[0][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[0][9]$_DFFE_PN0P_  (.D(_00307_),
    .Q(\samples_imag[0][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][0]$_DFFE_PN0P_  (.D(_00308_),
    .Q(\samples_imag[1][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[1][10]$_DFFE_PN0P_  (.D(_00309_),
    .Q(\samples_imag[1][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[1][11]$_DFFE_PN0P_  (.D(_00310_),
    .Q(\samples_imag[1][11] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][12]$_DFFE_PN0P_  (.D(_00311_),
    .Q(\samples_imag[1][12] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[1][13]$_DFFE_PN0P_  (.D(_00312_),
    .Q(\samples_imag[1][13] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][14]$_DFFE_PN0P_  (.D(_00313_),
    .Q(\samples_imag[1][14] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][15]$_DFFE_PN0P_  (.D(_00314_),
    .Q(\samples_imag[1][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \samples_imag[1][1]$_DFFE_PN0P_  (.D(_00315_),
    .Q(\samples_imag[1][1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][2]$_DFFE_PN0P_  (.D(_00316_),
    .Q(\samples_imag[1][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][3]$_DFFE_PN0P_  (.D(_00317_),
    .Q(\samples_imag[1][3] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \samples_imag[1][4]$_DFFE_PN0P_  (.D(_00318_),
    .Q(\samples_imag[1][4] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][5]$_DFFE_PN0P_  (.D(_00319_),
    .Q(\samples_imag[1][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][6]$_DFFE_PN0P_  (.D(_00320_),
    .Q(\samples_imag[1][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][7]$_DFFE_PN0P_  (.D(_00321_),
    .Q(\samples_imag[1][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][8]$_DFFE_PN0P_  (.D(_00322_),
    .Q(\samples_imag[1][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[1][9]$_DFFE_PN0P_  (.D(_00323_),
    .Q(\samples_imag[1][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][0]$_DFFE_PN0P_  (.D(_00324_),
    .Q(\samples_imag[2][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][10]$_DFFE_PN0P_  (.D(_00325_),
    .Q(\samples_imag[2][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][11]$_DFFE_PN0P_  (.D(_00326_),
    .Q(\samples_imag[2][11] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][12]$_DFFE_PN0P_  (.D(_00327_),
    .Q(\samples_imag[2][12] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[2][13]$_DFFE_PN0P_  (.D(_00328_),
    .Q(\samples_imag[2][13] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][14]$_DFFE_PN0P_  (.D(_00329_),
    .Q(\samples_imag[2][14] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][15]$_DFFE_PN0P_  (.D(_00330_),
    .Q(\samples_imag[2][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][1]$_DFFE_PN0P_  (.D(_00331_),
    .Q(\samples_imag[2][1] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][2]$_DFFE_PN0P_  (.D(_00332_),
    .Q(\samples_imag[2][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][3]$_DFFE_PN0P_  (.D(_00333_),
    .Q(\samples_imag[2][3] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][4]$_DFFE_PN0P_  (.D(_00334_),
    .Q(\samples_imag[2][4] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][5]$_DFFE_PN0P_  (.D(_00335_),
    .Q(\samples_imag[2][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][6]$_DFFE_PN0P_  (.D(_00336_),
    .Q(\samples_imag[2][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][7]$_DFFE_PN0P_  (.D(_00337_),
    .Q(\samples_imag[2][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][8]$_DFFE_PN0P_  (.D(_00338_),
    .Q(\samples_imag[2][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[2][9]$_DFFE_PN0P_  (.D(_00339_),
    .Q(\samples_imag[2][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][0]$_DFFE_PN0P_  (.D(_00340_),
    .Q(\samples_imag[3][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][10]$_DFFE_PN0P_  (.D(_00341_),
    .Q(\samples_imag[3][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][11]$_DFFE_PN0P_  (.D(_00342_),
    .Q(\samples_imag[3][11] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][12]$_DFFE_PN0P_  (.D(_00343_),
    .Q(\samples_imag[3][12] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][13]$_DFFE_PN0P_  (.D(_00344_),
    .Q(\samples_imag[3][13] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][14]$_DFFE_PN0P_  (.D(_00345_),
    .Q(\samples_imag[3][14] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][15]$_DFFE_PN0P_  (.D(_00346_),
    .Q(\samples_imag[3][15] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][1]$_DFFE_PN0P_  (.D(_00347_),
    .Q(\samples_imag[3][1] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][2]$_DFFE_PN0P_  (.D(_00348_),
    .Q(\samples_imag[3][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][3]$_DFFE_PN0P_  (.D(_00349_),
    .Q(\samples_imag[3][3] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][4]$_DFFE_PN0P_  (.D(_00350_),
    .Q(\samples_imag[3][4] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][5]$_DFFE_PN0P_  (.D(_00351_),
    .Q(\samples_imag[3][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][6]$_DFFE_PN0P_  (.D(_00352_),
    .Q(\samples_imag[3][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][7]$_DFFE_PN0P_  (.D(_00353_),
    .Q(\samples_imag[3][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][8]$_DFFE_PN0P_  (.D(_00354_),
    .Q(\samples_imag[3][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[3][9]$_DFFE_PN0P_  (.D(_00355_),
    .Q(\samples_imag[3][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][0]$_DFFE_PN0P_  (.D(_00356_),
    .Q(\samples_imag[4][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][10]$_DFFE_PN0P_  (.D(_00357_),
    .Q(\samples_imag[4][10] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][11]$_DFFE_PN0P_  (.D(_00358_),
    .Q(\samples_imag[4][11] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[4][12]$_DFFE_PN0P_  (.D(_00359_),
    .Q(\samples_imag[4][12] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][13]$_DFFE_PN0P_  (.D(_00360_),
    .Q(\samples_imag[4][13] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][14]$_DFFE_PN0P_  (.D(_00361_),
    .Q(\samples_imag[4][14] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][15]$_DFFE_PN0P_  (.D(_00362_),
    .Q(\samples_imag[4][15] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][1]$_DFFE_PN0P_  (.D(_00363_),
    .Q(\samples_imag[4][1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][2]$_DFFE_PN0P_  (.D(_00364_),
    .Q(\samples_imag[4][2] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[4][3]$_DFFE_PN0P_  (.D(_00365_),
    .Q(\samples_imag[4][3] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][4]$_DFFE_PN0P_  (.D(_00366_),
    .Q(\samples_imag[4][4] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][5]$_DFFE_PN0P_  (.D(_00367_),
    .Q(\samples_imag[4][5] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][6]$_DFFE_PN0P_  (.D(_00368_),
    .Q(\samples_imag[4][6] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[4][7]$_DFFE_PN0P_  (.D(_00369_),
    .Q(\samples_imag[4][7] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][8]$_DFFE_PN0P_  (.D(_00370_),
    .Q(\samples_imag[4][8] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[4][9]$_DFFE_PN0P_  (.D(_00371_),
    .Q(\samples_imag[4][9] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][0]$_DFFE_PN0P_  (.D(_00372_),
    .Q(\samples_imag[5][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][10]$_DFFE_PN0P_  (.D(_00373_),
    .Q(\samples_imag[5][10] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][11]$_DFFE_PN0P_  (.D(_00374_),
    .Q(\samples_imag[5][11] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][12]$_DFFE_PN0P_  (.D(_00375_),
    .Q(\samples_imag[5][12] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][13]$_DFFE_PN0P_  (.D(_00376_),
    .Q(\samples_imag[5][13] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][14]$_DFFE_PN0P_  (.D(_00377_),
    .Q(\samples_imag[5][14] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][15]$_DFFE_PN0P_  (.D(_00378_),
    .Q(\samples_imag[5][15] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][1]$_DFFE_PN0P_  (.D(_00379_),
    .Q(\samples_imag[5][1] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][2]$_DFFE_PN0P_  (.D(_00380_),
    .Q(\samples_imag[5][2] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][3]$_DFFE_PN0P_  (.D(_00381_),
    .Q(\samples_imag[5][3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[5][4]$_DFFE_PN0P_  (.D(_00382_),
    .Q(\samples_imag[5][4] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][5]$_DFFE_PN0P_  (.D(_00383_),
    .Q(\samples_imag[5][5] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[5][6]$_DFFE_PN0P_  (.D(_00384_),
    .Q(\samples_imag[5][6] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[5][7]$_DFFE_PN0P_  (.D(_00385_),
    .Q(\samples_imag[5][7] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[5][8]$_DFFE_PN0P_  (.D(_00386_),
    .Q(\samples_imag[5][8] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[5][9]$_DFFE_PN0P_  (.D(_00387_),
    .Q(\samples_imag[5][9] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][0]$_DFFE_PN0P_  (.D(_00388_),
    .Q(\samples_imag[6][0] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][10]$_DFFE_PN0P_  (.D(_00389_),
    .Q(\samples_imag[6][10] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][11]$_DFFE_PN0P_  (.D(_00390_),
    .Q(\samples_imag[6][11] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][12]$_DFFE_PN0P_  (.D(_00391_),
    .Q(\samples_imag[6][12] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][13]$_DFFE_PN0P_  (.D(_00392_),
    .Q(\samples_imag[6][13] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][14]$_DFFE_PN0P_  (.D(_00393_),
    .Q(\samples_imag[6][14] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[6][15]$_DFFE_PN0P_  (.D(_00394_),
    .Q(\samples_imag[6][15] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][1]$_DFFE_PN0P_  (.D(_00395_),
    .Q(\samples_imag[6][1] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][2]$_DFFE_PN0P_  (.D(_00396_),
    .Q(\samples_imag[6][2] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][3]$_DFFE_PN0P_  (.D(_00397_),
    .Q(\samples_imag[6][3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][4]$_DFFE_PN0P_  (.D(_00398_),
    .Q(\samples_imag[6][4] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][5]$_DFFE_PN0P_  (.D(_00399_),
    .Q(\samples_imag[6][5] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][6]$_DFFE_PN0P_  (.D(_00400_),
    .Q(\samples_imag[6][6] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][7]$_DFFE_PN0P_  (.D(_00401_),
    .Q(\samples_imag[6][7] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][8]$_DFFE_PN0P_  (.D(_00402_),
    .Q(\samples_imag[6][8] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[6][9]$_DFFE_PN0P_  (.D(_00403_),
    .Q(\samples_imag[6][9] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][0]$_DFFE_PN0P_  (.D(_00404_),
    .Q(\samples_imag[7][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][10]$_DFFE_PN0P_  (.D(_00405_),
    .Q(\samples_imag[7][10] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][11]$_DFFE_PN0P_  (.D(_00406_),
    .Q(\samples_imag[7][11] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][12]$_DFFE_PN0P_  (.D(_00407_),
    .Q(\samples_imag[7][12] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][13]$_DFFE_PN0P_  (.D(_00408_),
    .Q(\samples_imag[7][13] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][14]$_DFFE_PN0P_  (.D(_00409_),
    .Q(\samples_imag[7][14] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][15]$_DFFE_PN0P_  (.D(_00410_),
    .Q(\samples_imag[7][15] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][1]$_DFFE_PN0P_  (.D(_00411_),
    .Q(\samples_imag[7][1] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][2]$_DFFE_PN0P_  (.D(_00412_),
    .Q(\samples_imag[7][2] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][3]$_DFFE_PN0P_  (.D(_00413_),
    .Q(\samples_imag[7][3] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][4]$_DFFE_PN0P_  (.D(_00414_),
    .Q(\samples_imag[7][4] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][5]$_DFFE_PN0P_  (.D(_00415_),
    .Q(\samples_imag[7][5] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][6]$_DFFE_PN0P_  (.D(_00416_),
    .Q(\samples_imag[7][6] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[7][7]$_DFFE_PN0P_  (.D(_00417_),
    .Q(\samples_imag[7][7] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_imag[7][8]$_DFFE_PN0P_  (.D(_00418_),
    .Q(\samples_imag[7][8] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_imag[7][9]$_DFFE_PN0P_  (.D(_00419_),
    .Q(\samples_imag[7][9] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][0]$_DFFE_PN0P_  (.D(_00420_),
    .Q(\samples_real[0][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][10]$_DFFE_PN0P_  (.D(_00421_),
    .Q(\samples_real[0][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][11]$_DFFE_PN0P_  (.D(_00422_),
    .Q(\samples_real[0][11] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][12]$_DFFE_PN0P_  (.D(_00423_),
    .Q(\samples_real[0][12] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][13]$_DFFE_PN0P_  (.D(_00424_),
    .Q(\samples_real[0][13] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][14]$_DFFE_PN0P_  (.D(_00425_),
    .Q(\samples_real[0][14] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][15]$_DFFE_PN0P_  (.D(_00426_),
    .Q(\samples_real[0][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][1]$_DFFE_PN0P_  (.D(_00427_),
    .Q(\samples_real[0][1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][2]$_DFFE_PN0P_  (.D(_00428_),
    .Q(\samples_real[0][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][3]$_DFFE_PN0P_  (.D(_00429_),
    .Q(\samples_real[0][3] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][4]$_DFFE_PN0P_  (.D(_00430_),
    .Q(\samples_real[0][4] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][5]$_DFFE_PN0P_  (.D(_00431_),
    .Q(\samples_real[0][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][6]$_DFFE_PN0P_  (.D(_00432_),
    .Q(\samples_real[0][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][7]$_DFFE_PN0P_  (.D(_00433_),
    .Q(\samples_real[0][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][8]$_DFFE_PN0P_  (.D(_00434_),
    .Q(\samples_real[0][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[0][9]$_DFFE_PN0P_  (.D(_00435_),
    .Q(\samples_real[0][9] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][0]$_DFFE_PN0P_  (.D(_00436_),
    .Q(\samples_real[1][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][10]$_DFFE_PN0P_  (.D(_00437_),
    .Q(\samples_real[1][10] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][11]$_DFFE_PN0P_  (.D(_00438_),
    .Q(\samples_real[1][11] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][12]$_DFFE_PN0P_  (.D(_00439_),
    .Q(\samples_real[1][12] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][13]$_DFFE_PN0P_  (.D(_00440_),
    .Q(\samples_real[1][13] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][14]$_DFFE_PN0P_  (.D(_00441_),
    .Q(\samples_real[1][14] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][15]$_DFFE_PN0P_  (.D(_00442_),
    .Q(\samples_real[1][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][1]$_DFFE_PN0P_  (.D(_00443_),
    .Q(\samples_real[1][1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[1][2]$_DFFE_PN0P_  (.D(_00444_),
    .Q(\samples_real[1][2] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[1][3]$_DFFE_PN0P_  (.D(_00445_),
    .Q(\samples_real[1][3] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[1][4]$_DFFE_PN0P_  (.D(_00446_),
    .Q(\samples_real[1][4] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[1][5]$_DFFE_PN0P_  (.D(_00447_),
    .Q(\samples_real[1][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][6]$_DFFE_PN0P_  (.D(_00448_),
    .Q(\samples_real[1][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][7]$_DFFE_PN0P_  (.D(_00449_),
    .Q(\samples_real[1][7] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[1][8]$_DFFE_PN0P_  (.D(_00450_),
    .Q(\samples_real[1][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[1][9]$_DFFE_PN0P_  (.D(_00451_),
    .Q(\samples_real[1][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][0]$_DFFE_PN0P_  (.D(_00452_),
    .Q(\samples_real[2][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][10]$_DFFE_PN0P_  (.D(_00453_),
    .Q(\samples_real[2][10] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][11]$_DFFE_PN0P_  (.D(_00454_),
    .Q(\samples_real[2][11] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][12]$_DFFE_PN0P_  (.D(_00455_),
    .Q(\samples_real[2][12] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][13]$_DFFE_PN0P_  (.D(_00456_),
    .Q(\samples_real[2][13] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][14]$_DFFE_PN0P_  (.D(_00457_),
    .Q(\samples_real[2][14] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][15]$_DFFE_PN0P_  (.D(_00458_),
    .Q(\samples_real[2][15] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][1]$_DFFE_PN0P_  (.D(_00459_),
    .Q(\samples_real[2][1] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][2]$_DFFE_PN0P_  (.D(_00460_),
    .Q(\samples_real[2][2] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[2][3]$_DFFE_PN0P_  (.D(_00461_),
    .Q(\samples_real[2][3] ),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[2][4]$_DFFE_PN0P_  (.D(_00462_),
    .Q(\samples_real[2][4] ),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[2][5]$_DFFE_PN0P_  (.D(_00463_),
    .Q(\samples_real[2][5] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][6]$_DFFE_PN0P_  (.D(_00464_),
    .Q(\samples_real[2][6] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][7]$_DFFE_PN0P_  (.D(_00465_),
    .Q(\samples_real[2][7] ),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[2][8]$_DFFE_PN0P_  (.D(_00466_),
    .Q(\samples_real[2][8] ),
    .RESET_B(net92),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[2][9]$_DFFE_PN0P_  (.D(_00467_),
    .Q(\samples_real[2][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][0]$_DFFE_PN0P_  (.D(_00468_),
    .Q(\samples_real[3][0] ),
    .RESET_B(net353),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][10]$_DFFE_PN0P_  (.D(_00469_),
    .Q(\samples_real[3][10] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[3][11]$_DFFE_PN0P_  (.D(_00470_),
    .Q(\samples_real[3][11] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[3][12]$_DFFE_PN0P_  (.D(_00471_),
    .Q(\samples_real[3][12] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][13]$_DFFE_PN0P_  (.D(_00472_),
    .Q(\samples_real[3][13] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][14]$_DFFE_PN0P_  (.D(_00473_),
    .Q(\samples_real[3][14] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[3][15]$_DFFE_PN0P_  (.D(_00474_),
    .Q(\samples_real[3][15] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][1]$_DFFE_PN0P_  (.D(_00475_),
    .Q(\samples_real[3][1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][2]$_DFFE_PN0P_  (.D(_00476_),
    .Q(\samples_real[3][2] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][3]$_DFFE_PN0P_  (.D(_00477_),
    .Q(\samples_real[3][3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \samples_real[3][4]$_DFFE_PN0P_  (.D(_00478_),
    .Q(\samples_real[3][4] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][5]$_DFFE_PN0P_  (.D(_00479_),
    .Q(\samples_real[3][5] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][6]$_DFFE_PN0P_  (.D(_00480_),
    .Q(\samples_real[3][6] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[3][7]$_DFFE_PN0P_  (.D(_00481_),
    .Q(\samples_real[3][7] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[3][8]$_DFFE_PN0P_  (.D(_00482_),
    .Q(\samples_real[3][8] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[3][9]$_DFFE_PN0P_  (.D(_00483_),
    .Q(\samples_real[3][9] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][0]$_DFFE_PN0P_  (.D(_00484_),
    .Q(\samples_real[4][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][10]$_DFFE_PN0P_  (.D(_00485_),
    .Q(\samples_real[4][10] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][11]$_DFFE_PN0P_  (.D(_00486_),
    .Q(\samples_real[4][11] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][12]$_DFFE_PN0P_  (.D(_00487_),
    .Q(\samples_real[4][12] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][13]$_DFFE_PN0P_  (.D(_00488_),
    .Q(\samples_real[4][13] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][14]$_DFFE_PN0P_  (.D(_00489_),
    .Q(\samples_real[4][14] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][15]$_DFFE_PN0P_  (.D(_00490_),
    .Q(\samples_real[4][15] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][1]$_DFFE_PN0P_  (.D(_00491_),
    .Q(\samples_real[4][1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][2]$_DFFE_PN0P_  (.D(_00492_),
    .Q(\samples_real[4][2] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][3]$_DFFE_PN0P_  (.D(_00493_),
    .Q(\samples_real[4][3] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][4]$_DFFE_PN0P_  (.D(_00494_),
    .Q(\samples_real[4][4] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][5]$_DFFE_PN0P_  (.D(_00495_),
    .Q(\samples_real[4][5] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][6]$_DFFE_PN0P_  (.D(_00496_),
    .Q(\samples_real[4][6] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][7]$_DFFE_PN0P_  (.D(_00497_),
    .Q(\samples_real[4][7] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][8]$_DFFE_PN0P_  (.D(_00498_),
    .Q(\samples_real[4][8] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[4][9]$_DFFE_PN0P_  (.D(_00499_),
    .Q(\samples_real[4][9] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][0]$_DFFE_PN0P_  (.D(_00500_),
    .Q(\samples_real[5][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][10]$_DFFE_PN0P_  (.D(_00501_),
    .Q(\samples_real[5][10] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][11]$_DFFE_PN0P_  (.D(_00502_),
    .Q(\samples_real[5][11] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][12]$_DFFE_PN0P_  (.D(_00503_),
    .Q(\samples_real[5][12] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][13]$_DFFE_PN0P_  (.D(_00504_),
    .Q(\samples_real[5][13] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][14]$_DFFE_PN0P_  (.D(_00505_),
    .Q(\samples_real[5][14] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][15]$_DFFE_PN0P_  (.D(_00506_),
    .Q(\samples_real[5][15] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][1]$_DFFE_PN0P_  (.D(_00507_),
    .Q(\samples_real[5][1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][2]$_DFFE_PN0P_  (.D(_00508_),
    .Q(\samples_real[5][2] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][3]$_DFFE_PN0P_  (.D(_00509_),
    .Q(\samples_real[5][3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][4]$_DFFE_PN0P_  (.D(_00510_),
    .Q(\samples_real[5][4] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[5][5]$_DFFE_PN0P_  (.D(_00511_),
    .Q(\samples_real[5][5] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][6]$_DFFE_PN0P_  (.D(_00512_),
    .Q(\samples_real[5][6] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][7]$_DFFE_PN0P_  (.D(_00513_),
    .Q(\samples_real[5][7] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][8]$_DFFE_PN0P_  (.D(_00514_),
    .Q(\samples_real[5][8] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[5][9]$_DFFE_PN0P_  (.D(_00515_),
    .Q(\samples_real[5][9] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][0]$_DFFE_PN0P_  (.D(_00516_),
    .Q(\samples_real[6][0] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][10]$_DFFE_PN0P_  (.D(_00517_),
    .Q(\samples_real[6][10] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][11]$_DFFE_PN0P_  (.D(_00518_),
    .Q(\samples_real[6][11] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][12]$_DFFE_PN0P_  (.D(_00519_),
    .Q(\samples_real[6][12] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][13]$_DFFE_PN0P_  (.D(_00520_),
    .Q(\samples_real[6][13] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][14]$_DFFE_PN0P_  (.D(_00521_),
    .Q(\samples_real[6][14] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][15]$_DFFE_PN0P_  (.D(_00522_),
    .Q(\samples_real[6][15] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][1]$_DFFE_PN0P_  (.D(_00523_),
    .Q(\samples_real[6][1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][2]$_DFFE_PN0P_  (.D(_00524_),
    .Q(\samples_real[6][2] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][3]$_DFFE_PN0P_  (.D(_00525_),
    .Q(\samples_real[6][3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][4]$_DFFE_PN0P_  (.D(_00526_),
    .Q(\samples_real[6][4] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][5]$_DFFE_PN0P_  (.D(_00527_),
    .Q(\samples_real[6][5] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][6]$_DFFE_PN0P_  (.D(_00528_),
    .Q(\samples_real[6][6] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][7]$_DFFE_PN0P_  (.D(_00529_),
    .Q(\samples_real[6][7] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][8]$_DFFE_PN0P_  (.D(_00530_),
    .Q(\samples_real[6][8] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[6][9]$_DFFE_PN0P_  (.D(_00531_),
    .Q(\samples_real[6][9] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][0]$_DFFE_PN0P_  (.D(_00532_),
    .Q(\samples_real[7][0] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][10]$_DFFE_PN0P_  (.D(_00533_),
    .Q(\samples_real[7][10] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][11]$_DFFE_PN0P_  (.D(_00534_),
    .Q(\samples_real[7][11] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][12]$_DFFE_PN0P_  (.D(_00535_),
    .Q(\samples_real[7][12] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[7][13]$_DFFE_PN0P_  (.D(_00536_),
    .Q(\samples_real[7][13] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_2 \samples_real[7][14]$_DFFE_PN0P_  (.D(_00537_),
    .Q(\samples_real[7][14] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][15]$_DFFE_PN0P_  (.D(_00538_),
    .Q(\samples_real[7][15] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][1]$_DFFE_PN0P_  (.D(_00539_),
    .Q(\samples_real[7][1] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][2]$_DFFE_PN0P_  (.D(_00540_),
    .Q(\samples_real[7][2] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][3]$_DFFE_PN0P_  (.D(_00541_),
    .Q(\samples_real[7][3] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][4]$_DFFE_PN0P_  (.D(_00542_),
    .Q(\samples_real[7][4] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][5]$_DFFE_PN0P_  (.D(_00543_),
    .Q(\samples_real[7][5] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][6]$_DFFE_PN0P_  (.D(_00544_),
    .Q(\samples_real[7][6] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][7]$_DFFE_PN0P_  (.D(_00545_),
    .Q(\samples_real[7][7] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][8]$_DFFE_PN0P_  (.D(_00546_),
    .Q(\samples_real[7][8] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \samples_real[7][9]$_DFFE_PN0P_  (.D(_00547_),
    .Q(\samples_real[7][9] ),
    .RESET_B(net356),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_4 \stage[0]$_DFFE_PN0P_  (.D(_00548_),
    .Q(\stage[0] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \stage[1]$_DFFE_PN0P_  (.D(_00549_),
    .Q(\stage[1] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \stage[2]$_DFFE_PN0P_  (.D(_00550_),
    .Q(\stage[2] ),
    .RESET_B(net354),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfstp_1 \state[0]$_DFF_PN1_  (.D(_00004_),
    .Q(\state[0] ),
    .SET_B(net355),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \state[1]$_DFF_PN0_  (.D(_00005_),
    .Q(\state[1] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[2]$_DFF_PN0_  (.D(_00006_),
    .Q(\state[2] ),
    .RESET_B(net355),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[3]$_DFF_PN0_  (.D(_00003_),
    .Q(\state[3] ),
    .RESET_B(net357),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \temp_imag[0]$_DFFE_PP_  (.D(_00019_),
    .DE(_00007_),
    .Q(\temp_imag[0] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \temp_real[0]$_DFFE_PP_  (.D(_00018_),
    .DE(_00007_),
    .Q(\temp_real[0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \twiddle_idx[0]$_DFFE_PP_  (.D(_05877_),
    .DE(_00007_),
    .Q(\twiddle_idx[0] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \twiddle_idx[1]$_DFFE_PP_  (.D(_05878_),
    .DE(_00007_),
    .Q(\twiddle_idx[1] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__nor3_2 clone1 (.A(_02623_),
    .B(_02559_),
    .C(_02621_),
    .Y(net1));
 sky130_fd_sc_hd__nor3_4 clone2 (.A(_02206_),
    .B(_02306_),
    .C(_02229_),
    .Y(net2));
 sky130_fd_sc_hd__a211oi_2 clone3 (.A1(_02356_),
    .A2(_02359_),
    .B1(_02374_),
    .C1(_02371_),
    .Y(net3));
 sky130_fd_sc_hd__nand3_4 clone4 (.A(_01107_),
    .B(_01105_),
    .C(_01056_),
    .Y(net4));
 sky130_fd_sc_hd__clkbuf_2 clone11 (.A(_01972_),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 clone12 (.A(_02387_),
    .X(net12));
 sky130_fd_sc_hd__nor2_2 clone13 (.A(_02389_),
    .B(_02388_),
    .Y(net13));
 sky130_fd_sc_hd__inv_6 clone14 (.A(_07667_),
    .Y(net14));
 sky130_fd_sc_hd__buf_2 clone15 (.A(_01215_),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 clone16 (.A(_02136_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 clone17 (.A(_01376_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 clone19 (.A(_02600_),
    .X(net19));
 sky130_fd_sc_hd__buf_2 clone20 (.A(_01607_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 clone21 (.A(_01201_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 clone22 (.A(_01008_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 clone23 (.A(_02390_),
    .X(net23));
 sky130_fd_sc_hd__inv_4 clone24 (.A(_07667_),
    .Y(net24));
 sky130_fd_sc_hd__clkbuf_2 clone25 (.A(_01819_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 clone26 (.A(_00652_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 clone28 (.A(_01878_),
    .X(net28));
 sky130_fd_sc_hd__buf_2 clone29 (.A(_01877_),
    .X(net29));
 sky130_fd_sc_hd__buf_6 clone30 (.A(_00819_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 clone31 (.A(_00818_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 clone32 (.A(_01006_),
    .X(net32));
 sky130_fd_sc_hd__nand2_2 clone33 (.A(_01658_),
    .B(_01730_),
    .Y(net33));
 sky130_fd_sc_hd__buf_6 clone35 (.A(_02978_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 clone37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkinv_2 clone38 (.A(net404),
    .Y(net38));
 sky130_fd_sc_hd__clkbuf_2 clone39 (.A(_01497_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 clone42 (.A(net443),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 clone44 (.A(_03299_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 clone45 (.A(_03238_),
    .X(net45));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1611 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in_imag[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in_imag[10]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in_imag[11]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(data_in_imag[12]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in_imag[13]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in_imag[14]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(data_in_imag[15]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in_imag[1]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_in_imag[2]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(data_in_imag[3]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(data_in_imag[4]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(data_in_imag[5]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in_imag[6]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(data_in_imag[7]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(data_in_imag[8]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(data_in_imag[9]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(data_in_real[0]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_in_real[10]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(data_in_real[11]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(data_in_real[12]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(data_in_real[13]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(data_in_real[14]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(data_in_real[15]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(data_in_real[1]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(data_in_real[2]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(data_in_real[3]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(data_in_real[4]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(data_in_real[5]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(data_in_real[6]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(data_in_real[7]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(data_in_real[8]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(data_in_real[9]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(net649),
    .X(net91));
 sky130_fd_sc_hd__buf_16 input34 (.A(net648),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(start),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net94),
    .X(busy));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net95),
    .X(data_out_imag[0]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net96),
    .X(data_out_imag[100]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net97),
    .X(data_out_imag[101]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net98),
    .X(data_out_imag[102]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net99),
    .X(data_out_imag[103]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net100),
    .X(data_out_imag[104]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net101),
    .X(data_out_imag[105]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net102),
    .X(data_out_imag[106]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net103),
    .X(data_out_imag[107]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net104),
    .X(data_out_imag[108]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net105),
    .X(data_out_imag[109]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net106),
    .X(data_out_imag[10]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net107),
    .X(data_out_imag[110]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net108),
    .X(data_out_imag[111]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net109),
    .X(data_out_imag[112]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net110),
    .X(data_out_imag[113]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net111),
    .X(data_out_imag[114]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net112),
    .X(data_out_imag[115]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net113),
    .X(data_out_imag[116]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net114),
    .X(data_out_imag[117]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net115),
    .X(data_out_imag[118]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net116),
    .X(data_out_imag[119]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net117),
    .X(data_out_imag[11]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net118),
    .X(data_out_imag[120]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net119),
    .X(data_out_imag[121]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net120),
    .X(data_out_imag[122]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net121),
    .X(data_out_imag[123]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net122),
    .X(data_out_imag[124]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net123),
    .X(data_out_imag[125]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net124),
    .X(data_out_imag[126]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net125),
    .X(data_out_imag[127]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net126),
    .X(data_out_imag[12]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net127),
    .X(data_out_imag[13]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net128),
    .X(data_out_imag[14]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net129),
    .X(data_out_imag[15]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net130),
    .X(data_out_imag[16]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net131),
    .X(data_out_imag[17]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net132),
    .X(data_out_imag[18]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net133),
    .X(data_out_imag[19]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net134),
    .X(data_out_imag[1]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net135),
    .X(data_out_imag[20]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net136),
    .X(data_out_imag[21]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net137),
    .X(data_out_imag[22]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net138),
    .X(data_out_imag[23]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net139),
    .X(data_out_imag[24]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net140),
    .X(data_out_imag[25]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net141),
    .X(data_out_imag[26]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net142),
    .X(data_out_imag[27]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net143),
    .X(data_out_imag[28]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net144),
    .X(data_out_imag[29]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net145),
    .X(data_out_imag[2]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net146),
    .X(data_out_imag[30]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net147),
    .X(data_out_imag[31]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net148),
    .X(data_out_imag[32]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net149),
    .X(data_out_imag[33]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net150),
    .X(data_out_imag[34]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net151),
    .X(data_out_imag[35]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net152),
    .X(data_out_imag[36]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net153),
    .X(data_out_imag[37]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net154),
    .X(data_out_imag[38]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net155),
    .X(data_out_imag[39]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net156),
    .X(data_out_imag[3]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net157),
    .X(data_out_imag[40]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net158),
    .X(data_out_imag[41]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net159),
    .X(data_out_imag[42]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net160),
    .X(data_out_imag[43]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net161),
    .X(data_out_imag[44]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net162),
    .X(data_out_imag[45]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net163),
    .X(data_out_imag[46]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net164),
    .X(data_out_imag[47]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net165),
    .X(data_out_imag[48]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net166),
    .X(data_out_imag[49]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net167),
    .X(data_out_imag[4]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net168),
    .X(data_out_imag[50]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net169),
    .X(data_out_imag[51]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net170),
    .X(data_out_imag[52]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net171),
    .X(data_out_imag[53]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net172),
    .X(data_out_imag[54]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net173),
    .X(data_out_imag[55]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net174),
    .X(data_out_imag[56]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net175),
    .X(data_out_imag[57]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net176),
    .X(data_out_imag[58]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net177),
    .X(data_out_imag[59]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net178),
    .X(data_out_imag[5]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net179),
    .X(data_out_imag[60]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net180),
    .X(data_out_imag[61]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net181),
    .X(data_out_imag[62]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net182),
    .X(data_out_imag[63]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net183),
    .X(data_out_imag[64]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net184),
    .X(data_out_imag[65]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net185),
    .X(data_out_imag[66]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net186),
    .X(data_out_imag[67]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net187),
    .X(data_out_imag[68]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net188),
    .X(data_out_imag[69]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net189),
    .X(data_out_imag[6]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net190),
    .X(data_out_imag[70]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net191),
    .X(data_out_imag[71]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net192),
    .X(data_out_imag[72]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net193),
    .X(data_out_imag[73]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net194),
    .X(data_out_imag[74]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net195),
    .X(data_out_imag[75]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net196),
    .X(data_out_imag[76]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net197),
    .X(data_out_imag[77]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net198),
    .X(data_out_imag[78]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net199),
    .X(data_out_imag[79]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net200),
    .X(data_out_imag[7]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net201),
    .X(data_out_imag[80]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net202),
    .X(data_out_imag[81]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net203),
    .X(data_out_imag[82]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net204),
    .X(data_out_imag[83]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net205),
    .X(data_out_imag[84]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net206),
    .X(data_out_imag[85]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net207),
    .X(data_out_imag[86]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net208),
    .X(data_out_imag[87]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net209),
    .X(data_out_imag[88]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net210),
    .X(data_out_imag[89]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net211),
    .X(data_out_imag[8]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net212),
    .X(data_out_imag[90]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net213),
    .X(data_out_imag[91]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net214),
    .X(data_out_imag[92]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net215),
    .X(data_out_imag[93]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net216),
    .X(data_out_imag[94]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net217),
    .X(data_out_imag[95]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net218),
    .X(data_out_imag[96]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net219),
    .X(data_out_imag[97]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net220),
    .X(data_out_imag[98]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net221),
    .X(data_out_imag[99]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net222),
    .X(data_out_imag[9]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net223),
    .X(data_out_real[0]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net224),
    .X(data_out_real[100]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net225),
    .X(data_out_real[101]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net226),
    .X(data_out_real[102]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net227),
    .X(data_out_real[103]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net228),
    .X(data_out_real[104]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net229),
    .X(data_out_real[105]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net230),
    .X(data_out_real[106]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net231),
    .X(data_out_real[107]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net232),
    .X(data_out_real[108]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net233),
    .X(data_out_real[109]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net234),
    .X(data_out_real[10]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net235),
    .X(data_out_real[110]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net236),
    .X(data_out_real[111]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net237),
    .X(data_out_real[112]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net238),
    .X(data_out_real[113]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net239),
    .X(data_out_real[114]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net240),
    .X(data_out_real[115]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net241),
    .X(data_out_real[116]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net242),
    .X(data_out_real[117]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net243),
    .X(data_out_real[118]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net244),
    .X(data_out_real[119]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net245),
    .X(data_out_real[11]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net246),
    .X(data_out_real[120]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net247),
    .X(data_out_real[121]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net248),
    .X(data_out_real[122]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net249),
    .X(data_out_real[123]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net250),
    .X(data_out_real[124]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net251),
    .X(data_out_real[125]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net252),
    .X(data_out_real[126]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net253),
    .X(data_out_real[127]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net254),
    .X(data_out_real[12]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net255),
    .X(data_out_real[13]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net256),
    .X(data_out_real[14]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net257),
    .X(data_out_real[15]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net258),
    .X(data_out_real[16]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net259),
    .X(data_out_real[17]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net260),
    .X(data_out_real[18]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net261),
    .X(data_out_real[19]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net262),
    .X(data_out_real[1]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net263),
    .X(data_out_real[20]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net264),
    .X(data_out_real[21]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net265),
    .X(data_out_real[22]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net266),
    .X(data_out_real[23]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net267),
    .X(data_out_real[24]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net268),
    .X(data_out_real[25]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net269),
    .X(data_out_real[26]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net270),
    .X(data_out_real[27]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net271),
    .X(data_out_real[28]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net272),
    .X(data_out_real[29]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net273),
    .X(data_out_real[2]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net274),
    .X(data_out_real[30]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net275),
    .X(data_out_real[31]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net276),
    .X(data_out_real[32]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net277),
    .X(data_out_real[33]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net278),
    .X(data_out_real[34]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net279),
    .X(data_out_real[35]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net280),
    .X(data_out_real[36]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net281),
    .X(data_out_real[37]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net282),
    .X(data_out_real[38]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net283),
    .X(data_out_real[39]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net284),
    .X(data_out_real[3]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net285),
    .X(data_out_real[40]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net286),
    .X(data_out_real[41]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net287),
    .X(data_out_real[42]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net288),
    .X(data_out_real[43]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net289),
    .X(data_out_real[44]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net290),
    .X(data_out_real[45]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net291),
    .X(data_out_real[46]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net292),
    .X(data_out_real[47]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net293),
    .X(data_out_real[48]));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net294),
    .X(data_out_real[49]));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net295),
    .X(data_out_real[4]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net296),
    .X(data_out_real[50]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net297),
    .X(data_out_real[51]));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net298),
    .X(data_out_real[52]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net299),
    .X(data_out_real[53]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net300),
    .X(data_out_real[54]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net301),
    .X(data_out_real[55]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net302),
    .X(data_out_real[56]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net303),
    .X(data_out_real[57]));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net304),
    .X(data_out_real[58]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net305),
    .X(data_out_real[59]));
 sky130_fd_sc_hd__clkbuf_1 output248 (.A(net306),
    .X(data_out_real[5]));
 sky130_fd_sc_hd__clkbuf_1 output249 (.A(net307),
    .X(data_out_real[60]));
 sky130_fd_sc_hd__clkbuf_1 output250 (.A(net308),
    .X(data_out_real[61]));
 sky130_fd_sc_hd__clkbuf_1 output251 (.A(net309),
    .X(data_out_real[62]));
 sky130_fd_sc_hd__clkbuf_1 output252 (.A(net310),
    .X(data_out_real[63]));
 sky130_fd_sc_hd__clkbuf_1 output253 (.A(net311),
    .X(data_out_real[64]));
 sky130_fd_sc_hd__clkbuf_1 output254 (.A(net312),
    .X(data_out_real[65]));
 sky130_fd_sc_hd__clkbuf_1 output255 (.A(net313),
    .X(data_out_real[66]));
 sky130_fd_sc_hd__clkbuf_1 output256 (.A(net314),
    .X(data_out_real[67]));
 sky130_fd_sc_hd__clkbuf_1 output257 (.A(net315),
    .X(data_out_real[68]));
 sky130_fd_sc_hd__clkbuf_1 output258 (.A(net316),
    .X(data_out_real[69]));
 sky130_fd_sc_hd__clkbuf_1 output259 (.A(net317),
    .X(data_out_real[6]));
 sky130_fd_sc_hd__clkbuf_1 output260 (.A(net318),
    .X(data_out_real[70]));
 sky130_fd_sc_hd__clkbuf_1 output261 (.A(net319),
    .X(data_out_real[71]));
 sky130_fd_sc_hd__clkbuf_1 output262 (.A(net320),
    .X(data_out_real[72]));
 sky130_fd_sc_hd__clkbuf_1 output263 (.A(net321),
    .X(data_out_real[73]));
 sky130_fd_sc_hd__clkbuf_1 output264 (.A(net322),
    .X(data_out_real[74]));
 sky130_fd_sc_hd__clkbuf_1 output265 (.A(net323),
    .X(data_out_real[75]));
 sky130_fd_sc_hd__clkbuf_1 output266 (.A(net324),
    .X(data_out_real[76]));
 sky130_fd_sc_hd__clkbuf_1 output267 (.A(net325),
    .X(data_out_real[77]));
 sky130_fd_sc_hd__clkbuf_1 output268 (.A(net326),
    .X(data_out_real[78]));
 sky130_fd_sc_hd__clkbuf_1 output269 (.A(net327),
    .X(data_out_real[79]));
 sky130_fd_sc_hd__clkbuf_1 output270 (.A(net328),
    .X(data_out_real[7]));
 sky130_fd_sc_hd__clkbuf_1 output271 (.A(net329),
    .X(data_out_real[80]));
 sky130_fd_sc_hd__clkbuf_1 output272 (.A(net330),
    .X(data_out_real[81]));
 sky130_fd_sc_hd__clkbuf_1 output273 (.A(net331),
    .X(data_out_real[82]));
 sky130_fd_sc_hd__clkbuf_1 output274 (.A(net332),
    .X(data_out_real[83]));
 sky130_fd_sc_hd__clkbuf_1 output275 (.A(net333),
    .X(data_out_real[84]));
 sky130_fd_sc_hd__clkbuf_1 output276 (.A(net334),
    .X(data_out_real[85]));
 sky130_fd_sc_hd__clkbuf_1 output277 (.A(net335),
    .X(data_out_real[86]));
 sky130_fd_sc_hd__clkbuf_1 output278 (.A(net336),
    .X(data_out_real[87]));
 sky130_fd_sc_hd__clkbuf_1 output279 (.A(net337),
    .X(data_out_real[88]));
 sky130_fd_sc_hd__clkbuf_1 output280 (.A(net338),
    .X(data_out_real[89]));
 sky130_fd_sc_hd__clkbuf_1 output281 (.A(net339),
    .X(data_out_real[8]));
 sky130_fd_sc_hd__clkbuf_1 output282 (.A(net340),
    .X(data_out_real[90]));
 sky130_fd_sc_hd__clkbuf_1 output283 (.A(net341),
    .X(data_out_real[91]));
 sky130_fd_sc_hd__clkbuf_1 output284 (.A(net342),
    .X(data_out_real[92]));
 sky130_fd_sc_hd__clkbuf_1 output285 (.A(net343),
    .X(data_out_real[93]));
 sky130_fd_sc_hd__clkbuf_1 output286 (.A(net344),
    .X(data_out_real[94]));
 sky130_fd_sc_hd__clkbuf_1 output287 (.A(net345),
    .X(data_out_real[95]));
 sky130_fd_sc_hd__clkbuf_1 output288 (.A(net346),
    .X(data_out_real[96]));
 sky130_fd_sc_hd__clkbuf_1 output289 (.A(net347),
    .X(data_out_real[97]));
 sky130_fd_sc_hd__clkbuf_1 output290 (.A(net348),
    .X(data_out_real[98]));
 sky130_fd_sc_hd__clkbuf_1 output291 (.A(net349),
    .X(data_out_real[99]));
 sky130_fd_sc_hd__clkbuf_1 output292 (.A(net350),
    .X(data_out_real[9]));
 sky130_fd_sc_hd__clkbuf_1 output293 (.A(net351),
    .X(data_ready));
 sky130_fd_sc_hd__clkbuf_1 output294 (.A(net352),
    .X(data_valid_out));
 sky130_fd_sc_hd__buf_16 load_slew295 (.A(net92),
    .X(net353));
 sky130_fd_sc_hd__buf_16 load_slew296 (.A(net92),
    .X(net354));
 sky130_fd_sc_hd__buf_16 load_slew297 (.A(net357),
    .X(net355));
 sky130_fd_sc_hd__buf_16 load_slew298 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__buf_16 load_slew299 (.A(net92),
    .X(net357));
 sky130_fd_sc_hd__conb_1 _15301__300 (.LO(net358));
 sky130_fd_sc_hd__conb_1 _15305__301 (.LO(net359));
 sky130_fd_sc_hd__conb_1 _15310__302 (.LO(net360));
 sky130_fd_sc_hd__conb_1 _15312__303 (.LO(net361));
 sky130_fd_sc_hd__conb_1 _15323__304 (.LO(net362));
 sky130_fd_sc_hd__conb_1 _15330__305 (.LO(net363));
 sky130_fd_sc_hd__conb_1 _15338__306 (.LO(net364));
 sky130_fd_sc_hd__conb_1 _15345__307 (.LO(net365));
 sky130_fd_sc_hd__conb_1 _15351__308 (.LO(net366));
 sky130_fd_sc_hd__conb_1 _15359__309 (.LO(net367));
 sky130_fd_sc_hd__conb_1 _15364__310 (.LO(net368));
 sky130_fd_sc_hd__conb_1 _15373__311 (.LO(net369));
 sky130_fd_sc_hd__conb_1 _15380__312 (.LO(net370));
 sky130_fd_sc_hd__conb_1 _15387__313 (.LO(net371));
 sky130_fd_sc_hd__conb_1 _15388__314 (.LO(net372));
 sky130_fd_sc_hd__conb_1 _15396__315 (.LO(net373));
 sky130_fd_sc_hd__conb_1 _15404__316 (.LO(net374));
 sky130_fd_sc_hd__conb_1 _15412__317 (.LO(net375));
 sky130_fd_sc_hd__conb_1 _15420__318 (.LO(net376));
 sky130_fd_sc_hd__conb_1 _15428__319 (.LO(net377));
 sky130_fd_sc_hd__conb_1 _15436__320 (.LO(net378));
 sky130_fd_sc_hd__conb_1 _15443__321 (.LO(net379));
 sky130_fd_sc_hd__conb_1 _15444__322 (.LO(net380));
 sky130_fd_sc_hd__conb_1 _15452__323 (.LO(net381));
 sky130_fd_sc_hd__conb_1 _15459__324 (.LO(net382));
 sky130_fd_sc_hd__conb_1 _15470__325 (.LO(net383));
 sky130_fd_sc_hd__conb_1 _15475__326 (.LO(net384));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_1 clkload2 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_1 clkload7 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload9 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload11 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__bufinv_16 clkload14 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_4 clkload15 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload16 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload17 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload18 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload19 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload20 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload21 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload22 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__bufinv_16 clkload26 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload27 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__bufinv_16 clkload28 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload29 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_2 clkload30 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload32 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_2 clkload33 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_2 clkload34 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_2 clkload35 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload36 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload37 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__bufinv_16 clkload38 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload39 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__bufinv_16 clkload41 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__bufinv_16 clkload44 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload45 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload47 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload48 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__inv_6 clkload50 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload51 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__inv_6 clkload52 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__inv_8 clkload53 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_07667_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(_07667_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net411),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_02780_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_02701_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer6 (.A(_02963_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net407),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(_02784_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net393),
    .X(net394));
 sky130_fd_sc_hd__buf_2 rebuffer10 (.A(_02978_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(_02700_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(_07677_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(net418),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net398),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(_02778_),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_16 clone34 (.A(_01390_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(_02785_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer36 (.A(_02861_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(_02861_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net404),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net405),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(_02962_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer42 (.A(_02960_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(_02958_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer50 (.A(net414),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer51 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer53 (.A(net421),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_2 rebuffer54 (.A(_07677_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer55 (.A(net433),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(_02862_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer57 (.A(net423),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer58 (.A(_02862_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer59 (.A(_02862_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(_07675_),
    .X(net427));
 sky130_fd_sc_hd__buf_4 rebuffer61 (.A(_01960_),
    .X(net428));
 sky130_fd_sc_hd__buf_2 rebuffer75 (.A(_03463_),
    .X(net442));
 sky130_fd_sc_hd__buf_6 rebuffer76 (.A(\idx2[2] ),
    .X(net443));
 sky130_fd_sc_hd__buf_2 rebuffer77 (.A(net443),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net443),
    .X(net445));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer79 (.A(net445),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net443),
    .X(net447));
 sky130_fd_sc_hd__buf_2 rebuffer81 (.A(_06041_),
    .X(net448));
 sky130_fd_sc_hd__buf_2 rebuffer82 (.A(_06041_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(_06041_),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_16 clone84 (.A(_03237_),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_16 clone85 (.A(net470),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer86 (.A(_05962_),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 rebuffer87 (.A(_05962_),
    .X(net454));
 sky130_fd_sc_hd__buf_6 rebuffer88 (.A(_03442_),
    .X(net455));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer89 (.A(net455),
    .X(net456));
 sky130_fd_sc_hd__buf_12 rebuffer93 (.A(_03342_),
    .X(net462));
 sky130_fd_sc_hd__buf_6 rebuffer104 (.A(_08146_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer105 (.A(net471),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer106 (.A(net471),
    .X(net473));
 sky130_fd_sc_hd__buf_1 rebuffer107 (.A(\idx2[0] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer108 (.A(net474),
    .X(net475));
 sky130_fd_sc_hd__buf_2 rebuffer109 (.A(_03269_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer110 (.A(net476),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer111 (.A(_03324_),
    .X(net478));
 sky130_fd_sc_hd__buf_6 rebuffer112 (.A(_03354_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer113 (.A(net479),
    .X(net480));
 sky130_fd_sc_hd__buf_4 rebuffer114 (.A(net480),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer115 (.A(_03277_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer116 (.A(_03378_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer117 (.A(net483),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer118 (.A(_03378_),
    .X(net485));
 sky130_fd_sc_hd__buf_6 rebuffer119 (.A(_06729_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer120 (.A(net486),
    .X(net487));
 sky130_fd_sc_hd__buf_6 rebuffer121 (.A(net486),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer122 (.A(net488),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer123 (.A(net488),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer124 (.A(net490),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer125 (.A(net486),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_2 rebuffer126 (.A(\idx2[1] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer127 (.A(net493),
    .X(net494));
 sky130_fd_sc_hd__buf_6 rebuffer128 (.A(_03308_),
    .X(net495));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer129 (.A(net495),
    .X(net496));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer130 (.A(net495),
    .X(net497));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer131 (.A(_03415_),
    .X(net498));
 sky130_fd_sc_hd__buf_2 rebuffer132 (.A(net440),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer133 (.A(net499),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer134 (.A(net499),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer135 (.A(_03393_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer136 (.A(net502),
    .X(net503));
 sky130_fd_sc_hd__buf_6 rebuffer137 (.A(_03386_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer138 (.A(net504),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer139 (.A(_03277_),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_2 rebuffer140 (.A(\idx2[0] ),
    .X(net507));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer141 (.A(_03325_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer142 (.A(_03242_),
    .X(net509));
 sky130_fd_sc_hd__buf_6 rebuffer147 (.A(\idx1[1] ),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_2 rebuffer148 (.A(net514),
    .X(net515));
 sky130_fd_sc_hd__buf_6 rebuffer149 (.A(net579),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer150 (.A(net635),
    .X(net517));
 sky130_fd_sc_hd__buf_12 rebuffer151 (.A(_03923_),
    .X(net518));
 sky130_fd_sc_hd__buf_6 rebuffer152 (.A(\idx1[2] ),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_2 rebuffer153 (.A(net519),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer154 (.A(net519),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer155 (.A(net521),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer156 (.A(net531),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer157 (.A(_03922_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer158 (.A(_03922_),
    .X(net525));
 sky130_fd_sc_hd__buf_6 rebuffer159 (.A(\idx1[0] ),
    .X(net526));
 sky130_fd_sc_hd__buf_2 rebuffer231 (.A(net601),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer161 (.A(net572),
    .X(net528));
 sky130_fd_sc_hd__buf_2 rebuffer162 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_1 rebuffer163 (.A(net532),
    .X(net530));
 sky130_fd_sc_hd__buf_1 rebuffer165 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__buf_1 rebuffer166 (.A(net537),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer168 (.A(_03156_),
    .X(net535));
 sky130_fd_sc_hd__buf_4 rebuffer169 (.A(_03156_),
    .X(net536));
 sky130_fd_sc_hd__buf_1 rebuffer170 (.A(net558),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer171 (.A(_03155_),
    .X(net538));
 sky130_fd_sc_hd__buf_2 clone172 (.A(net540),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer173 (.A(_03154_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer174 (.A(_03913_),
    .X(net541));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer175 (.A(_03990_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer176 (.A(_03917_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer177 (.A(_03909_),
    .X(net544));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer178 (.A(_03947_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer179 (.A(net633),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer180 (.A(_03196_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer181 (.A(net547),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer182 (.A(net596),
    .X(net549));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer183 (.A(net549),
    .X(net550));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer184 (.A(net549),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer185 (.A(_03161_),
    .X(net552));
 sky130_fd_sc_hd__buf_6 rebuffer186 (.A(net595),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer187 (.A(_03951_),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_2 rebuffer188 (.A(_03160_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer189 (.A(net598),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer190 (.A(_03955_),
    .X(net557));
 sky130_fd_sc_hd__buf_1 rebuffer191 (.A(net602),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer192 (.A(_03152_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer193 (.A(_03152_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer194 (.A(_03152_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer195 (.A(net561),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer196 (.A(_03963_),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 rebuffer198 (.A(_05039_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer199 (.A(net565),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 rebuffer200 (.A(net611),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_16 clone201 (.A(_05040_),
    .X(net568));
 sky130_fd_sc_hd__buf_2 rebuffer202 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_1 rebuffer203 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_1 rebuffer204 (.A(net585),
    .X(net571));
 sky130_fd_sc_hd__buf_6 rebuffer205 (.A(net526),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer206 (.A(_05032_),
    .X(net573));
 sky130_fd_sc_hd__buf_4 rebuffer207 (.A(_03167_),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 rebuffer208 (.A(_03153_),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 rebuffer209 (.A(_03153_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer210 (.A(_05092_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer211 (.A(_05885_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_2 rebuffer212 (.A(net514),
    .X(net579));
 sky130_fd_sc_hd__buf_4 rebuffer213 (.A(_03167_),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 rebuffer214 (.A(_05082_),
    .X(net581));
 sky130_fd_sc_hd__buf_8 rebuffer215 (.A(_03167_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer216 (.A(net582),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer217 (.A(_03175_),
    .X(net584));
 sky130_fd_sc_hd__buf_1 rebuffer218 (.A(net512),
    .X(net585));
 sky130_fd_sc_hd__buf_4 rebuffer219 (.A(_03164_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer220 (.A(net586),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer221 (.A(_05887_),
    .X(net588));
 sky130_fd_sc_hd__buf_2 rebuffer222 (.A(_03149_),
    .X(net589));
 sky130_fd_sc_hd__buf_8 rebuffer223 (.A(_03149_),
    .X(net590));
 sky130_fd_sc_hd__buf_4 rebuffer224 (.A(_03153_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer225 (.A(_05070_),
    .X(net592));
 sky130_fd_sc_hd__buf_1 rebuffer235 (.A(net637),
    .X(net602));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer229 (.A(_03170_),
    .X(net600));
 sky130_fd_sc_hd__buf_6 rebuffer243 (.A(_07732_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer246 (.A(_03202_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer247 (.A(net613),
    .X(net614));
 sky130_fd_sc_hd__buf_6 rebuffer248 (.A(_03161_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer249 (.A(_03967_),
    .X(net616));
 sky130_fd_sc_hd__buf_2 rebuffer266 (.A(net65),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer267 (.A(net516),
    .X(net634));
 sky130_fd_sc_hd__buf_2 rebuffer268 (.A(net634),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer269 (.A(net635),
    .X(net636));
 sky130_fd_sc_hd__buf_8 rebuffer270 (.A(_07846_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer271 (.A(_03934_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer272 (.A(_04016_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer273 (.A(_03209_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer274 (.A(_03959_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer275 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_16 clone276 (.A(net591),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer277 (.A(_03930_),
    .X(net644));
 sky130_fd_sc_hd__buf_8 rebuffer279 (.A(_04045_),
    .X(net646));
 sky130_fd_sc_hd__buf_6 rebuffer280 (.A(_04097_),
    .X(net647));
 sky130_fd_sc_hd__buf_16 load_slew1 (.A(\temp_real[0] ),
    .X(net53));
 sky130_fd_sc_hd__nor2_4 clone40 (.A(_01870_),
    .B(_01886_),
    .Y(net410));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer43 (.A(_02692_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(_07674_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer64 (.A(net431),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer65 (.A(_02957_),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_16 clone67 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_2 rebuffer68 (.A(_02863_),
    .X(net435));
 sky130_fd_sc_hd__buf_8 rebuffer71 (.A(_03362_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(net438),
    .X(net439));
 sky130_fd_sc_hd__buf_6 rebuffer73 (.A(_03415_),
    .X(net440));
 sky130_fd_sc_hd__buf_6 rebuffer74 (.A(_03269_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer84 (.A(net441),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer85 (.A(_06713_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(_06713_),
    .X(net460));
 sky130_fd_sc_hd__buf_6 rebuffer92 (.A(_03607_),
    .X(net461));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer94 (.A(net462),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer95 (.A(net463),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 rebuffer96 (.A(_03319_),
    .X(net465));
 sky130_fd_sc_hd__buf_6 rebuffer97 (.A(_06631_),
    .X(net466));
 sky130_fd_sc_hd__buf_6 rebuffer98 (.A(_03463_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer99 (.A(_03463_),
    .X(net468));
 sky130_fd_sc_hd__buf_4 rebuffer100 (.A(_03238_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer101 (.A(_03235_),
    .X(net470));
 sky130_fd_sc_hd__buf_6 rebuffer102 (.A(_03286_),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_2 rebuffer143 (.A(_07732_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer144 (.A(_05045_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer145 (.A(_05057_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer146 (.A(_05039_),
    .X(net593));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer172 (.A(_05887_),
    .X(net594));
 sky130_fd_sc_hd__buf_6 rebuffer197 (.A(_03161_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer201 (.A(_03161_),
    .X(net596));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer226 (.A(_05074_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer227 (.A(_03160_),
    .X(net598));
 sky130_fd_sc_hd__buf_2 rebuffer228 (.A(_05078_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer232 (.A(_03165_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer233 (.A(_03165_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer234 (.A(net605),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer236 (.A(_03164_),
    .X(net607));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer239 (.A(_05105_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer240 (.A(_07792_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer241 (.A(_07792_),
    .X(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_04194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\samples_imag[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\samples_imag[1][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\samples_imag[2][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\samples_imag[2][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\samples_imag[3][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\samples_imag[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\samples_imag[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\samples_real[0][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\samples_real[0][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\samples_real[0][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\samples_real[0][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\samples_real[0][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\samples_real[0][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\samples_real[1][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\samples_real[2][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\samples_real[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\samples_real[7][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\samples_real[7][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\samples_imag[0][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\samples_real[0][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\samples_real[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\samples_real[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\samples_real[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net163));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_752 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_654 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_632 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_752 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
endmodule
