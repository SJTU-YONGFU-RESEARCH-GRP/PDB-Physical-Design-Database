module parameterized_self_correcting_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net7;

 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _15_ (.A1(net4),
    .A2(net5),
    .B(net6),
    .ZN(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _16_ (.A1(net2),
    .A2(_04_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _17_ (.I(net2),
    .ZN(_06_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _18_ (.I0(_05_),
    .I1(_06_),
    .S(net3),
    .Z(_00_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _19_ (.I(net6),
    .ZN(_07_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _20_ (.A1(net3),
    .A2(_07_),
    .A3(net2),
    .Z(_08_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _21_ (.A1(net3),
    .A2(net6),
    .B(net2),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _22_ (.I0(_08_),
    .I1(_09_),
    .S(net4),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _23_ (.A1(net3),
    .A2(net4),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _24_ (.A1(_07_),
    .A2(net2),
    .A3(_10_),
    .Z(_11_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _25_ (.A1(net6),
    .A2(_10_),
    .B(net2),
    .ZN(_12_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _26_ (.I0(_11_),
    .I1(_12_),
    .S(net5),
    .Z(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _27_ (.A1(net5),
    .A2(net2),
    .A3(_10_),
    .Z(_13_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _28_ (.A1(net3),
    .A2(net4),
    .A3(net5),
    .B(net2),
    .ZN(_14_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _29_ (.I0(_13_),
    .I1(_14_),
    .S(net6),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \counter_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 hold1 (.I(net7),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_46 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_47 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_48 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_50 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_55 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input1 (.I(enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output2 (.I(net3),
    .Z(count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net4),
    .Z(count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output4 (.I(net5),
    .Z(count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output5 (.I(net6),
    .Z(count[3]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_196 ();
endmodule
