
* cell configurable_lfsr
* pin parallel_out[2]
* pin seed[1]
* pin parallel_out[1]
* pin seed[0]
* pin parallel_out[0]
* pin rst_n
* pin serial_out
* pin seed[2]
* pin tap_pattern[0]
* pin tap_pattern[1]
* pin enable
* pin tap_pattern[2]
* pin seed[3]
* pin parallel_out[3]
* pin tap_pattern[3]
* pin tap_pattern[7]
* pin load_seed
* pin parallel_out[4]
* pin parallel_out[7]
* pin seed[4]
* pin seed[7]
* pin seed[5]
* pin clk
* pin tap_pattern[4]
* pin parallel_out[5]
* pin tap_pattern[6]
* pin seed[6]
* pin parallel_out[6]
* pin tap_pattern[5]
.SUBCKT configurable_lfsr 1 2 3 4 17 18 20 28 29 30 35 39 41 42 52 55 65 66 69
+ 75 78 82 83 98 99 100 102 103 104
* net 1 parallel_out[2]
* net 2 seed[1]
* net 3 parallel_out[1]
* net 4 seed[0]
* net 17 parallel_out[0]
* net 18 rst_n
* net 20 serial_out
* net 28 seed[2]
* net 29 tap_pattern[0]
* net 30 tap_pattern[1]
* net 35 enable
* net 39 tap_pattern[2]
* net 41 seed[3]
* net 42 parallel_out[3]
* net 52 tap_pattern[3]
* net 55 tap_pattern[7]
* net 65 load_seed
* net 66 parallel_out[4]
* net 69 parallel_out[7]
* net 75 seed[4]
* net 78 seed[7]
* net 82 seed[5]
* net 83 clk
* net 98 tap_pattern[4]
* net 99 parallel_out[5]
* net 100 tap_pattern[6]
* net 102 seed[6]
* net 103 parallel_out[6]
* net 104 tap_pattern[5]
* cell instance $3 r0 *1 23.46,2.72
X$3 7 5 1 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $5 r0 *1 27.6,2.72
X$5 7 2 8 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $8 m0 *1 32.2,8.16
X$8 7 15 3 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $12 r0 *1 31.28,2.72
X$12 7 4 9 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $19 r0 *1 10.12,19.04
X$19 6 21 5 37 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $22 m0 *1 6.44,24.48
X$22 6 23 5 45 32 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $25 r0 *1 26.68,19.04
X$25 6 27 15 5 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $27 r0 *1 47.84,24.48
X$27 7 5 38 51 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $135 r0 *1 27.6,13.6
X$135 7 10 8 12 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $137 r0 *1 30.82,13.6
X$137 7 10 9 11 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $153 m0 *1 4.14,19.04
X$153 7 28 13 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $155 m0 *1 5.98,19.04
X$155 7 10 13 31 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $163 m0 *1 27.14,19.04
X$163 7 10 27 12 7 14 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $165 m0 *1 29.44,19.04
X$165 6 23 15 19 14 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $170 m0 *1 53.36,19.04
X$170 7 16 17 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $171 m0 *1 54.74,19.04
X$171 7 25 16 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $172 r0 *1 1.38,19.04
X$172 7 18 7 24 6 6 sky130_fd_sc_hd__dlygate4sd3_1
* cell instance $173 r0 *1 5.06,19.04
X$173 7 24 6 23 7 6 sky130_fd_sc_hd__clkbuf_4
* cell instance $174 r0 *1 7.82,19.04
X$174 7 10 21 31 7 32 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $183 r0 *1 30.36,19.04
X$183 7 10 36 11 7 26 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $184 r0 *1 32.2,19.04
X$184 6 23 25 19 26 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $193 r0 *1 53.36,19.04
X$193 7 29 33 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $194 r0 *1 54.74,19.04
X$194 7 25 20 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $211 m0 *1 34.5,24.48
X$211 6 36 25 15 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $213 m0 *1 39.1,24.48
X$213 7 15 34 40 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $216 m0 *1 42.78,24.48
X$216 7 30 34 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $219 m0 *1 49.68,24.48
X$219 7 33 25 44 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $220 m0 *1 51.06,24.48
X$220 7 35 6 22 7 6 sky130_fd_sc_hd__clkbuf_4
* cell instance $224 r0 *1 1.84,24.48
X$224 7 37 42 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $225 r0 *1 3.22,24.48
X$225 6 23 37 45 64 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $236 r0 *1 31.74,24.48
X$236 7 47 6 19 7 6 sky130_fd_sc_hd__clkbuf_4
* cell instance $238 r0 *1 36.34,24.48
X$238 7 44 40 7 46 6 6 sky130_fd_sc_hd__xor2_1
* cell instance $247 r0 *1 51.06,24.48
X$247 7 39 38 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $249 m0 *1 1.38,29.92
X$249 7 41 53 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $250 m0 *1 2.76,29.92
X$250 7 52 56 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $252 m0 *1 4.6,29.92
X$252 7 10 53 70 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $253 m0 *1 5.98,29.92
X$253 7 47 6 45 7 6 sky130_fd_sc_hd__clkbuf_4
* cell instance $254 m0 *1 8.74,29.92
X$254 6 23 43 45 58 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $257 m0 *1 17.94,29.92
X$257 7 83 6 47 7 6 sky130_fd_sc_hd__clkbuf_4
* cell instance $265 m0 *1 37.72,29.92
X$265 7 48 59 57 7 6 6 sky130_fd_sc_hd__xnor2_1
* cell instance $266 m0 *1 40.94,29.92
X$266 7 49 46 48 7 6 6 sky130_fd_sc_hd__xnor2_1
* cell instance $271 m0 *1 46.92,29.92
X$271 7 51 54 49 7 6 6 sky130_fd_sc_hd__xnor2_1
* cell instance $273 m0 *1 50.6,29.92
X$273 7 63 50 54 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $275 m0 *1 52.9,29.92
X$275 7 55 50 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $278 r0 *1 1.84,29.92
X$278 7 43 66 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $280 r0 *1 4.14,29.92
X$280 7 67 60 70 7 64 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $281 r0 *1 5.98,29.92
X$281 7 37 56 61 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $283 r0 *1 7.82,29.92
X$283 7 67 68 79 7 58 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $284 r0 *1 9.66,29.92
X$284 6 60 37 43 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $288 r0 *1 15.64,29.92
X$288 6 68 43 73 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $291 r0 *1 22.08,29.92
X$291 7 61 90 7 74 6 6 sky130_fd_sc_hd__xor2_1
* cell instance $294 r0 *1 29.9,29.92
X$294 6 23 63 19 62 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $295 r0 *1 39.1,29.92
X$295 7 57 80 72 7 62 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $297 r0 *1 41.4,29.92
X$297 7 67 22 71 6 7 6 sky130_fd_sc_hd__nor2_1
* cell instance $303 r0 *1 51.52,29.92
X$303 7 63 69 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $311 m0 *1 1.38,35.36
X$311 7 65 7 6 67 6 sky130_fd_sc_hd__clkbuf_2
* cell instance $312 m0 *1 3.22,35.36
X$312 7 75 76 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $315 m0 *1 5.98,35.36
X$315 7 10 76 79 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $318 m0 *1 10.12,35.36
X$318 6 23 73 45 86 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $321 m0 *1 23.46,35.36
X$321 7 67 6 10 7 6 sky130_fd_sc_hd__buf_2
* cell instance $322 m0 *1 25.3,35.36
X$322 7 93 74 59 7 6 6 sky130_fd_sc_hd__xnor2_1
* cell instance $326 m0 *1 29.9,35.36
X$326 6 23 81 19 87 7 7 6 sky130_fd_sc_hd__dfrtp_1
* cell instance $328 m0 *1 39.56,35.36
X$328 7 22 67 80 6 7 6 sky130_fd_sc_hd__nand2b_1
* cell instance $329 m0 *1 41.86,35.36
X$329 7 63 71 67 77 7 72 6 6 sky130_fd_sc_hd__a22oi_1
* cell instance $331 m0 *1 46.46,35.36
X$331 7 78 77 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $337 r0 *1 5.52,35.36
X$337 7 82 88 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $340 r0 *1 8.28,35.36
X$340 7 10 88 89 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $341 r0 *1 9.66,35.36
X$341 7 67 84 89 7 86 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $348 r0 *1 20.7,35.36
X$348 6 84 73 81 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $349 r0 *1 24.38,35.36
X$349 7 43 97 92 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $352 r0 *1 30.36,35.36
X$352 7 10 101 91 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $353 r0 *1 31.74,35.36
X$353 7 67 85 91 7 87 6 6 sky130_fd_sc_hd__o21ai_0
* cell instance $356 r0 *1 37.72,35.36
X$356 6 85 81 63 22 7 7 6 sky130_fd_sc_hd__mux2i_1
* cell instance $374 m0 *1 22.54,40.8
X$374 7 73 96 90 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $375 m0 *1 23.92,40.8
X$375 7 92 95 93 7 6 6 sky130_fd_sc_hd__xnor2_1
* cell instance $450 m0 *1 23,51.68
X$450 7 104 96 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $453 m0 *1 24.38,51.68
X$453 7 98 97 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $454 r0 *1 24.38,46.24
X$454 7 81 94 95 7 6 6 sky130_fd_sc_hd__nand2_1
* cell instance $493 r0 *1 22.54,51.68
X$493 7 73 99 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $496 r0 *1 25.3,51.68
X$496 7 100 94 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $502 r0 *1 30.82,51.68
X$502 7 102 101 6 7 6 sky130_fd_sc_hd__clkbuf_1
* cell instance $506 r0 *1 38.64,51.68
X$506 7 81 103 6 7 6 sky130_fd_sc_hd__clkbuf_1
.ENDS configurable_lfsr

* cell sky130_fd_sc_hd__dlygate4sd3_1
* pin VPB
* pin A
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__dlygate4sd3_1 1 3 5 7 8 9
* net 1 VPB
* net 3 A
* net 5 VPWR
* net 7 X
* net 8 VGND
* device instance $1 r0 *1 2.465,2.275 pfet_01v8_hvt
M$1 6 2 5 1 pfet_01v8_hvt L=500000U W=420000U AS=140750000000P AD=109200000000P
+ PS=1325000U PD=1360000U
* device instance $2 r0 *1 3.115,1.985 pfet_01v8_hvt
M$2 7 6 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $3 r0 *1 0.58,2.275 pfet_01v8_hvt
M$3 5 3 4 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $4 r0 *1 1.175,2.275 pfet_01v8_hvt
M$4 2 4 5 1 pfet_01v8_hvt L=500000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $5 r0 *1 2.465,0.445 nfet_01v8
M$5 8 2 6 9 nfet_01v8 L=500000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $6 r0 *1 3.115,0.56 nfet_01v8
M$6 7 6 8 9 nfet_01v8 L=150000U W=650000U AS=97000000000P AD=169000000000P
+ PS=975000U PD=1820000U
* device instance $7 r0 *1 0.58,0.445 nfet_01v8
M$7 8 3 4 9 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $8 r0 *1 1.175,0.445 nfet_01v8
M$8 2 4 8 9 nfet_01v8 L=500000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__dlygate4sd3_1

* cell sky130_fd_sc_hd__buf_2
* pin VPB
* pin A
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__buf_2 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 VGND
* net 5 X
* net 6 VPWR
* device instance $1 r0 *1 0.47,2.125 pfet_01v8_hvt
M$1 2 3 6 1 pfet_01v8_hvt L=150000U W=640000U AS=149000000000P AD=166400000000P
+ PS=1325000U PD=1800000U
* device instance $2 r0 *1 0.945,1.985 pfet_01v8_hvt
M$2 5 2 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=284000000000P
+ AD=400000000000P PS=2595000U PD=3800000U
* device instance $4 r0 *1 0.47,0.445 nfet_01v8
M$4 4 3 2 7 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $5 r0 *1 0.945,0.56 nfet_01v8
M$5 5 2 4 7 nfet_01v8 L=150000U W=1300000U AS=184750000000P AD=260000000000P
+ PS=1895000U PD=2750000U
.ENDS sky130_fd_sc_hd__buf_2

* cell sky130_fd_sc_hd__xor2_1
* pin VPB
* pin B
* pin A
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__xor2_1 1 2 3 6 7 8 9
* net 1 VPB
* net 2 B
* net 3 A
* net 6 VPWR
* net 7 X
* net 8 VGND
* device instance $1 r0 *1 2.71,1.985 pfet_01v8_hvt
M$1 7 4 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=300000000000P PS=2520000U PD=2600000U
* device instance $2 r0 *1 0.51,1.985 pfet_01v8_hvt
M$2 10 2 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $3 r0 *1 0.93,1.985 pfet_01v8_hvt
M$3 6 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $4 r0 *1 1.35,1.985 pfet_01v8_hvt
M$4 5 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $5 r0 *1 1.77,1.985 pfet_01v8_hvt
M$5 6 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $6 r0 *1 0.51,0.56 nfet_01v8
M$6 4 2 8 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 0.93,0.56 nfet_01v8
M$7 8 3 4 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $8 r0 *1 1.35,0.56 nfet_01v8
M$8 11 3 8 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $9 r0 *1 1.77,0.56 nfet_01v8
M$9 7 2 11 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=250250000000P
+ PS=920000U PD=1420000U
* device instance $10 r0 *1 2.69,0.56 nfet_01v8
M$10 8 4 7 9 nfet_01v8 L=150000U W=650000U AS=250250000000P AD=208000000000P
+ PS=1420000U PD=1940000U
.ENDS sky130_fd_sc_hd__xor2_1

* cell sky130_fd_sc_hd__clkbuf_2
* pin VPB
* pin A
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_2 1 2 3 4 6 7
* net 1 VPB
* net 2 A
* net 3 VPWR
* net 4 VGND
* net 6 X
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 3 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=162500000000P PS=2530000U PD=1325000U
* device instance $2 r0 *1 0.95,1.985 pfet_01v8_hvt
M$2 6 5 3 1 pfet_01v8_hvt L=150000U W=2000000U AS=297500000000P
+ AD=395000000000P PS=2595000U PD=3790000U
* device instance $4 r0 *1 0.475,0.445 nfet_01v8
M$4 4 2 5 7 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=68250000000P
+ PS=1370000U PD=745000U
* device instance $5 r0 *1 0.95,0.445 nfet_01v8
M$5 6 5 4 7 nfet_01v8 L=150000U W=840000U AS=124950000000P AD=165900000000P
+ PS=1435000U PD=2050000U
.ENDS sky130_fd_sc_hd__clkbuf_2

* cell sky130_fd_sc_hd__a22oi_1
* pin VPB
* pin B2
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a22oi_1 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 7 VPWR
* net 8 Y
* net 9 VGND
* device instance $1 r0 *1 1.83,1.985 pfet_01v8_hvt
M$1 6 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.25,1.985 pfet_01v8_hvt
M$2 7 5 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=300000000000P PS=1270000U PD=2600000U
* device instance $3 r0 *1 0.47,1.985 pfet_01v8_hvt
M$3 6 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $4 r0 *1 0.89,1.985 pfet_01v8_hvt
M$4 8 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $5 r0 *1 1.83,0.56 nfet_01v8
M$5 11 4 8 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=68250000000P
+ PS=1820000U PD=860000U
* device instance $6 r0 *1 2.19,0.56 nfet_01v8
M$6 9 5 11 10 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=234000000000P
+ PS=860000U PD=2020000U
* device instance $7 r0 *1 0.47,0.56 nfet_01v8
M$7 12 2 9 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=74750000000P
+ PS=1820000U PD=880000U
* device instance $8 r0 *1 0.85,0.56 nfet_01v8
M$8 8 3 12 10 nfet_01v8 L=150000U W=650000U AS=74750000000P AD=169000000000P
+ PS=880000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22oi_1

* cell sky130_fd_sc_hd__nor2_1
* pin VPB
* pin A
* pin B
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor2_1 1 2 3 4 5 6 7
* net 1 VPB
* net 2 A
* net 3 B
* net 4 Y
* net 5 VGND
* net 6 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 3 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=105000000000P PS=2520000U PD=1210000U
* device instance $2 r0 *1 0.83,1.985 pfet_01v8_hvt
M$2 6 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $3 r0 *1 0.47,0.56 nfet_01v8
M$3 4 3 5 7 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $4 r0 *1 0.89,0.56 nfet_01v8
M$4 5 2 4 7 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2_1

* cell sky130_fd_sc_hd__nand2b_1
* pin VPB
* pin B
* pin A_N
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nand2b_1 1 2 4 5 6 7 8
* net 1 VPB
* net 2 B
* net 4 A_N
* net 5 Y
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 7 4 3 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=145750000000P
+ PS=1360000U PD=1335000U
* device instance $2 r0 *1 0.955,1.985 pfet_01v8_hvt
M$2 5 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=145750000000P
+ AD=135000000000P PS=1335000U PD=1270000U
* device instance $3 r0 *1 1.375,1.985 pfet_01v8_hvt
M$3 7 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=265000000000P PS=1270000U PD=2530000U
* device instance $4 r0 *1 0.47,0.675 nfet_01v8
M$4 3 4 6 8 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
* device instance $5 r0 *1 0.955,0.56 nfet_01v8
M$5 9 2 6 8 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=87750000000P
+ PS=985000U PD=920000U
* device instance $6 r0 *1 1.375,0.56 nfet_01v8
M$6 5 3 9 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2b_1

* cell sky130_fd_sc_hd__dfrtp_1
* pin VGND
* pin RESET_B
* pin Q
* pin CLK
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__dfrtp_1 1 6 9 14 15 17 18 21
* net 1 VGND
* net 6 RESET_B
* net 9 Q
* net 14 CLK
* net 15 D
* net 17 VPWR
* net 18 VPB
* device instance $1 r0 *1 8.73,1.985 pfet_01v8_hvt
M$1 9 8 17 18 pfet_01v8_hvt L=150000U W=1000000U AS=301200000000P
+ AD=260000000000P PS=2660000U PD=2520000U
* device instance $2 r0 *1 5.35,2.065 pfet_01v8_hvt
M$2 16 5 17 18 pfet_01v8_hvt L=150000U W=840000U AS=218400000000P
+ AD=129150000000P PS=2200000U PD=1185000U
* device instance $3 r0 *1 5.845,2.275 pfet_01v8_hvt
M$3 7 2 16 18 pfet_01v8_hvt L=150000U W=420000U AS=129150000000P
+ AD=58800000000P PS=1185000U PD=700000U
* device instance $4 r0 *1 6.275,2.275 pfet_01v8_hvt
M$4 20 3 7 18 pfet_01v8_hvt L=150000U W=420000U AS=58800000000P AD=56700000000P
+ PS=700000U PD=690000U
* device instance $5 r0 *1 6.695,2.275 pfet_01v8_hvt
M$5 17 8 20 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=81900000000P PS=690000U PD=810000U
* device instance $6 r0 *1 7.235,2.275 pfet_01v8_hvt
M$6 8 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=81900000000P AD=56700000000P
+ PS=810000U PD=690000U
* device instance $7 r0 *1 7.655,2.275 pfet_01v8_hvt
M$7 17 7 8 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=113400000000P PS=690000U PD=1380000U
* device instance $8 r0 *1 2.225,2.275 pfet_01v8_hvt
M$8 4 15 17 18 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=65100000000P PS=1360000U PD=730000U
* device instance $9 r0 *1 2.685,2.275 pfet_01v8_hvt
M$9 5 3 4 18 pfet_01v8_hvt L=150000U W=420000U AS=65100000000P AD=72450000000P
+ PS=730000U PD=765000U
* device instance $10 r0 *1 3.18,2.275 pfet_01v8_hvt
M$10 19 2 5 18 pfet_01v8_hvt L=150000U W=420000U AS=72450000000P
+ AD=115500000000P PS=765000U PD=970000U
* device instance $11 r0 *1 3.88,2.275 pfet_01v8_hvt
M$11 17 16 19 18 pfet_01v8_hvt L=150000U W=420000U AS=115500000000P
+ AD=70350000000P PS=970000U PD=755000U
* device instance $12 r0 *1 4.365,2.275 pfet_01v8_hvt
M$12 19 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=70350000000P
+ AD=109200000000P PS=755000U PD=1360000U
* device instance $13 r0 *1 0.47,2.135 pfet_01v8_hvt
M$13 17 14 2 18 pfet_01v8_hvt L=150000U W=640000U AS=166400000000P
+ AD=86400000000P PS=1800000U PD=910000U
* device instance $14 r0 *1 0.89,2.135 pfet_01v8_hvt
M$14 3 2 17 18 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=166400000000P PS=910000U PD=1800000U
* device instance $15 r0 *1 8.73,0.56 nfet_01v8
M$15 9 8 1 21 nfet_01v8 L=150000U W=650000U AS=208700000000P AD=169000000000P
+ PS=2020000U PD=1820000U
* device instance $16 r0 *1 0.47,0.445 nfet_01v8
M$16 1 14 2 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $17 r0 *1 0.89,0.445 nfet_01v8
M$17 3 2 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $18 r0 *1 2.64,0.415 nfet_01v8
M$18 5 2 4 21 nfet_01v8 L=150000U W=360000U AS=66000000000P AD=59400000000P
+ PS=745000U PD=690000U
* device instance $19 r0 *1 3.12,0.415 nfet_01v8
M$19 12 3 5 21 nfet_01v8 L=150000U W=360000U AS=59400000000P AD=140100000000P
+ PS=690000U PD=1100000U
* device instance $20 r0 *1 5.465,0.415 nfet_01v8
M$20 7 3 16 21 nfet_01v8 L=150000U W=360000U AS=99900000000P AD=71100000000P
+ PS=985000U PD=755000U
* device instance $21 r0 *1 6.01,0.415 nfet_01v8
M$21 11 2 7 21 nfet_01v8 L=150000U W=360000U AS=71100000000P AD=66900000000P
+ PS=755000U PD=750000U
* device instance $22 r0 *1 2.165,0.445 nfet_01v8
M$22 4 15 1 21 nfet_01v8 L=150000U W=420000U AS=220500000000P AD=66000000000P
+ PS=1890000U PD=745000U
* device instance $23 r0 *1 3.95,0.445 nfet_01v8
M$23 13 16 12 21 nfet_01v8 L=150000U W=420000U AS=140100000000P AD=44100000000P
+ PS=1100000U PD=630000U
* device instance $24 r0 *1 4.31,0.445 nfet_01v8
M$24 1 6 13 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=134600000000P
+ PS=630000U PD=1150000U
* device instance $25 r0 *1 6.49,0.445 nfet_01v8
M$25 1 8 11 21 nfet_01v8 L=150000U W=420000U AS=66900000000P AD=124950000000P
+ PS=750000U PD=1015000U
* device instance $26 r0 *1 7.235,0.445 nfet_01v8
M$26 10 6 1 21 nfet_01v8 L=150000U W=420000U AS=124950000000P AD=64050000000P
+ PS=1015000U PD=725000U
* device instance $27 r0 *1 7.69,0.445 nfet_01v8
M$27 8 7 10 21 nfet_01v8 L=150000U W=420000U AS=64050000000P AD=109200000000P
+ PS=725000U PD=1360000U
* device instance $28 r0 *1 4.97,0.555 nfet_01v8
M$28 16 5 1 21 nfet_01v8 L=150000U W=640000U AS=134600000000P AD=99900000000P
+ PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_1

* cell sky130_fd_sc_hd__clkbuf_1
* pin VPB
* pin A
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_1 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 X
* net 5 VGND
* net 6 VPWR
* device instance $1 r0 *1 0.47,2.09 pfet_01v8_hvt
M$1 6 2 4 1 pfet_01v8_hvt L=150000U W=790000U AS=205400000000P AD=114550000000P
+ PS=2100000U PD=1080000U
* device instance $2 r0 *1 0.91,2.09 pfet_01v8_hvt
M$2 2 3 6 1 pfet_01v8_hvt L=150000U W=790000U AS=114550000000P AD=205400000000P
+ PS=1080000U PD=2100000U
* device instance $3 r0 *1 0.47,0.495 nfet_01v8
M$3 5 2 4 7 nfet_01v8 L=150000U W=520000U AS=135200000000P AD=75400000000P
+ PS=1560000U PD=810000U
* device instance $4 r0 *1 0.91,0.495 nfet_01v8
M$4 2 3 5 7 nfet_01v8 L=150000U W=520000U AS=75400000000P AD=135200000000P
+ PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

* cell sky130_fd_sc_hd__xnor2_1
* pin VPB
* pin B
* pin A
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__xnor2_1 1 2 3 4 5 7 9
* net 1 VPB
* net 2 B
* net 3 A
* net 4 Y
* net 5 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.51,1.985 pfet_01v8_hvt
M$1 8 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=300000000000P
+ AD=135000000000P PS=2600000U PD=1270000U
* device instance $2 r0 *1 0.93,1.985 pfet_01v8_hvt
M$2 5 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=365000000000P PS=1270000U PD=1730000U
* device instance $3 r0 *1 1.81,1.985 pfet_01v8_hvt
M$3 10 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=365000000000P
+ AD=105000000000P PS=1730000U PD=1210000U
* device instance $4 r0 *1 2.17,1.985 pfet_01v8_hvt
M$4 4 2 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=165000000000P PS=1210000U PD=1330000U
* device instance $5 r0 *1 2.65,1.985 pfet_01v8_hvt
M$5 5 8 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=360000000000P PS=1330000U PD=2720000U
* device instance $6 r0 *1 2.29,0.56 nfet_01v8
M$6 6 2 7 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 2.71,0.56 nfet_01v8
M$7 4 8 6 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=195000000000P
+ PS=920000U PD=1900000U
* device instance $8 r0 *1 0.57,0.56 nfet_01v8
M$8 11 2 8 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=68250000000P
+ PS=1820000U PD=860000U
* device instance $9 r0 *1 0.93,0.56 nfet_01v8
M$9 7 3 11 9 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=87750000000P
+ PS=860000U PD=920000U
* device instance $10 r0 *1 1.35,0.56 nfet_01v8
M$10 6 3 7 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__xnor2_1

* cell sky130_fd_sc_hd__o21ai_0
* pin VPB
* pin A1
* pin A2
* pin B1
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o21ai_0 1 2 3 4 5 6 8 9
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 B1
* net 5 VPWR
* net 6 Y
* net 8 VGND
* device instance $1 r0 *1 0.525,2.165 pfet_01v8_hvt
M$1 10 2 5 1 pfet_01v8_hvt L=150000U W=640000U AS=169600000000P AD=76800000000P
+ PS=1810000U PD=880000U
* device instance $2 r0 *1 0.915,2.165 pfet_01v8_hvt
M$2 6 3 10 1 pfet_01v8_hvt L=150000U W=640000U AS=76800000000P AD=89600000000P
+ PS=880000U PD=920000U
* device instance $3 r0 *1 1.345,2.165 pfet_01v8_hvt
M$3 5 4 6 1 pfet_01v8_hvt L=150000U W=640000U AS=89600000000P AD=182400000000P
+ PS=920000U PD=1850000U
* device instance $4 r0 *1 0.5,0.445 nfet_01v8
M$4 8 2 7 9 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=58800000000P
+ PS=1370000U PD=700000U
* device instance $5 r0 *1 0.93,0.445 nfet_01v8
M$5 7 3 8 9 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=58800000000P
+ PS=700000U PD=700000U
* device instance $6 r0 *1 1.36,0.445 nfet_01v8
M$6 6 4 7 9 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=111300000000P
+ PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__o21ai_0

* cell sky130_fd_sc_hd__nand2_1
* pin VPB
* pin A
* pin B
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__nand2_1 1 2 3 4 5 6 7
* net 1 VPB
* net 2 A
* net 3 B
* net 4 Y
* net 5 VPWR
* net 6 VGND
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 4 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.91,1.985 pfet_01v8_hvt
M$2 5 2 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $3 r0 *1 0.49,0.56 nfet_01v8
M$3 8 3 6 7 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $4 r0 *1 0.91,0.56 nfet_01v8
M$4 4 2 8 7 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2_1

* cell sky130_fd_sc_hd__mux2i_1
* pin VGND
* pin Y
* pin A0
* pin A1
* pin S
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2i_1 1 3 6 7 8 10 11 13
* net 1 VGND
* net 3 Y
* net 6 A0
* net 7 A1
* net 8 S
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 3.21,1.985 pfet_01v8_hvt
M$1 10 8 5 11 pfet_01v8_hvt L=150000U W=1000000U AS=290000000000P
+ AD=260000000000P PS=2580000U PD=2520000U
* device instance $2 r0 *1 0.49,1.985 pfet_01v8_hvt
M$2 3 6 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=152500000000P PS=2560000U PD=1305000U
* device instance $3 r0 *1 0.945,1.985 pfet_01v8_hvt
M$3 12 7 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=197500000000P PS=1305000U PD=1395000U
* device instance $4 r0 *1 1.49,1.985 pfet_01v8_hvt
M$4 10 5 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=197500000000P
+ AD=300000000000P PS=1395000U PD=1600000U
* device instance $5 r0 *1 2.24,1.985 pfet_01v8_hvt
M$5 9 8 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=300000000000P
+ AD=260000000000P PS=1600000U PD=2520000U
* device instance $6 r0 *1 3.21,0.56 nfet_01v8
M$6 1 8 5 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
* device instance $7 r0 *1 1.85,0.56 nfet_01v8
M$7 1 5 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 2.27,0.56 nfet_01v8
M$8 4 8 1 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 3 6 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $10 r0 *1 0.89,0.56 nfet_01v8
M$10 4 7 3 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=182000000000P
+ PS=920000U PD=1860000U
.ENDS sky130_fd_sc_hd__mux2i_1

* cell sky130_fd_sc_hd__clkbuf_4
* pin VPB
* pin A
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_4 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 VGND
* net 5 X
* net 6 VPWR
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 6 3 2 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=165000000000P PS=2530000U PD=1330000U
* device instance $2 r0 *1 0.955,1.985 pfet_01v8_hvt
M$2 5 2 6 1 pfet_01v8_hvt L=150000U W=4000000U AS=585000000000P
+ AD=720000000000P PS=5170000U PD=6440000U
* device instance $6 r0 *1 0.475,0.445 nfet_01v8
M$6 4 3 2 7 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=70350000000P
+ PS=1370000U PD=755000U
* device instance $7 r0 *1 0.96,0.445 nfet_01v8
M$7 5 2 4 7 nfet_01v8 L=150000U W=1680000U AS=246750000000P AD=298200000000P
+ PS=2855000U PD=3520000U
.ENDS sky130_fd_sc_hd__clkbuf_4
