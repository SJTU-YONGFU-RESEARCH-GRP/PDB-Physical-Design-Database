module clock_divider (clk_in,
    clk_out,
    rst_n,
    div_ratio,
    duty_cycle);
 input clk_in;
 output clk_out;
 input rst_n;
 input [7:0] div_ratio;
 input [7:0] duty_cycle;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire net81;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire net83;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire net2;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire net1;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk_in;
 wire clknet_1_0__leaf_clk_in;
 wire clknet_1_1__leaf_clk_in;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net82;
 wire net84;
 wire net85;
 wire net86;

 BUF_X2 _0882_ (.A(duty_cycle[7]),
    .Z(_0017_));
 BUF_X8 _0883_ (.A(net5),
    .Z(_0018_));
 AND2_X1 _0884_ (.A1(_0017_),
    .A2(net2),
    .ZN(_0748_));
 BUF_X2 _0885_ (.A(duty_cycle[6]),
    .Z(_0019_));
 CLKBUF_X1 hold71 (.A(rst_n),
    .Z(net81));
 AND2_X1 _0887_ (.A1(_0019_),
    .A2(net6),
    .ZN(_0749_));
 AND2_X1 _0888_ (.A1(_0017_),
    .A2(net6),
    .ZN(_0745_));
 BUF_X2 _0889_ (.A(duty_cycle[5]),
    .Z(_0021_));
 AND2_X1 _0890_ (.A1(net2),
    .A2(_0021_),
    .ZN(_0754_));
 BUF_X2 _0891_ (.A(duty_cycle[4]),
    .Z(_0022_));
 AND2_X1 _0892_ (.A1(net6),
    .A2(_0022_),
    .ZN(_0755_));
 AND2_X1 _0893_ (.A1(net2),
    .A2(_0019_),
    .ZN(_0584_));
 BUF_X4 _0894_ (.A(div_ratio[5]),
    .Z(_0023_));
 AND2_X1 _0895_ (.A1(_0017_),
    .A2(_0023_),
    .ZN(_0585_));
 AND2_X1 _0896_ (.A1(net6),
    .A2(_0021_),
    .ZN(_0753_));
 BUF_X4 _0897_ (.A(duty_cycle[3]),
    .Z(_0024_));
 AND2_X1 _0898_ (.A1(_0018_),
    .A2(_0024_),
    .ZN(_0761_));
 BUF_X4 _0899_ (.A(duty_cycle[2]),
    .Z(_0025_));
 AND2_X1 _0900_ (.A1(net6),
    .A2(_0025_),
    .ZN(_0762_));
 AND2_X1 _0901_ (.A1(_0018_),
    .A2(_0022_),
    .ZN(_0756_));
 AND2_X1 _0902_ (.A1(_0021_),
    .A2(_0023_),
    .ZN(_0757_));
 AND2_X1 _0903_ (.A1(_0019_),
    .A2(_0023_),
    .ZN(_0596_));
 BUF_X8 _0904_ (.A(div_ratio[4]),
    .Z(_0026_));
 AND2_X1 _0905_ (.A1(_0017_),
    .A2(_0026_),
    .ZN(_0597_));
 AND2_X1 _0906_ (.A1(_0018_),
    .A2(_0025_),
    .ZN(_0629_));
 BUF_X8 _0907_ (.A(duty_cycle[1]),
    .Z(_0027_));
 AND2_X1 _0908_ (.A1(net6),
    .A2(_0027_),
    .ZN(_0630_));
 AND2_X1 _0909_ (.A1(_0022_),
    .A2(_0023_),
    .ZN(_0763_));
 AND2_X1 _0910_ (.A1(_0021_),
    .A2(_0026_),
    .ZN(_0764_));
 AND2_X1 _0911_ (.A1(_0019_),
    .A2(_0026_),
    .ZN(_0612_));
 BUF_X4 _0912_ (.A(net4),
    .Z(_0028_));
 AND2_X1 _0913_ (.A1(_0017_),
    .A2(_0028_),
    .ZN(_0613_));
 AND2_X1 _0914_ (.A1(_0023_),
    .A2(_0025_),
    .ZN(_0650_));
 AND2_X1 _0915_ (.A1(_0027_),
    .A2(_0018_),
    .ZN(_0651_));
 AND2_X1 _0916_ (.A1(_0022_),
    .A2(_0026_),
    .ZN(_0765_));
 AND2_X1 _0917_ (.A1(_0021_),
    .A2(_0028_),
    .ZN(_0766_));
 AND2_X1 _0918_ (.A1(_0025_),
    .A2(_0026_),
    .ZN(_0674_));
 AND2_X1 _0919_ (.A1(_0023_),
    .A2(_0027_),
    .ZN(_0675_));
 BUF_X2 _0920_ (.A(duty_cycle[0]),
    .Z(_0029_));
 AND2_X1 _0921_ (.A1(net6),
    .A2(_0029_),
    .ZN(_0653_));
 AND2_X1 _0922_ (.A1(_0022_),
    .A2(_0028_),
    .ZN(_0654_));
 BUF_X4 _0923_ (.A(net3),
    .Z(_0030_));
 AND2_X1 _0924_ (.A1(_0021_),
    .A2(_0030_),
    .ZN(_0655_));
 AND2_X1 _0925_ (.A1(_0019_),
    .A2(_0030_),
    .ZN(_0658_));
 BUF_X2 _0926_ (.A(div_ratio[1]),
    .Z(_0031_));
 AND2_X1 _0927_ (.A1(_0017_),
    .A2(_0031_),
    .ZN(_0659_));
 AND2_X1 _0928_ (.A1(_0025_),
    .A2(_0028_),
    .ZN(_0698_));
 AND2_X1 _0929_ (.A1(_0026_),
    .A2(_0027_),
    .ZN(_0699_));
 AND2_X1 _0930_ (.A1(_0018_),
    .A2(_0029_),
    .ZN(_0677_));
 AND2_X1 _0931_ (.A1(_0022_),
    .A2(_0030_),
    .ZN(_0678_));
 AND2_X1 _0932_ (.A1(_0021_),
    .A2(_0031_),
    .ZN(_0679_));
 AND2_X1 _0933_ (.A1(_0019_),
    .A2(_0031_),
    .ZN(_0682_));
 BUF_X2 _0934_ (.A(div_ratio[0]),
    .Z(_0032_));
 AND2_X1 _0935_ (.A1(_0017_),
    .A2(_0032_),
    .ZN(_0683_));
 AND2_X1 _0936_ (.A1(_0025_),
    .A2(_0030_),
    .ZN(_0719_));
 AND2_X1 _0937_ (.A1(_0027_),
    .A2(_0028_),
    .ZN(_0718_));
 AND2_X1 _0938_ (.A1(_0023_),
    .A2(_0029_),
    .ZN(_0703_));
 AND2_X1 _0939_ (.A1(_0022_),
    .A2(_0031_),
    .ZN(_0702_));
 AND2_X1 _0940_ (.A1(_0021_),
    .A2(_0032_),
    .ZN(_0701_));
 AND2_X1 _0941_ (.A1(_0019_),
    .A2(_0032_),
    .ZN(_0771_));
 NAND2_X1 _0942_ (.A1(_0024_),
    .A2(_0032_),
    .ZN(_0733_));
 AND2_X1 _0943_ (.A1(_0026_),
    .A2(_0029_),
    .ZN(_0773_));
 AND2_X1 _0944_ (.A1(_0022_),
    .A2(_0032_),
    .ZN(_0772_));
 AND2_X1 _0945_ (.A1(_0027_),
    .A2(_0031_),
    .ZN(_0791_));
 AND2_X1 _0946_ (.A1(_0025_),
    .A2(_0032_),
    .ZN(_0790_));
 AND2_X1 _0947_ (.A1(_0030_),
    .A2(_0029_),
    .ZN(_0800_));
 AND2_X1 _0948_ (.A1(_0029_),
    .A2(_0031_),
    .ZN(_0823_));
 AND2_X1 _0949_ (.A1(_0027_),
    .A2(_0032_),
    .ZN(_0822_));
 CLKBUF_X2 _0950_ (.A(_0752_),
    .Z(_0033_));
 INV_X2 _0951_ (.A(_0033_),
    .ZN(_0034_));
 CLKBUF_X2 _0952_ (.A(_0746_),
    .Z(_0035_));
 CLKBUF_X3 _0953_ (.A(_0760_),
    .Z(_0036_));
 INV_X1 _0954_ (.A(_0036_),
    .ZN(_0037_));
 NOR3_X2 _0955_ (.A1(_0034_),
    .A2(_0035_),
    .A3(_0037_),
    .ZN(_0038_));
 CLKBUF_X3 _0956_ (.A(_0770_),
    .Z(_0039_));
 BUF_X4 _0957_ (.A(_0805_),
    .Z(_0040_));
 NAND2_X2 _0958_ (.A1(_0039_),
    .A2(_0040_),
    .ZN(_0041_));
 CLKBUF_X3 _0959_ (.A(_0808_),
    .Z(_0042_));
 CLKBUF_X3 _0960_ (.A(_0812_),
    .Z(_0043_));
 BUF_X4 _0961_ (.A(_0809_),
    .Z(_0044_));
 AOI21_X4 _0962_ (.A(_0042_),
    .B1(_0043_),
    .B2(_0044_),
    .ZN(_0045_));
 BUF_X4 _0963_ (.A(_0813_),
    .Z(_0046_));
 NAND4_X4 _0964_ (.A1(_0039_),
    .A2(_0044_),
    .A3(_0040_),
    .A4(_0046_),
    .ZN(_0047_));
 BUF_X1 rebuffer71 (.A(_0265_),
    .Z(net83));
 BUF_X4 _0966_ (.A(_0777_),
    .Z(_0049_));
 AOI21_X4 _0967_ (.A(_0776_),
    .B1(net84),
    .B2(_0049_),
    .ZN(_0050_));
 OAI22_X4 _0968_ (.A1(_0041_),
    .A2(_0045_),
    .B1(_0047_),
    .B2(_0050_),
    .ZN(_0051_));
 BUF_X4 _0969_ (.A(_0783_),
    .Z(_0052_));
 AOI211_X4 _0970_ (.A(_0052_),
    .B(_0793_),
    .C1(_0741_),
    .C2(_0794_),
    .ZN(_0053_));
 BUF_X4 _0971_ (.A(_0816_),
    .Z(_0054_));
 CLKBUF_X3 _0972_ (.A(_0784_),
    .Z(_0055_));
 OAI211_X4 _0973_ (.A(_0054_),
    .B(_0049_),
    .C1(_0052_),
    .C2(_0055_),
    .ZN(_0056_));
 NOR3_X2 _0974_ (.A1(_0047_),
    .A2(_0053_),
    .A3(_0056_),
    .ZN(_0057_));
 OAI21_X2 _0975_ (.A(_0038_),
    .B1(_0051_),
    .B2(_0057_),
    .ZN(_0058_));
 INV_X1 _0976_ (.A(_0751_),
    .ZN(_0059_));
 BUF_X2 _0977_ (.A(_0759_),
    .Z(_0060_));
 OAI21_X1 _0978_ (.A(_0033_),
    .B1(_0036_),
    .B2(_0060_),
    .ZN(_0061_));
 AND3_X1 _0979_ (.A1(_0035_),
    .A2(_0059_),
    .A3(_0061_),
    .ZN(_0062_));
 NAND3_X1 _0980_ (.A1(_0039_),
    .A2(_0036_),
    .A3(_0804_),
    .ZN(_0063_));
 AOI21_X1 _0981_ (.A(_0060_),
    .B1(_0769_),
    .B2(_0036_),
    .ZN(_0064_));
 NAND2_X1 _0982_ (.A1(_0063_),
    .A2(_0064_),
    .ZN(_0065_));
 NOR2_X1 _0983_ (.A1(_0034_),
    .A2(_0035_),
    .ZN(_0066_));
 INV_X1 _0984_ (.A(_0035_),
    .ZN(_0067_));
 AOI221_X2 _0985_ (.A(_0062_),
    .B1(_0065_),
    .B2(_0066_),
    .C1(_0067_),
    .C2(_0751_),
    .ZN(_0068_));
 NAND4_X1 _0986_ (.A1(_0035_),
    .A2(_0059_),
    .A3(_0063_),
    .A4(_0064_),
    .ZN(_0069_));
 OR3_X2 _0987_ (.A1(_0057_),
    .A2(_0051_),
    .A3(_0069_),
    .ZN(_0070_));
 NAND3_X4 _0988_ (.A1(_0058_),
    .A2(_0068_),
    .A3(_0070_),
    .ZN(_0071_));
 OAI21_X2 _0989_ (.A(_0050_),
    .B1(_0056_),
    .B2(_0053_),
    .ZN(_0072_));
 XOR2_X2 _0990_ (.A(_0072_),
    .B(_0046_),
    .Z(_0073_));
 BUF_X4 _0991_ (.A(_0073_),
    .Z(_0074_));
 INV_X1 _0992_ (.A(_0049_),
    .ZN(_0075_));
 AOI211_X2 _0993_ (.A(_0815_),
    .B(_0052_),
    .C1(_0055_),
    .C2(_0742_),
    .ZN(_0076_));
 NOR2_X1 _0994_ (.A1(_0054_),
    .A2(_0815_),
    .ZN(_0077_));
 OR3_X2 _0995_ (.A1(_0075_),
    .A2(net34),
    .A3(_0077_),
    .ZN(_0078_));
 OAI21_X2 _0996_ (.A(_0075_),
    .B1(net34),
    .B2(_0077_),
    .ZN(_0079_));
 AND2_X2 _0997_ (.A1(_0078_),
    .A2(_0079_),
    .ZN(_0080_));
 AOI21_X4 _0998_ (.A(_0043_),
    .B1(_0776_),
    .B2(_0046_),
    .ZN(_0081_));
 XNOR2_X2 _0999_ (.A(_0044_),
    .B(_0081_),
    .ZN(_0082_));
 AND3_X2 _1000_ (.A1(_0074_),
    .A2(_0080_),
    .A3(_0082_),
    .ZN(_0083_));
 NAND2_X2 _1001_ (.A1(_0071_),
    .A2(_0083_),
    .ZN(_0084_));
 INV_X1 _1002_ (.A(_0060_),
    .ZN(_0085_));
 AOI21_X2 _1003_ (.A(_0769_),
    .B1(_0804_),
    .B2(_0039_),
    .ZN(_0086_));
 NAND3_X1 _1004_ (.A1(_0039_),
    .A2(_0040_),
    .A3(_0042_),
    .ZN(_0087_));
 AND4_X1 _1005_ (.A1(_0033_),
    .A2(_0085_),
    .A3(_0086_),
    .A4(_0087_),
    .ZN(_0088_));
 AND3_X1 _1006_ (.A1(_0039_),
    .A2(_0044_),
    .A3(_0040_),
    .ZN(_0089_));
 AND3_X1 _1007_ (.A1(_0034_),
    .A2(_0036_),
    .A3(_0089_),
    .ZN(_0090_));
 OAI211_X4 _1008_ (.A(_0049_),
    .B(_0046_),
    .C1(_0054_),
    .C2(net84),
    .ZN(_0091_));
 OAI21_X4 _1009_ (.A(_0081_),
    .B1(_0091_),
    .B2(net34),
    .ZN(_0092_));
 MUX2_X2 _1010_ (.A(_0088_),
    .B(_0090_),
    .S(_0092_),
    .Z(_0093_));
 NOR2_X1 _1011_ (.A1(_0033_),
    .A2(_0037_),
    .ZN(_0094_));
 NOR3_X1 _1012_ (.A1(_0034_),
    .A2(_0060_),
    .A3(_0089_),
    .ZN(_0095_));
 AND2_X1 _1013_ (.A1(_0086_),
    .A2(_0087_),
    .ZN(_0096_));
 MUX2_X2 _1014_ (.A(_0094_),
    .B(_0095_),
    .S(_0096_),
    .Z(_0097_));
 NOR3_X4 _1015_ (.A1(_0034_),
    .A2(_0036_),
    .A3(_0060_),
    .ZN(_0098_));
 NOR2_X2 _1016_ (.A1(_0033_),
    .A2(_0085_),
    .ZN(_0099_));
 OR4_X4 _1017_ (.A1(_0097_),
    .A2(_0093_),
    .A3(_0098_),
    .A4(_0099_),
    .ZN(_0100_));
 BUF_X8 clone2 (.A(net5),
    .Z(net2));
 OAI21_X2 _1019_ (.A(_0086_),
    .B1(_0045_),
    .B2(_0041_),
    .ZN(_0102_));
 INV_X1 _1020_ (.A(_0047_),
    .ZN(_0103_));
 AOI21_X4 _1021_ (.A(_0102_),
    .B1(_0072_),
    .B2(_0103_),
    .ZN(_0104_));
 XNOR2_X2 _1022_ (.A(_0036_),
    .B(_0104_),
    .ZN(_0105_));
 BUF_X4 _1023_ (.A(_0105_),
    .Z(_0106_));
 AOI21_X4 _1024_ (.A(_0804_),
    .B1(_0042_),
    .B2(_0040_),
    .ZN(_0107_));
 OAI211_X2 _1025_ (.A(_0081_),
    .B(_0107_),
    .C1(_0091_),
    .C2(net34),
    .ZN(_0108_));
 INV_X1 _1026_ (.A(_0039_),
    .ZN(_0109_));
 NAND2_X1 _1027_ (.A1(_0044_),
    .A2(_0040_),
    .ZN(_0110_));
 AOI21_X1 _1028_ (.A(_0109_),
    .B1(_0107_),
    .B2(_0110_),
    .ZN(_0111_));
 AND2_X1 _1029_ (.A1(_0044_),
    .A2(_0040_),
    .ZN(_0112_));
 NOR2_X1 _1030_ (.A1(_0039_),
    .A2(_0112_),
    .ZN(_0113_));
 OR2_X2 _1031_ (.A1(net34),
    .A2(_0091_),
    .ZN(_0114_));
 INV_X1 _1032_ (.A(_0043_),
    .ZN(_0115_));
 NAND2_X1 _1033_ (.A1(_0046_),
    .A2(_0776_),
    .ZN(_0116_));
 AND4_X1 _1034_ (.A1(_0109_),
    .A2(_0115_),
    .A3(_0116_),
    .A4(_0107_),
    .ZN(_0117_));
 AOI222_X2 _1035_ (.A1(_0108_),
    .A2(_0111_),
    .B1(_0113_),
    .B2(_0107_),
    .C1(_0114_),
    .C2(_0117_),
    .ZN(_0118_));
 BUF_X4 _1036_ (.A(_0118_),
    .Z(_0119_));
 NOR2_X1 _1037_ (.A1(_0042_),
    .A2(_0043_),
    .ZN(_0120_));
 OAI211_X2 _1038_ (.A(_0050_),
    .B(_0120_),
    .C1(_0053_),
    .C2(_0056_),
    .ZN(_0121_));
 INV_X1 _1039_ (.A(_0040_),
    .ZN(_0122_));
 INV_X1 _1040_ (.A(_0042_),
    .ZN(_0123_));
 OAI21_X1 _1041_ (.A(_0044_),
    .B1(_0046_),
    .B2(_0043_),
    .ZN(_0124_));
 AOI21_X1 _1042_ (.A(_0122_),
    .B1(_0123_),
    .B2(_0124_),
    .ZN(_0125_));
 NOR2_X1 _1043_ (.A1(_0040_),
    .A2(_0042_),
    .ZN(_0126_));
 AND3_X1 _1044_ (.A1(_0115_),
    .A2(_0050_),
    .A3(_0126_),
    .ZN(_0127_));
 OR2_X2 _1045_ (.A1(_0056_),
    .A2(_0053_),
    .ZN(_0128_));
 AOI222_X2 _1046_ (.A1(_0121_),
    .A2(_0125_),
    .B1(_0126_),
    .B2(_0124_),
    .C1(_0128_),
    .C2(_0127_),
    .ZN(_0129_));
 BUF_X4 _1047_ (.A(_0129_),
    .Z(_0130_));
 AND2_X4 _1048_ (.A1(_0130_),
    .A2(_0119_),
    .ZN(_0131_));
 NAND3_X4 _1049_ (.A1(net61),
    .A2(_0106_),
    .A3(net68),
    .ZN(_0132_));
 NOR2_X2 _1050_ (.A1(_0084_),
    .A2(_0132_),
    .ZN(_0133_));
 INV_X2 _1051_ (.A(_0133_),
    .ZN(_0825_));
 AND3_X1 _1052_ (.A1(_0058_),
    .A2(_0068_),
    .A3(_0070_),
    .ZN(_0134_));
 BUF_X4 _1053_ (.A(_0134_),
    .Z(_0135_));
 NAND3_X4 _1054_ (.A1(net35),
    .A2(_0080_),
    .A3(_0082_),
    .ZN(_0136_));
 NOR2_X2 _1055_ (.A1(_0135_),
    .A2(_0136_),
    .ZN(_0137_));
 NOR4_X4 _1056_ (.A1(_0097_),
    .A2(_0093_),
    .A3(_0098_),
    .A4(_0099_),
    .ZN(_0138_));
 XNOR2_X2 _1057_ (.A(_0037_),
    .B(_0104_),
    .ZN(_0139_));
 NAND2_X4 _1058_ (.A1(net23),
    .A2(_0119_),
    .ZN(_0140_));
 NOR3_X4 _1059_ (.A1(_0140_),
    .A2(_0139_),
    .A3(net14),
    .ZN(_0141_));
 INV_X1 _1060_ (.A(_0054_),
    .ZN(_0142_));
 NOR2_X2 _1061_ (.A1(_0055_),
    .A2(_0052_),
    .ZN(_0143_));
 OAI21_X4 _1062_ (.A(_0142_),
    .B1(_0053_),
    .B2(_0143_),
    .ZN(_0144_));
 OR3_X4 _1063_ (.A1(_0142_),
    .A2(_0053_),
    .A3(_0143_),
    .ZN(_0145_));
 AND4_X4 _1064_ (.A1(_0078_),
    .A2(_0079_),
    .A3(_0144_),
    .A4(_0145_),
    .ZN(_0146_));
 AND3_X4 _1065_ (.A1(net35),
    .A2(_0082_),
    .A3(_0146_),
    .ZN(_0147_));
 NAND4_X4 _1066_ (.A1(_0131_),
    .A2(_0105_),
    .A3(_0100_),
    .A4(_0147_),
    .ZN(_0148_));
 AOI22_X4 _1067_ (.A1(net12),
    .A2(_0137_),
    .B1(net86),
    .B2(_0135_),
    .ZN(_0149_));
 INV_X1 _1068_ (.A(_0149_),
    .ZN(_0829_));
 NAND2_X2 _1069_ (.A1(_0106_),
    .A2(net68),
    .ZN(_0150_));
 NAND3_X2 _1070_ (.A1(_0071_),
    .A2(_0083_),
    .A3(net61),
    .ZN(_0151_));
 NAND2_X1 _1071_ (.A1(_0135_),
    .A2(_0147_),
    .ZN(_0152_));
 AOI21_X4 _1072_ (.A(_0150_),
    .B1(_0151_),
    .B2(_0152_),
    .ZN(_0153_));
 NAND3_X4 _1073_ (.A1(net35),
    .A2(_0082_),
    .A3(_0146_),
    .ZN(_0154_));
 NOR2_X4 _1074_ (.A1(_0140_),
    .A2(_0154_),
    .ZN(_0155_));
 AOI21_X4 _1075_ (.A(net62),
    .B1(_0106_),
    .B2(_0155_),
    .ZN(_0156_));
 NOR2_X4 _1076_ (.A1(_0153_),
    .A2(_0156_),
    .ZN(_0157_));
 AND2_X1 _1077_ (.A1(_0144_),
    .A2(_0145_),
    .ZN(_0158_));
 CLKBUF_X3 _1078_ (.A(_0158_),
    .Z(_0159_));
 XNOR2_X2 _1079_ (.A(_0149_),
    .B(_0159_),
    .ZN(_0160_));
 BUF_X4 _1080_ (.A(_0071_),
    .Z(_0161_));
 AND4_X1 _1081_ (.A1(_0074_),
    .A2(_0080_),
    .A3(_0082_),
    .A4(_0119_),
    .ZN(_0162_));
 NAND4_X2 _1082_ (.A1(_0161_),
    .A2(net61),
    .A3(_0106_),
    .A4(_0162_),
    .ZN(_0163_));
 BUF_X4 _1083_ (.A(_0135_),
    .Z(_0164_));
 OAI21_X1 _1084_ (.A(_0164_),
    .B1(net19),
    .B2(_0139_),
    .ZN(_0165_));
 NAND3_X2 _1085_ (.A1(_0155_),
    .A2(_0163_),
    .A3(_0165_),
    .ZN(_0166_));
 AOI221_X2 _1086_ (.A(_0804_),
    .B1(_0092_),
    .B2(_0112_),
    .C1(_0042_),
    .C2(_0040_),
    .ZN(_0167_));
 XNOR2_X2 _1087_ (.A(_0109_),
    .B(_0167_),
    .ZN(_0168_));
 NAND4_X4 _1088_ (.A1(_0074_),
    .A2(_0082_),
    .A3(_0130_),
    .A4(_0146_),
    .ZN(_0169_));
 OAI21_X2 _1089_ (.A(_0168_),
    .B1(_0169_),
    .B2(_0164_),
    .ZN(_0170_));
 NAND4_X2 _1090_ (.A1(_0161_),
    .A2(_0083_),
    .A3(net61),
    .A4(net69),
    .ZN(_0171_));
 XOR2_X2 _1091_ (.A(_0055_),
    .B(_0742_),
    .Z(_0172_));
 AND4_X2 _1092_ (.A1(_0106_),
    .A2(_0170_),
    .A3(_0171_),
    .A4(_0172_),
    .ZN(_0173_));
 NAND2_X4 _1093_ (.A1(_0166_),
    .A2(_0173_),
    .ZN(_0174_));
 NOR2_X4 _1094_ (.A1(net17),
    .A2(_0139_),
    .ZN(_0175_));
 NAND2_X1 _1095_ (.A1(_0130_),
    .A2(_0159_),
    .ZN(_0176_));
 AOI211_X4 _1096_ (.A(_0136_),
    .B(_0168_),
    .C1(_0176_),
    .C2(_0135_),
    .ZN(_0177_));
 AND3_X1 _1097_ (.A1(_0074_),
    .A2(_0080_),
    .A3(_0130_),
    .ZN(_0178_));
 NAND2_X4 _1098_ (.A1(_0144_),
    .A2(_0145_),
    .ZN(_0179_));
 OAI21_X2 _1099_ (.A(_0178_),
    .B1(_0179_),
    .B2(_0135_),
    .ZN(_0180_));
 NAND2_X1 _1100_ (.A1(_0078_),
    .A2(_0079_),
    .ZN(_0181_));
 AND3_X1 _1101_ (.A1(_0074_),
    .A2(_0181_),
    .A3(_0130_),
    .ZN(_0182_));
 NAND3_X2 _1102_ (.A1(_0161_),
    .A2(_0159_),
    .A3(_0182_),
    .ZN(_0183_));
 AOI22_X4 _1103_ (.A1(_0175_),
    .A2(_0177_),
    .B1(_0180_),
    .B2(_0183_),
    .ZN(_0184_));
 NAND2_X1 _1104_ (.A1(_0080_),
    .A2(_0159_),
    .ZN(_0185_));
 XNOR2_X2 _1105_ (.A(_0044_),
    .B(_0092_),
    .ZN(_0186_));
 INV_X1 _1106_ (.A(_0186_),
    .ZN(_0187_));
 NOR3_X2 _1107_ (.A1(_0164_),
    .A2(_0185_),
    .A3(_0187_),
    .ZN(_0188_));
 NAND2_X1 _1108_ (.A1(_0164_),
    .A2(_0187_),
    .ZN(_0189_));
 NOR4_X4 _1109_ (.A1(_0140_),
    .A2(_0139_),
    .A3(net15),
    .A4(_0154_),
    .ZN(_0190_));
 OAI222_X2 _1110_ (.A1(_0084_),
    .A2(_0132_),
    .B1(_0146_),
    .B2(_0186_),
    .C1(_0189_),
    .C2(_0190_),
    .ZN(_0191_));
 OAI21_X4 _1111_ (.A(_0184_),
    .B1(_0191_),
    .B2(_0188_),
    .ZN(_0192_));
 NOR3_X4 _1112_ (.A1(net63),
    .A2(_0174_),
    .A3(net36),
    .ZN(_0193_));
 NOR2_X1 _1113_ (.A1(_0157_),
    .A2(_0193_),
    .ZN(_0832_));
 NOR2_X1 _1114_ (.A1(_0139_),
    .A2(_0140_),
    .ZN(_0194_));
 NOR3_X2 _1115_ (.A1(_0135_),
    .A2(_0136_),
    .A3(net16),
    .ZN(_0195_));
 NOR2_X1 _1116_ (.A1(_0071_),
    .A2(_0154_),
    .ZN(_0196_));
 OAI21_X4 _1117_ (.A(_0194_),
    .B1(_0195_),
    .B2(_0196_),
    .ZN(_0197_));
 OAI21_X4 _1118_ (.A(net14),
    .B1(_0150_),
    .B2(_0154_),
    .ZN(_0198_));
 NAND2_X1 _1119_ (.A1(net61),
    .A2(_0106_),
    .ZN(_0199_));
 AND2_X1 _1120_ (.A1(_0083_),
    .A2(net1),
    .ZN(_0200_));
 NOR2_X1 _1121_ (.A1(_0057_),
    .A2(_0051_),
    .ZN(_0201_));
 NOR3_X1 _1122_ (.A1(_0067_),
    .A2(_0751_),
    .A3(_0065_),
    .ZN(_0202_));
 AND4_X1 _1123_ (.A1(_0201_),
    .A2(_0202_),
    .A3(_0144_),
    .A4(_0145_),
    .ZN(_0203_));
 NAND3_X1 _1124_ (.A1(_0038_),
    .A2(_0144_),
    .A3(_0145_),
    .ZN(_0204_));
 OAI22_X2 _1125_ (.A1(_0068_),
    .A2(_0179_),
    .B1(_0204_),
    .B2(_0201_),
    .ZN(_0205_));
 XNOR2_X2 _1126_ (.A(_0055_),
    .B(_0742_),
    .ZN(_0206_));
 AND4_X1 _1127_ (.A1(_0058_),
    .A2(_0068_),
    .A3(_0070_),
    .A4(_0179_),
    .ZN(_0207_));
 NOR4_X4 _1128_ (.A1(_0207_),
    .A2(_0205_),
    .A3(_0206_),
    .A4(_0203_),
    .ZN(_0208_));
 AND4_X1 _1129_ (.A1(_0199_),
    .A2(_0119_),
    .A3(_0200_),
    .A4(_0208_),
    .ZN(_0209_));
 AND3_X2 _1130_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0209_),
    .ZN(_0210_));
 NAND3_X1 _1131_ (.A1(net61),
    .A2(net68),
    .A3(_0147_),
    .ZN(_0211_));
 AOI21_X2 _1132_ (.A(_0161_),
    .B1(_0106_),
    .B2(_0211_),
    .ZN(_0212_));
 OAI211_X2 _1133_ (.A(_0161_),
    .B(_0083_),
    .C1(net61),
    .C2(_0159_),
    .ZN(_0213_));
 OAI22_X2 _1134_ (.A1(_0106_),
    .A2(_0155_),
    .B1(_0150_),
    .B2(_0213_),
    .ZN(_0214_));
 NOR2_X2 _1135_ (.A1(_0212_),
    .A2(_0214_),
    .ZN(_0215_));
 NOR2_X2 _1136_ (.A1(_0210_),
    .A2(_0215_),
    .ZN(_0216_));
 NOR2_X4 _1137_ (.A1(_0193_),
    .A2(_0216_),
    .ZN(_0217_));
 XNOR2_X1 _1138_ (.A(_0179_),
    .B(_0149_),
    .ZN(_0218_));
 AOI21_X1 _1139_ (.A(_0186_),
    .B1(net12),
    .B2(_0137_),
    .ZN(_0219_));
 AND2_X1 _1140_ (.A1(_0074_),
    .A2(_0146_),
    .ZN(_0220_));
 OAI221_X2 _1141_ (.A(_0220_),
    .B1(_0190_),
    .B2(_0161_),
    .C1(_0084_),
    .C2(_0132_),
    .ZN(_0221_));
 MUX2_X1 _1142_ (.A(_0186_),
    .B(_0219_),
    .S(_0221_),
    .Z(_0222_));
 BUF_X4 _1143_ (.A(_0222_),
    .Z(_0223_));
 BUF_X4 _1144_ (.A(_0743_),
    .Z(_0224_));
 OAI21_X2 _1145_ (.A(_0080_),
    .B1(_0179_),
    .B2(_0164_),
    .ZN(_0225_));
 NAND3_X2 _1146_ (.A1(_0161_),
    .A2(_0181_),
    .A3(_0159_),
    .ZN(_0226_));
 AOI21_X4 _1147_ (.A(_0136_),
    .B1(_0179_),
    .B2(_0135_),
    .ZN(_0227_));
 AOI22_X4 _1148_ (.A1(_0225_),
    .A2(_0226_),
    .B1(_0227_),
    .B2(net13),
    .ZN(_0228_));
 AND3_X2 _1149_ (.A1(_0224_),
    .A2(_0206_),
    .A3(_0228_),
    .ZN(_0229_));
 NAND3_X1 _1150_ (.A1(_0218_),
    .A2(_0223_),
    .A3(_0229_),
    .ZN(_0230_));
 BUF_X4 _1151_ (.A(_0218_),
    .Z(_0231_));
 AND3_X2 _1152_ (.A1(_0224_),
    .A2(_0172_),
    .A3(_0228_),
    .ZN(_0232_));
 NAND3_X1 _1153_ (.A1(_0231_),
    .A2(_0223_),
    .A3(_0232_),
    .ZN(_0233_));
 AND3_X1 _1154_ (.A1(_0155_),
    .A2(_0163_),
    .A3(_0165_),
    .ZN(_0234_));
 NAND4_X4 _1155_ (.A1(_0106_),
    .A2(_0170_),
    .A3(_0171_),
    .A4(_0172_),
    .ZN(_0235_));
 NOR2_X2 _1156_ (.A1(_0234_),
    .A2(_0235_),
    .ZN(_0236_));
 NAND3_X1 _1157_ (.A1(_0161_),
    .A2(_0146_),
    .A3(_0186_),
    .ZN(_0237_));
 NOR2_X1 _1158_ (.A1(_0071_),
    .A2(_0186_),
    .ZN(_0238_));
 AOI222_X2 _1159_ (.A1(_0137_),
    .A2(_0141_),
    .B1(_0185_),
    .B2(_0187_),
    .C1(_0148_),
    .C2(_0238_),
    .ZN(_0239_));
 AOI222_X2 _1160_ (.A1(_0175_),
    .A2(_0177_),
    .B1(_0180_),
    .B2(_0183_),
    .C1(_0239_),
    .C2(_0237_),
    .ZN(_0240_));
 AOI21_X4 _1161_ (.A(_0157_),
    .B1(net78),
    .B2(_0236_),
    .ZN(_0241_));
 MUX2_X2 _1162_ (.A(_0230_),
    .B(_0233_),
    .S(_0241_),
    .Z(_0242_));
 NOR2_X1 _1163_ (.A1(_0164_),
    .A2(_0169_),
    .ZN(_0243_));
 NAND2_X1 _1164_ (.A1(_0164_),
    .A2(_0179_),
    .ZN(_0244_));
 OAI22_X2 _1165_ (.A1(net18),
    .A2(_0139_),
    .B1(_0179_),
    .B2(_0164_),
    .ZN(_0245_));
 NAND3_X2 _1166_ (.A1(_0200_),
    .A2(_0244_),
    .A3(_0245_),
    .ZN(_0246_));
 MUX2_X2 _1167_ (.A(_0243_),
    .B(_0246_),
    .S(net30),
    .Z(_0247_));
 NAND2_X2 _1168_ (.A1(_0161_),
    .A2(_0147_),
    .ZN(_0248_));
 OR2_X1 _1169_ (.A1(net1),
    .A2(_0248_),
    .ZN(_0249_));
 NAND2_X1 _1170_ (.A1(net1),
    .A2(_0248_),
    .ZN(_0250_));
 AND3_X1 _1171_ (.A1(_0175_),
    .A2(_0119_),
    .A3(_0227_),
    .ZN(_0251_));
 OAI21_X2 _1172_ (.A(_0249_),
    .B1(_0250_),
    .B2(_0251_),
    .ZN(_0252_));
 NAND2_X1 _1173_ (.A1(_0164_),
    .A2(_0154_),
    .ZN(_0253_));
 AOI21_X4 _1174_ (.A(_0136_),
    .B1(net33),
    .B2(_0253_),
    .ZN(_0254_));
 AND4_X2 _1175_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0208_),
    .A4(_0254_),
    .ZN(_0255_));
 AOI22_X4 _1176_ (.A1(_0197_),
    .A2(_0198_),
    .B1(_0166_),
    .B2(_0173_),
    .ZN(_0256_));
 NAND3_X2 _1177_ (.A1(_0184_),
    .A2(_0208_),
    .A3(_0254_),
    .ZN(_0257_));
 OAI221_X2 _1178_ (.A(_0247_),
    .B1(_0252_),
    .B2(_0255_),
    .C1(_0256_),
    .C2(_0257_),
    .ZN(_0258_));
 OAI221_X2 _1179_ (.A(_0146_),
    .B1(net22),
    .B2(_0161_),
    .C1(_0084_),
    .C2(_0132_),
    .ZN(_0259_));
 XOR2_X2 _1180_ (.A(_0074_),
    .B(_0259_),
    .Z(_0260_));
 OAI21_X2 _1181_ (.A(_0080_),
    .B1(_0084_),
    .B2(_0132_),
    .ZN(_0261_));
 OR3_X1 _1182_ (.A1(_0153_),
    .A2(_0156_),
    .A3(_0261_),
    .ZN(_0262_));
 NAND2_X1 _1183_ (.A1(_0159_),
    .A2(_0172_),
    .ZN(_0263_));
 NAND2_X1 _1184_ (.A1(_0179_),
    .A2(_0172_),
    .ZN(_0264_));
 MUX2_X2 _1185_ (.A(_0263_),
    .B(_0264_),
    .S(_0149_),
    .Z(_0265_));
 OAI22_X4 _1186_ (.A1(_0133_),
    .A2(_0260_),
    .B1(_0262_),
    .B2(_0265_),
    .ZN(_0266_));
 NAND2_X1 _1187_ (.A1(_0074_),
    .A2(_0228_),
    .ZN(_0267_));
 OR2_X2 _1188_ (.A1(_0265_),
    .A2(_0267_),
    .ZN(_0268_));
 OAI21_X4 _1189_ (.A(_0266_),
    .B1(net25),
    .B2(_0268_),
    .ZN(_0269_));
 NOR3_X4 _1190_ (.A1(net39),
    .A2(_0258_),
    .A3(net29),
    .ZN(_0270_));
 NOR2_X1 _1191_ (.A1(_0217_),
    .A2(_0270_),
    .ZN(_0835_));
 NOR3_X2 _1192_ (.A1(_0164_),
    .A2(net30),
    .A3(_0169_),
    .ZN(_0271_));
 AOI21_X4 _1193_ (.A(_0271_),
    .B1(_0246_),
    .B2(net30),
    .ZN(_0272_));
 AND3_X2 _1194_ (.A1(_0184_),
    .A2(_0208_),
    .A3(_0254_),
    .ZN(_0273_));
 OAI22_X4 _1195_ (.A1(_0153_),
    .A2(_0156_),
    .B1(_0234_),
    .B2(_0235_),
    .ZN(_0274_));
 NAND2_X1 _1196_ (.A1(_0273_),
    .A2(_0274_),
    .ZN(_0275_));
 XNOR2_X2 _1197_ (.A(_0272_),
    .B(_0275_),
    .ZN(_0276_));
 NAND2_X1 _1198_ (.A1(_0231_),
    .A2(_0229_),
    .ZN(_0277_));
 NAND2_X1 _1199_ (.A1(_0231_),
    .A2(_0232_),
    .ZN(_0278_));
 MUX2_X2 _1200_ (.A(_0277_),
    .B(_0278_),
    .S(_0241_),
    .Z(_0279_));
 OAI221_X2 _1201_ (.A(net79),
    .B1(_0255_),
    .B2(_0252_),
    .C1(_0256_),
    .C2(_0257_),
    .ZN(_0280_));
 AOI21_X1 _1202_ (.A(_0140_),
    .B1(_0248_),
    .B2(net14),
    .ZN(_0281_));
 AOI21_X1 _1203_ (.A(_0139_),
    .B1(_0227_),
    .B2(_0281_),
    .ZN(_0282_));
 NOR3_X1 _1204_ (.A1(_0106_),
    .A2(_0140_),
    .A3(_0248_),
    .ZN(_0283_));
 OAI33_X1 _1205_ (.A1(_0160_),
    .A2(_0174_),
    .A3(_0192_),
    .B1(_0210_),
    .B2(_0282_),
    .B3(_0283_),
    .ZN(_0284_));
 OR2_X2 _1206_ (.A1(net10),
    .A2(_0255_),
    .ZN(_0285_));
 OR4_X2 _1207_ (.A1(_0279_),
    .A2(_0269_),
    .A3(_0280_),
    .A4(_0285_),
    .ZN(_0286_));
 AOI21_X4 _1208_ (.A(_0270_),
    .B1(_0286_),
    .B2(_0276_),
    .ZN(_0287_));
 NOR2_X4 _1209_ (.A1(_0224_),
    .A2(_0217_),
    .ZN(_0288_));
 INV_X1 _1210_ (.A(_0224_),
    .ZN(_0289_));
 NAND4_X4 _1211_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0208_),
    .A4(_0254_),
    .ZN(_0290_));
 NOR2_X1 _1212_ (.A1(net1),
    .A2(_0248_),
    .ZN(_0291_));
 AND2_X1 _1213_ (.A1(net1),
    .A2(_0248_),
    .ZN(_0292_));
 NAND3_X2 _1214_ (.A1(_0175_),
    .A2(net30),
    .A3(_0227_),
    .ZN(_0293_));
 AOI21_X4 _1215_ (.A(_0291_),
    .B1(_0292_),
    .B2(_0293_),
    .ZN(_0294_));
 AOI22_X4 _1216_ (.A1(_0290_),
    .A2(_0294_),
    .B1(_0274_),
    .B2(_0273_),
    .ZN(_0295_));
 NAND3_X1 _1217_ (.A1(_0224_),
    .A2(_0247_),
    .A3(_0295_),
    .ZN(_0296_));
 OAI33_X1 _1218_ (.A1(_0289_),
    .A2(_0193_),
    .A3(_0216_),
    .B1(_0269_),
    .B2(_0242_),
    .B3(_0296_),
    .ZN(_0297_));
 CLKBUF_X3 _1219_ (.A(_0828_),
    .Z(_0298_));
 NOR3_X4 _1220_ (.A1(_0153_),
    .A2(_0156_),
    .A3(_0206_),
    .ZN(_0299_));
 NOR2_X2 _1221_ (.A1(_0157_),
    .A2(_0172_),
    .ZN(_0300_));
 NOR3_X4 _1222_ (.A1(_0193_),
    .A2(_0299_),
    .A3(_0300_),
    .ZN(_0301_));
 NAND2_X2 _1223_ (.A1(_0298_),
    .A2(_0301_),
    .ZN(_0302_));
 OR3_X4 _1224_ (.A1(net9),
    .A2(_0302_),
    .A3(_0288_),
    .ZN(_0303_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 AND3_X1 _1226_ (.A1(_0231_),
    .A2(_0223_),
    .A3(_0229_),
    .ZN(_0305_));
 AND3_X1 _1227_ (.A1(_0231_),
    .A2(_0223_),
    .A3(_0232_),
    .ZN(_0306_));
 MUX2_X2 _1228_ (.A(_0305_),
    .B(_0306_),
    .S(net50),
    .Z(_0307_));
 XNOR2_X2 _1229_ (.A(_0074_),
    .B(_0259_),
    .ZN(_0308_));
 NOR3_X2 _1230_ (.A1(_0153_),
    .A2(_0156_),
    .A3(_0261_),
    .ZN(_0309_));
 NOR2_X1 _1231_ (.A1(_0179_),
    .A2(_0206_),
    .ZN(_0310_));
 NOR2_X1 _1232_ (.A1(_0159_),
    .A2(_0206_),
    .ZN(_0311_));
 MUX2_X2 _1233_ (.A(_0310_),
    .B(_0311_),
    .S(_0149_),
    .Z(_0312_));
 AOI22_X4 _1234_ (.A1(_0825_),
    .A2(_0308_),
    .B1(_0309_),
    .B2(_0312_),
    .ZN(_0313_));
 NAND2_X2 _1235_ (.A1(_0197_),
    .A2(_0198_),
    .ZN(_0314_));
 OAI21_X4 _1236_ (.A(_0314_),
    .B1(_0174_),
    .B2(net36),
    .ZN(_0315_));
 NOR2_X2 _1237_ (.A1(_0265_),
    .A2(_0267_),
    .ZN(_0316_));
 AOI211_X2 _1238_ (.A(_0313_),
    .B(_0258_),
    .C1(_0315_),
    .C2(_0316_),
    .ZN(_0317_));
 NAND3_X1 _1239_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0209_),
    .ZN(_0318_));
 OR2_X1 _1240_ (.A1(_0212_),
    .A2(_0214_),
    .ZN(_0319_));
 AOI21_X2 _1241_ (.A(_0289_),
    .B1(_0318_),
    .B2(_0319_),
    .ZN(_0320_));
 OAI221_X2 _1242_ (.A(_0160_),
    .B1(_0320_),
    .B2(_0299_),
    .C1(_0172_),
    .C2(_0157_),
    .ZN(_0321_));
 NAND2_X1 _1243_ (.A1(_0236_),
    .A2(net78),
    .ZN(_0322_));
 NOR2_X1 _1244_ (.A1(_0160_),
    .A2(_0299_),
    .ZN(_0323_));
 OAI21_X2 _1245_ (.A(_0224_),
    .B1(_0210_),
    .B2(_0215_),
    .ZN(_0324_));
 OAI211_X2 _1246_ (.A(_0322_),
    .B(_0323_),
    .C1(_0300_),
    .C2(_0324_),
    .ZN(_0325_));
 AOI22_X4 _1247_ (.A1(_0307_),
    .A2(_0317_),
    .B1(_0321_),
    .B2(_0325_),
    .ZN(_0326_));
 AOI21_X4 _1248_ (.A(_0313_),
    .B1(_0316_),
    .B2(_0315_),
    .ZN(_0327_));
 AOI21_X2 _1249_ (.A(_0228_),
    .B1(_0312_),
    .B2(_0157_),
    .ZN(_0328_));
 NOR2_X2 _1250_ (.A1(_0265_),
    .A2(_0261_),
    .ZN(_0329_));
 AOI21_X4 _1251_ (.A(_0328_),
    .B1(_0329_),
    .B2(_0315_),
    .ZN(_0330_));
 AND3_X1 _1252_ (.A1(_0295_),
    .A2(_0327_),
    .A3(_0330_),
    .ZN(_0331_));
 AND2_X1 _1253_ (.A1(_0231_),
    .A2(_0229_),
    .ZN(_0332_));
 AND2_X1 _1254_ (.A1(_0231_),
    .A2(_0232_),
    .ZN(_0333_));
 MUX2_X2 _1255_ (.A(_0332_),
    .B(_0333_),
    .S(net26),
    .Z(_0334_));
 NAND3_X1 _1256_ (.A1(_0231_),
    .A2(_0236_),
    .A3(net78),
    .ZN(_0335_));
 XNOR2_X1 _1257_ (.A(_0186_),
    .B(net82),
    .ZN(_0336_));
 NAND4_X1 _1258_ (.A1(_0074_),
    .A2(_0197_),
    .A3(_0198_),
    .A4(_0228_),
    .ZN(_0337_));
 OAI22_X2 _1259_ (.A1(_0133_),
    .A2(_0336_),
    .B1(net83),
    .B2(_0337_),
    .ZN(_0338_));
 NAND3_X2 _1260_ (.A1(_0335_),
    .A2(_0338_),
    .A3(_0290_),
    .ZN(_0339_));
 OAI211_X2 _1261_ (.A(net79),
    .B(_0272_),
    .C1(_0252_),
    .C2(_0255_),
    .ZN(_0340_));
 OAI221_X2 _1262_ (.A(net10),
    .B1(_0272_),
    .B2(_0280_),
    .C1(_0340_),
    .C2(_0275_),
    .ZN(_0341_));
 AND3_X1 _1263_ (.A1(_0334_),
    .A2(_0339_),
    .A3(_0341_),
    .ZN(_0342_));
 OAI211_X2 _1264_ (.A(net80),
    .B(_0247_),
    .C1(_0256_),
    .C2(_0257_),
    .ZN(_0343_));
 NAND4_X1 _1265_ (.A1(_0223_),
    .A2(_0273_),
    .A3(_0272_),
    .A4(_0274_),
    .ZN(_0344_));
 NAND3_X1 _1266_ (.A1(net10),
    .A2(_0343_),
    .A3(_0344_),
    .ZN(_0345_));
 AOI21_X2 _1267_ (.A(_0339_),
    .B1(_0345_),
    .B2(_0334_),
    .ZN(_0346_));
 OAI211_X4 _1268_ (.A(_0326_),
    .B(_0331_),
    .C1(_0342_),
    .C2(_0346_),
    .ZN(_0347_));
 NOR2_X1 _1269_ (.A1(net45),
    .A2(_0347_),
    .ZN(_0348_));
 NOR2_X2 _1270_ (.A1(_0287_),
    .A2(_0348_),
    .ZN(_0838_));
 NOR2_X2 _1271_ (.A1(net27),
    .A2(_0280_),
    .ZN(_0349_));
 AND3_X1 _1272_ (.A1(net10),
    .A2(_0343_),
    .A3(_0344_),
    .ZN(_0350_));
 NOR2_X2 _1273_ (.A1(_0279_),
    .A2(_0350_),
    .ZN(_0351_));
 OR3_X2 _1274_ (.A1(_0242_),
    .A2(_0269_),
    .A3(_0285_),
    .ZN(_0352_));
 INV_X1 _1275_ (.A(_0295_),
    .ZN(_0353_));
 AOI22_X4 _1276_ (.A1(_0349_),
    .A2(_0351_),
    .B1(_0352_),
    .B2(_0353_),
    .ZN(_0354_));
 NAND3_X2 _1277_ (.A1(_0334_),
    .A2(_0327_),
    .A3(_0341_),
    .ZN(_0355_));
 OAI21_X2 _1278_ (.A(net27),
    .B1(_0285_),
    .B2(_0279_),
    .ZN(_0356_));
 AND3_X1 _1279_ (.A1(_0326_),
    .A2(_0355_),
    .A3(_0356_),
    .ZN(_0357_));
 OAI22_X2 _1280_ (.A1(net44),
    .A2(_0347_),
    .B1(_0354_),
    .B2(_0357_),
    .ZN(_0358_));
 NOR3_X4 _1281_ (.A1(_0288_),
    .A2(net11),
    .A3(_0302_),
    .ZN(_0359_));
 AND3_X1 _1282_ (.A1(_0334_),
    .A2(_0327_),
    .A3(_0341_),
    .ZN(_0360_));
 XNOR2_X2 _1283_ (.A(_0339_),
    .B(_0360_),
    .ZN(_0361_));
 NAND4_X4 _1284_ (.A1(_0287_),
    .A2(_0359_),
    .A3(_0330_),
    .A4(_0361_),
    .ZN(_0362_));
 NAND2_X1 _1285_ (.A1(_0353_),
    .A2(_0352_),
    .ZN(_0363_));
 NAND2_X1 _1286_ (.A1(_0349_),
    .A2(_0351_),
    .ZN(_0364_));
 NAND2_X2 _1287_ (.A1(_0363_),
    .A2(_0364_),
    .ZN(_0365_));
 AOI21_X4 _1288_ (.A(_0358_),
    .B1(_0362_),
    .B2(_0365_),
    .ZN(_0366_));
 NAND2_X4 _1289_ (.A1(_0355_),
    .A2(_0356_),
    .ZN(_0367_));
 NAND2_X1 _1290_ (.A1(_0295_),
    .A2(_0327_),
    .ZN(_0368_));
 AND3_X1 _1291_ (.A1(_0335_),
    .A2(_0338_),
    .A3(_0290_),
    .ZN(_0369_));
 OAI21_X1 _1292_ (.A(_0369_),
    .B1(_0350_),
    .B2(_0279_),
    .ZN(_0370_));
 NAND3_X1 _1293_ (.A1(_0334_),
    .A2(_0339_),
    .A3(_0341_),
    .ZN(_0371_));
 AOI21_X2 _1294_ (.A(_0368_),
    .B1(_0370_),
    .B2(_0371_),
    .ZN(_0372_));
 OAI21_X4 _1295_ (.A(_0359_),
    .B1(_0372_),
    .B2(_0287_),
    .ZN(_0373_));
 XNOR2_X2 _1296_ (.A(_0367_),
    .B(_0373_),
    .ZN(_0374_));
 AND2_X1 _1297_ (.A1(_0315_),
    .A2(_0329_),
    .ZN(_0375_));
 OR2_X2 _1298_ (.A1(_0375_),
    .A2(_0328_),
    .ZN(_0376_));
 AOI221_X2 _1299_ (.A(_0272_),
    .B1(_0294_),
    .B2(_0290_),
    .C1(_0274_),
    .C2(_0273_),
    .ZN(_0377_));
 OAI211_X2 _1300_ (.A(_0266_),
    .B(_0377_),
    .C1(net24),
    .C2(_0268_),
    .ZN(_0378_));
 NAND2_X1 _1301_ (.A1(_0157_),
    .A2(_0172_),
    .ZN(_0379_));
 AOI221_X2 _1302_ (.A(_0231_),
    .B1(_0324_),
    .B2(_0379_),
    .C1(_0206_),
    .C2(_0314_),
    .ZN(_0380_));
 NOR2_X1 _1303_ (.A1(_0174_),
    .A2(net37),
    .ZN(_0381_));
 OR2_X1 _1304_ (.A1(_0160_),
    .A2(_0299_),
    .ZN(_0382_));
 NAND2_X1 _1305_ (.A1(_0314_),
    .A2(_0206_),
    .ZN(_0383_));
 AOI211_X2 _1306_ (.A(_0381_),
    .B(_0382_),
    .C1(_0383_),
    .C2(_0320_),
    .ZN(_0384_));
 OAI22_X4 _1307_ (.A1(net39),
    .A2(_0378_),
    .B1(_0380_),
    .B2(_0384_),
    .ZN(_0385_));
 NOR2_X1 _1308_ (.A1(_0376_),
    .A2(_0385_),
    .ZN(_0386_));
 INV_X2 _1309_ (.A(_0386_),
    .ZN(_0387_));
 XNOR2_X2 _1310_ (.A(_0369_),
    .B(_0360_),
    .ZN(_0388_));
 CLKBUF_X3 _1311_ (.A(_0819_),
    .Z(_0389_));
 NOR2_X2 _1312_ (.A1(_0288_),
    .A2(net9),
    .ZN(_0390_));
 NAND3_X4 _1313_ (.A1(_0389_),
    .A2(_0390_),
    .A3(_0301_),
    .ZN(_0391_));
 INV_X1 _1314_ (.A(_0298_),
    .ZN(_0392_));
 NAND3_X4 _1315_ (.A1(_0307_),
    .A2(_0377_),
    .A3(_0327_),
    .ZN(_0393_));
 NOR4_X4 _1316_ (.A1(_0279_),
    .A2(net64),
    .A3(_0280_),
    .A4(_0285_),
    .ZN(_0394_));
 NAND2_X1 _1317_ (.A1(_0298_),
    .A2(_0276_),
    .ZN(_0395_));
 OAI22_X4 _1318_ (.A1(_0392_),
    .A2(_0393_),
    .B1(_0394_),
    .B2(_0395_),
    .ZN(_0396_));
 AOI221_X2 _1319_ (.A(_0298_),
    .B1(_0307_),
    .B2(_0317_),
    .C1(_0276_),
    .C2(_0286_),
    .ZN(_0397_));
 OAI22_X4 _1320_ (.A1(_0347_),
    .A2(net46),
    .B1(_0396_),
    .B2(_0397_),
    .ZN(_0398_));
 OR4_X4 _1321_ (.A1(_0398_),
    .A2(_0388_),
    .A3(_0391_),
    .A4(_0387_),
    .ZN(_0399_));
 NOR2_X4 _1322_ (.A1(net70),
    .A2(_0374_),
    .ZN(_0400_));
 NOR2_X1 _1323_ (.A1(_0366_),
    .A2(net72),
    .ZN(_0841_));
 OR2_X2 _1324_ (.A1(_0391_),
    .A2(_0398_),
    .ZN(_0401_));
 NOR4_X1 _1325_ (.A1(_0288_),
    .A2(net74),
    .A3(_0302_),
    .A4(_0385_),
    .ZN(_0402_));
 NAND3_X1 _1326_ (.A1(_0295_),
    .A2(_0327_),
    .A3(_0330_),
    .ZN(_0403_));
 AOI21_X1 _1327_ (.A(_0403_),
    .B1(_0371_),
    .B2(_0370_),
    .ZN(_0404_));
 OAI21_X1 _1328_ (.A(_0402_),
    .B1(_0404_),
    .B2(_0287_),
    .ZN(_0405_));
 AOI21_X1 _1329_ (.A(_0279_),
    .B1(_0393_),
    .B2(net10),
    .ZN(_0406_));
 NAND2_X1 _1330_ (.A1(_0224_),
    .A2(_0231_),
    .ZN(_0407_));
 NOR4_X1 _1331_ (.A1(_0381_),
    .A2(_0407_),
    .A3(_0299_),
    .A4(_0300_),
    .ZN(_0408_));
 OAI21_X1 _1332_ (.A(_0408_),
    .B1(_0270_),
    .B2(_0217_),
    .ZN(_0409_));
 AOI21_X2 _1333_ (.A(_0406_),
    .B1(_0409_),
    .B2(_0376_),
    .ZN(_0410_));
 XOR2_X1 _1334_ (.A(_0405_),
    .B(_0410_),
    .Z(_0411_));
 INV_X1 _1335_ (.A(_0276_),
    .ZN(_0412_));
 OAI21_X2 _1336_ (.A(_0393_),
    .B1(_0412_),
    .B2(_0394_),
    .ZN(_0413_));
 NOR4_X2 _1337_ (.A1(net44),
    .A2(_0413_),
    .A3(_0376_),
    .A4(_0388_),
    .ZN(_0414_));
 NAND2_X1 _1338_ (.A1(_0359_),
    .A2(_0372_),
    .ZN(_0415_));
 OAI221_X1 _1339_ (.A(_0357_),
    .B1(_0414_),
    .B2(_0354_),
    .C1(_0415_),
    .C2(_0376_),
    .ZN(_0416_));
 OR3_X2 _1340_ (.A1(_0401_),
    .A2(_0411_),
    .A3(_0416_),
    .ZN(_0417_));
 NOR3_X2 _1341_ (.A1(net28),
    .A2(_0387_),
    .A3(_0373_),
    .ZN(_0418_));
 XNOR2_X2 _1342_ (.A(_0361_),
    .B(_0418_),
    .ZN(_0419_));
 AOI21_X4 _1343_ (.A(_0400_),
    .B1(_0417_),
    .B2(_0419_),
    .ZN(_0420_));
 OR2_X1 _1344_ (.A1(_0387_),
    .A2(_0373_),
    .ZN(_0421_));
 XOR2_X2 _1345_ (.A(_0367_),
    .B(_0421_),
    .Z(_0422_));
 XNOR2_X2 _1346_ (.A(_0366_),
    .B(_0389_),
    .ZN(_0423_));
 BUF_X2 _1347_ (.A(_0821_),
    .Z(_0424_));
 INV_X1 _1348_ (.A(_0424_),
    .ZN(_0425_));
 OR2_X1 _1349_ (.A1(_0288_),
    .A2(net9),
    .ZN(_0426_));
 NOR3_X4 _1350_ (.A1(_0425_),
    .A2(_0426_),
    .A3(net85),
    .ZN(_0427_));
 NOR3_X1 _1351_ (.A1(_0413_),
    .A2(net47),
    .A3(_0326_),
    .ZN(_0428_));
 OAI21_X1 _1352_ (.A(_0359_),
    .B1(_0404_),
    .B2(_0287_),
    .ZN(_0429_));
 AND2_X1 _1353_ (.A1(_0326_),
    .A2(_0429_),
    .ZN(_0430_));
 OAI221_X2 _1354_ (.A(_0389_),
    .B1(net44),
    .B2(_0347_),
    .C1(_0354_),
    .C2(_0357_),
    .ZN(_0431_));
 AOI21_X4 _1355_ (.A(_0431_),
    .B1(_0362_),
    .B2(_0365_),
    .ZN(_0432_));
 OAI21_X1 _1356_ (.A(_0224_),
    .B1(_0217_),
    .B2(_0270_),
    .ZN(_0433_));
 OAI221_X2 _1357_ (.A(_0298_),
    .B1(_0224_),
    .B2(_0217_),
    .C1(_0412_),
    .C2(_0394_),
    .ZN(_0434_));
 OAI211_X2 _1358_ (.A(_0433_),
    .B(_0434_),
    .C1(_0347_),
    .C2(net75),
    .ZN(_0435_));
 XOR2_X2 _1359_ (.A(_0301_),
    .B(_0435_),
    .Z(_0436_));
 OAI221_X2 _1360_ (.A(_0427_),
    .B1(_0428_),
    .B2(_0430_),
    .C1(_0432_),
    .C2(_0436_),
    .ZN(_0437_));
 XNOR2_X1 _1361_ (.A(_0405_),
    .B(_0410_),
    .ZN(_0438_));
 OR2_X1 _1362_ (.A1(_0354_),
    .A2(_0357_),
    .ZN(_0439_));
 OAI221_X2 _1363_ (.A(_0439_),
    .B1(_0414_),
    .B2(_0354_),
    .C1(_0415_),
    .C2(_0387_),
    .ZN(_0440_));
 OAI221_X2 _1364_ (.A(_0438_),
    .B1(_0374_),
    .B2(_0399_),
    .C1(_0401_),
    .C2(_0440_),
    .ZN(_0441_));
 NOR4_X4 _1365_ (.A1(_0437_),
    .A2(_0423_),
    .A3(_0400_),
    .A4(_0441_),
    .ZN(_0442_));
 AOI21_X4 _1366_ (.A(_0420_),
    .B1(_0422_),
    .B2(_0442_),
    .ZN(_0844_));
 NAND2_X1 _1367_ (.A1(_0420_),
    .A2(net20),
    .ZN(_0443_));
 XOR2_X2 _1368_ (.A(_0367_),
    .B(_0373_),
    .Z(_0444_));
 NOR4_X4 _1369_ (.A1(_0387_),
    .A2(_0388_),
    .A3(_0391_),
    .A4(net49),
    .ZN(_0445_));
 NAND2_X2 _1370_ (.A1(_0444_),
    .A2(_0445_),
    .ZN(_0446_));
 NOR2_X1 _1371_ (.A1(_0391_),
    .A2(net48),
    .ZN(_0447_));
 NAND3_X1 _1372_ (.A1(_0386_),
    .A2(_0366_),
    .A3(_0447_),
    .ZN(_0448_));
 NAND3_X1 _1373_ (.A1(_0446_),
    .A2(_0421_),
    .A3(_0448_),
    .ZN(_0449_));
 XOR2_X2 _1374_ (.A(_0367_),
    .B(_0449_),
    .Z(_0450_));
 OAI21_X2 _1375_ (.A(_0443_),
    .B1(_0450_),
    .B2(_0442_),
    .ZN(_0451_));
 INV_X1 _1376_ (.A(_0451_),
    .ZN(_0452_));
 NOR3_X1 _1377_ (.A1(net73),
    .A2(_0423_),
    .A3(_0437_),
    .ZN(_0453_));
 NOR4_X1 _1378_ (.A1(_0385_),
    .A2(_0440_),
    .A3(_0391_),
    .A4(net49),
    .ZN(_0454_));
 NOR2_X1 _1379_ (.A1(_0400_),
    .A2(_0454_),
    .ZN(_0455_));
 MUX2_X1 _1380_ (.A(_0330_),
    .B(_0411_),
    .S(_0455_),
    .Z(_0456_));
 NAND3_X1 _1381_ (.A1(_0420_),
    .A2(_0453_),
    .A3(_0456_),
    .ZN(_0457_));
 OR3_X1 _1382_ (.A1(net71),
    .A2(_0423_),
    .A3(_0437_),
    .ZN(_0458_));
 NAND2_X1 _1383_ (.A1(_0417_),
    .A2(_0419_),
    .ZN(_0459_));
 NAND2_X1 _1384_ (.A1(_0446_),
    .A2(_0459_),
    .ZN(_0460_));
 AOI21_X1 _1385_ (.A(_0458_),
    .B1(_0450_),
    .B2(_0460_),
    .ZN(_0461_));
 OAI21_X2 _1386_ (.A(_0457_),
    .B1(_0461_),
    .B2(_0456_),
    .ZN(_0462_));
 AOI21_X2 _1387_ (.A(net71),
    .B1(_0447_),
    .B2(_0366_),
    .ZN(_0463_));
 OAI21_X1 _1388_ (.A(_0463_),
    .B1(_0838_),
    .B2(_0303_),
    .ZN(_0464_));
 XNOR2_X1 _1389_ (.A(_0326_),
    .B(_0464_),
    .ZN(_0465_));
 NAND2_X1 _1390_ (.A1(_0389_),
    .A2(_0366_),
    .ZN(_0466_));
 NOR3_X1 _1391_ (.A1(_0426_),
    .A2(_0398_),
    .A3(_0466_),
    .ZN(_0467_));
 OAI21_X2 _1392_ (.A(_0463_),
    .B1(_0467_),
    .B2(_0436_),
    .ZN(_0468_));
 NOR2_X1 _1393_ (.A1(_0396_),
    .A2(net21),
    .ZN(_0469_));
 NOR2_X2 _1394_ (.A1(_0348_),
    .A2(_0469_),
    .ZN(_0470_));
 NAND2_X1 _1395_ (.A1(_0446_),
    .A2(_0466_),
    .ZN(_0471_));
 OAI21_X1 _1396_ (.A(_0424_),
    .B1(_0374_),
    .B2(_0399_),
    .ZN(_0472_));
 AOI211_X2 _1397_ (.A(_0423_),
    .B(_0472_),
    .C1(_0417_),
    .C2(_0419_),
    .ZN(_0473_));
 AOI211_X2 _1398_ (.A(_0471_),
    .B(_0473_),
    .C1(_0422_),
    .C2(net20),
    .ZN(_0474_));
 OR2_X2 _1399_ (.A1(_0470_),
    .A2(_0474_),
    .ZN(_0475_));
 NAND2_X1 _1400_ (.A1(_0470_),
    .A2(_0474_),
    .ZN(_0476_));
 AOI211_X2 _1401_ (.A(_0465_),
    .B(_0468_),
    .C1(_0475_),
    .C2(_0476_),
    .ZN(_0477_));
 AOI211_X4 _1402_ (.A(_0459_),
    .B(_0423_),
    .C1(_0422_),
    .C2(_0442_),
    .ZN(_0478_));
 AND2_X1 _1403_ (.A1(_0417_),
    .A2(_0419_),
    .ZN(_0479_));
 NAND2_X1 _1404_ (.A1(_0424_),
    .A2(_0423_),
    .ZN(_0480_));
 NAND2_X1 _1405_ (.A1(_0425_),
    .A2(_0446_),
    .ZN(_0481_));
 OAI22_X2 _1406_ (.A1(_0479_),
    .A2(_0480_),
    .B1(_0481_),
    .B2(_0423_),
    .ZN(_0482_));
 OAI21_X4 _1407_ (.A(_0851_),
    .B1(_0478_),
    .B2(_0482_),
    .ZN(_0483_));
 OAI21_X2 _1408_ (.A(_0298_),
    .B1(_0287_),
    .B2(net40),
    .ZN(_0484_));
 AOI21_X2 _1409_ (.A(_0390_),
    .B1(net40),
    .B2(_0287_),
    .ZN(_0485_));
 AOI21_X2 _1410_ (.A(net41),
    .B1(_0445_),
    .B2(_0444_),
    .ZN(_0486_));
 OAI21_X2 _1411_ (.A(_0392_),
    .B1(_0413_),
    .B2(_0486_),
    .ZN(_0487_));
 AOI21_X2 _1412_ (.A(_0426_),
    .B1(_0838_),
    .B2(_0486_),
    .ZN(_0488_));
 AOI22_X4 _1413_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_0487_),
    .B2(_0488_),
    .ZN(_0489_));
 NOR2_X1 _1414_ (.A1(net71),
    .A2(_0423_),
    .ZN(_0490_));
 NAND3_X1 _1415_ (.A1(_0424_),
    .A2(_0470_),
    .A3(_0490_),
    .ZN(_0491_));
 OAI21_X2 _1416_ (.A(_0489_),
    .B1(_0491_),
    .B2(net42),
    .ZN(_0492_));
 OR3_X4 _1417_ (.A1(_0390_),
    .A2(net42),
    .A3(_0491_),
    .ZN(_0493_));
 AOI21_X4 _1418_ (.A(_0483_),
    .B1(_0492_),
    .B2(_0493_),
    .ZN(_0494_));
 AND2_X1 _1419_ (.A1(_0824_),
    .A2(_0490_),
    .ZN(_0495_));
 XNOR2_X2 _1420_ (.A(_0844_),
    .B(_0424_),
    .ZN(_0850_));
 NAND2_X1 _1421_ (.A1(_0029_),
    .A2(_0032_),
    .ZN(_0496_));
 AND4_X1 _1422_ (.A1(_0489_),
    .A2(_0495_),
    .A3(net76),
    .A4(_0496_),
    .ZN(_0497_));
 OAI211_X2 _1423_ (.A(_0462_),
    .B(_0477_),
    .C1(_0497_),
    .C2(_0494_),
    .ZN(_0498_));
 AND2_X2 _1424_ (.A1(_0498_),
    .A2(_0452_),
    .ZN(_0847_));
 INV_X1 _1425_ (.A(_0852_),
    .ZN(_0499_));
 NOR2_X1 _1426_ (.A1(_0478_),
    .A2(_0482_),
    .ZN(_0500_));
 XOR2_X1 _1427_ (.A(_0851_),
    .B(_0500_),
    .Z(_0501_));
 NOR4_X1 _1428_ (.A1(_0824_),
    .A2(_0499_),
    .A3(_0452_),
    .A4(_0501_),
    .ZN(_0502_));
 NAND2_X1 _1429_ (.A1(_0495_),
    .A2(net76),
    .ZN(_0503_));
 NOR2_X1 _1430_ (.A1(_0451_),
    .A2(_0503_),
    .ZN(_0504_));
 AOI21_X1 _1431_ (.A(_0502_),
    .B1(_0504_),
    .B2(_0498_),
    .ZN(_0505_));
 INV_X1 _1432_ (.A(_0023_),
    .ZN(_0506_));
 NOR3_X2 _1433_ (.A1(_0026_),
    .A2(net4),
    .A3(net3),
    .ZN(_0507_));
 NAND3_X2 _1434_ (.A1(_0506_),
    .A2(_0858_),
    .A3(_0507_),
    .ZN(_0508_));
 NOR3_X1 _1435_ (.A1(net5),
    .A2(net6),
    .A3(_0508_),
    .ZN(_0509_));
 NOR2_X1 _1436_ (.A1(_0826_),
    .A2(_0509_),
    .ZN(_0510_));
 INV_X1 _1437_ (.A(_0833_),
    .ZN(_0511_));
 INV_X1 _1438_ (.A(_0839_),
    .ZN(_0512_));
 AOI21_X2 _1439_ (.A(_0845_),
    .B1(_0848_),
    .B2(_0846_),
    .ZN(_0513_));
 INV_X2 _1440_ (.A(_0513_),
    .ZN(_0514_));
 AOI21_X4 _1441_ (.A(_0842_),
    .B1(_0843_),
    .B2(_0514_),
    .ZN(_0515_));
 INV_X1 _1442_ (.A(_0840_),
    .ZN(_0516_));
 OAI21_X4 _1443_ (.A(_0512_),
    .B1(_0515_),
    .B2(_0516_),
    .ZN(_0517_));
 AOI21_X4 _1444_ (.A(_0836_),
    .B1(_0517_),
    .B2(_0837_),
    .ZN(_0518_));
 INV_X1 _1445_ (.A(_0834_),
    .ZN(_0519_));
 OAI21_X4 _1446_ (.A(_0511_),
    .B1(_0519_),
    .B2(_0518_),
    .ZN(_0520_));
 AOI21_X4 _1447_ (.A(_0830_),
    .B1(_0520_),
    .B2(_0831_),
    .ZN(_0521_));
 INV_X1 _1448_ (.A(_0827_),
    .ZN(_0522_));
 OAI21_X4 _1449_ (.A(_0510_),
    .B1(_0521_),
    .B2(_0522_),
    .ZN(_0523_));
 OR2_X4 _1450_ (.A1(_0523_),
    .A2(\counter[0] ),
    .ZN(_0524_));
 OR3_X4 _1451_ (.A1(_0465_),
    .A2(_0524_),
    .A3(_0496_),
    .ZN(_0525_));
 AOI21_X4 _1452_ (.A(_0525_),
    .B1(_0492_),
    .B2(_0493_),
    .ZN(_0526_));
 NOR3_X1 _1453_ (.A1(_0452_),
    .A2(_0468_),
    .A3(_0503_),
    .ZN(_0527_));
 NAND4_X1 _1454_ (.A1(_0451_),
    .A2(_0489_),
    .A3(_0495_),
    .A4(net76),
    .ZN(_0528_));
 AOI22_X1 _1455_ (.A1(_0475_),
    .A2(_0476_),
    .B1(_0468_),
    .B2(_0528_),
    .ZN(_0529_));
 OAI21_X2 _1456_ (.A(_0526_),
    .B1(_0527_),
    .B2(_0529_),
    .ZN(_0530_));
 NAND4_X1 _1457_ (.A1(_0837_),
    .A2(_0843_),
    .A3(_0846_),
    .A4(_0849_),
    .ZN(_0531_));
 NAND4_X1 _1458_ (.A1(_0827_),
    .A2(_0840_),
    .A3(_0831_),
    .A4(_0834_),
    .ZN(_0532_));
 NOR2_X1 _1459_ (.A1(_0531_),
    .A2(_0532_),
    .ZN(_0533_));
 NAND3_X1 _1460_ (.A1(_0425_),
    .A2(_0489_),
    .A3(_0495_),
    .ZN(_0534_));
 NOR2_X1 _1461_ (.A1(_0844_),
    .A2(_0534_),
    .ZN(_0535_));
 AND4_X1 _1462_ (.A1(_0424_),
    .A2(net42),
    .A3(_0489_),
    .A4(_0495_),
    .ZN(_0536_));
 OAI221_X2 _1463_ (.A(net65),
    .B1(_0535_),
    .B2(_0536_),
    .C1(net38),
    .C2(_0451_),
    .ZN(_0537_));
 NOR2_X1 _1464_ (.A1(_0452_),
    .A2(_0462_),
    .ZN(_0538_));
 AND4_X1 _1465_ (.A1(_0477_),
    .A2(_0489_),
    .A3(_0495_),
    .A4(net77),
    .ZN(_0539_));
 AOI22_X2 _1466_ (.A1(_0462_),
    .A2(_0537_),
    .B1(_0538_),
    .B2(_0539_),
    .ZN(_0540_));
 OAI222_X2 _1467_ (.A1(_0530_),
    .A2(_0505_),
    .B1(_0533_),
    .B2(_0523_),
    .C1(_0540_),
    .C2(_0524_),
    .ZN(_0000_));
 NOR3_X1 _1468_ (.A1(_0030_),
    .A2(_0031_),
    .A3(_0032_),
    .ZN(_0541_));
 XNOR2_X1 _1469_ (.A(_0028_),
    .B(_0541_),
    .ZN(_0862_));
 XNOR2_X1 _1470_ (.A(_0030_),
    .B(_0858_),
    .ZN(_0865_));
 INV_X1 _1471_ (.A(_0031_),
    .ZN(_0857_));
 INV_X1 _1472_ (.A(_0032_),
    .ZN(_0854_));
 NAND3_X1 _1473_ (.A1(_0857_),
    .A2(_0854_),
    .A3(_0507_),
    .ZN(_0542_));
 NOR3_X1 _1474_ (.A1(net2),
    .A2(_0023_),
    .A3(_0542_),
    .ZN(_0543_));
 XNOR2_X1 _1475_ (.A(net6),
    .B(_0543_),
    .ZN(_0868_));
 XOR2_X2 _1476_ (.A(net2),
    .B(_0508_),
    .Z(_0871_));
 XNOR2_X1 _1477_ (.A(_0506_),
    .B(_0542_),
    .ZN(_0874_));
 INV_X1 _1478_ (.A(_0858_),
    .ZN(_0544_));
 NOR3_X1 _1479_ (.A1(_0028_),
    .A2(net3),
    .A3(_0544_),
    .ZN(_0545_));
 XNOR2_X1 _1480_ (.A(_0026_),
    .B(_0545_),
    .ZN(_0877_));
 INV_X1 _1481_ (.A(_0870_),
    .ZN(_0546_));
 INV_X1 _1482_ (.A(_0872_),
    .ZN(_0547_));
 INV_X1 _1483_ (.A(_0876_),
    .ZN(_0548_));
 INV_X1 _1484_ (.A(_0864_),
    .ZN(_0549_));
 INV_X1 _1485_ (.A(_0866_),
    .ZN(_0550_));
 INV_X1 _1486_ (.A(_0861_),
    .ZN(_0551_));
 INV_X1 _1487_ (.A(_0856_),
    .ZN(_0552_));
 AOI21_X1 _1488_ (.A(_0551_),
    .B1(_0855_),
    .B2(_0552_),
    .ZN(_0553_));
 OAI21_X1 _1489_ (.A(_0867_),
    .B1(_0860_),
    .B2(_0553_),
    .ZN(_0554_));
 AOI21_X1 _1490_ (.A(_0549_),
    .B1(_0550_),
    .B2(_0554_),
    .ZN(_0555_));
 OAI21_X1 _1491_ (.A(_0879_),
    .B1(_0863_),
    .B2(_0555_),
    .ZN(_0556_));
 INV_X1 _1492_ (.A(_0878_),
    .ZN(_0557_));
 AOI21_X1 _1493_ (.A(_0548_),
    .B1(_0556_),
    .B2(_0557_),
    .ZN(_0558_));
 OAI21_X1 _1494_ (.A(_0873_),
    .B1(_0875_),
    .B2(_0558_),
    .ZN(_0559_));
 AOI21_X1 _1495_ (.A(_0546_),
    .B1(_0547_),
    .B2(_0559_),
    .ZN(_0560_));
 INV_X1 _1496_ (.A(_0015_),
    .ZN(_0561_));
 OAI33_X1 _1497_ (.A1(net5),
    .A2(net6),
    .A3(_0508_),
    .B1(_0560_),
    .B2(_0561_),
    .B3(_0869_),
    .ZN(_0562_));
 INV_X2 _1498_ (.A(_0562_),
    .ZN(_0563_));
 NOR2_X1 _1499_ (.A1(\counter[0] ),
    .A2(_0563_),
    .ZN(_0001_));
 AND2_X1 _1500_ (.A1(_0881_),
    .A2(_0562_),
    .ZN(_0002_));
 XOR2_X1 _1501_ (.A(_0880_),
    .B(_0013_),
    .Z(_0564_));
 NOR2_X1 _1502_ (.A1(_0563_),
    .A2(_0564_),
    .ZN(_0003_));
 NAND3_X2 _1503_ (.A1(\counter[0] ),
    .A2(\counter[2] ),
    .A3(\counter[1] ),
    .ZN(_0565_));
 XNOR2_X1 _1504_ (.A(_0012_),
    .B(_0565_),
    .ZN(_0566_));
 NOR2_X1 _1505_ (.A1(_0563_),
    .A2(_0566_),
    .ZN(_0004_));
 AND2_X1 _1506_ (.A1(_0880_),
    .A2(\counter[2] ),
    .ZN(_0567_));
 NAND2_X1 _1507_ (.A1(\counter[3] ),
    .A2(_0567_),
    .ZN(_0568_));
 XNOR2_X1 _1508_ (.A(_0014_),
    .B(_0568_),
    .ZN(_0569_));
 NOR2_X1 _1509_ (.A1(_0563_),
    .A2(_0569_),
    .ZN(_0005_));
 INV_X1 _1510_ (.A(_0565_),
    .ZN(_0570_));
 NAND3_X1 _1511_ (.A1(\counter[3] ),
    .A2(\counter[4] ),
    .A3(_0570_),
    .ZN(_0571_));
 XNOR2_X1 _1512_ (.A(_0011_),
    .B(_0571_),
    .ZN(_0572_));
 NOR2_X1 _1513_ (.A1(_0563_),
    .A2(_0572_),
    .ZN(_0006_));
 NAND4_X1 _1514_ (.A1(\counter[3] ),
    .A2(\counter[4] ),
    .A3(\counter[5] ),
    .A4(_0567_),
    .ZN(_0573_));
 XNOR2_X1 _1515_ (.A(_0010_),
    .B(_0573_),
    .ZN(_0574_));
 NOR2_X1 _1516_ (.A1(_0563_),
    .A2(_0574_),
    .ZN(_0007_));
 NAND4_X1 _1517_ (.A1(\counter[3] ),
    .A2(\counter[4] ),
    .A3(\counter[5] ),
    .A4(\counter[6] ),
    .ZN(_0575_));
 NOR2_X1 _1518_ (.A1(_0565_),
    .A2(_0575_),
    .ZN(_0576_));
 XOR2_X1 _1519_ (.A(_0016_),
    .B(_0576_),
    .Z(_0577_));
 NOR2_X1 _1520_ (.A1(_0563_),
    .A2(_0577_),
    .ZN(_0008_));
 NAND2_X1 _1521_ (.A1(\counter[7] ),
    .A2(_0567_),
    .ZN(_0578_));
 NOR2_X1 _1522_ (.A1(_0575_),
    .A2(_0578_),
    .ZN(_0579_));
 XNOR2_X1 _1523_ (.A(_0561_),
    .B(_0579_),
    .ZN(_0580_));
 NOR2_X1 _1524_ (.A1(_0563_),
    .A2(_0580_),
    .ZN(_0009_));
 INV_X1 _1525_ (.A(_0767_),
    .ZN(_0632_));
 INV_X1 _1526_ (.A(_0622_),
    .ZN(_0637_));
 INV_X1 _1527_ (.A(_0774_),
    .ZN(_0727_));
 NAND2_X1 _1528_ (.A1(_0027_),
    .A2(_0030_),
    .ZN(_0731_));
 NAND2_X1 _1529_ (.A1(_0028_),
    .A2(_0029_),
    .ZN(_0735_));
 INV_X1 _1530_ (.A(_0594_),
    .ZN(_0589_));
 NAND2_X1 _1531_ (.A1(_0019_),
    .A2(_0028_),
    .ZN(_0633_));
 INV_X1 _1532_ (.A(_0684_),
    .ZN(_0686_));
 NAND2_X1 _1533_ (.A1(_0025_),
    .A2(_0031_),
    .ZN(_0732_));
 INV_X1 _1534_ (.A(_0781_),
    .ZN(_0736_));
 INV_X1 _1535_ (.A(_0586_),
    .ZN(_0590_));
 INV_X1 _1536_ (.A(_0614_),
    .ZN(_0617_));
 NAND2_X1 _1537_ (.A1(_0017_),
    .A2(_0030_),
    .ZN(_0634_));
 INV_X1 _1538_ (.A(_0660_),
    .ZN(_0663_));
 INV_X1 _1539_ (.A(_0615_),
    .ZN(_0621_));
 INV_X1 _1540_ (.A(_0627_),
    .ZN(_0642_));
 INV_X1 _1541_ (.A(_0631_),
    .ZN(_0645_));
 INV_X1 _1542_ (.A(_0648_),
    .ZN(_0666_));
 INV_X1 _1543_ (.A(_0652_),
    .ZN(_0670_));
 INV_X2 _1544_ (.A(_0672_),
    .ZN(_0690_));
 INV_X1 _1545_ (.A(_0676_),
    .ZN(_0694_));
 INV_X2 _1546_ (.A(_0693_),
    .ZN(_0708_));
 INV_X1 _1547_ (.A(_0696_),
    .ZN(_0713_));
 INV_X1 _1548_ (.A(_0700_),
    .ZN(_0716_));
 INV_X2 _1549_ (.A(_0710_),
    .ZN(_0814_));
 INV_X1 _1550_ (.A(_0714_),
    .ZN(_0778_));
 INV_X1 _1551_ (.A(_0717_),
    .ZN(_0724_));
 INV_X1 _1552_ (.A(_0726_),
    .ZN(_0786_));
 INV_X1 _1553_ (.A(_0626_),
    .ZN(_0620_));
 INV_X1 _1554_ (.A(_0641_),
    .ZN(_0638_));
 INV_X1 _1555_ (.A(_0668_),
    .ZN(_0662_));
 INV_X1 _1556_ (.A(_0692_),
    .ZN(_0687_));
 AND2_X1 _1557_ (.A1(net6),
    .A2(_0024_),
    .ZN(_0607_));
 INV_X1 _1558_ (.A(_0592_),
    .ZN(_0758_));
 AND2_X1 _1559_ (.A1(_0023_),
    .A2(_0024_),
    .ZN(_0628_));
 AND2_X1 _1560_ (.A1(_0024_),
    .A2(_0026_),
    .ZN(_0649_));
 AND2_X1 _1561_ (.A1(_0024_),
    .A2(_0028_),
    .ZN(_0673_));
 AND2_X1 _1562_ (.A1(_0024_),
    .A2(_0030_),
    .ZN(_0697_));
 INV_X1 _1563_ (.A(_0729_),
    .ZN(_0723_));
 INV_X1 _1564_ (.A(_0737_),
    .ZN(_0787_));
 INV_X1 _1565_ (.A(_0619_),
    .ZN(_0802_));
 INV_X1 _1566_ (.A(_0640_),
    .ZN(_0806_));
 INV_X1 _1567_ (.A(_0665_),
    .ZN(_0810_));
 INV_X1 _1568_ (.A(_0591_),
    .ZN(_0750_));
 INV_X1 _1569_ (.A(_0618_),
    .ZN(_0768_));
 AND2_X1 _1570_ (.A1(_0024_),
    .A2(_0031_),
    .ZN(_0720_));
 INV_X2 _1571_ (.A(_0689_),
    .ZN(_0775_));
 INV_X1 _1572_ (.A(_0730_),
    .ZN(_0788_));
 INV_X1 _1573_ (.A(_0738_),
    .ZN(_0798_));
 INV_X1 _1574_ (.A(_0639_),
    .ZN(_0803_));
 INV_X1 _1575_ (.A(_0664_),
    .ZN(_0807_));
 INV_X1 _1576_ (.A(_0688_),
    .ZN(_0811_));
 INV_X1 _1577_ (.A(_0593_),
    .ZN(_0588_));
 FA_X1 _1578_ (.A(_0583_),
    .B(_0584_),
    .CI(_0585_),
    .CO(_0586_),
    .S(_0587_));
 FA_X1 _1579_ (.A(_0588_),
    .B(_0589_),
    .CI(_0590_),
    .CO(_0591_),
    .S(_0592_));
 FA_X1 _1580_ (.A(_0595_),
    .B(_0596_),
    .CI(_0597_),
    .CO(_0598_),
    .S(_0599_));
 FA_X1 _1581_ (.A(_0600_),
    .B(_0601_),
    .CI(_0598_),
    .CO(_0602_),
    .S(_0603_));
 FA_X1 _1582_ (.A(_0604_),
    .B(_0605_),
    .CI(_0599_),
    .CO(_0601_),
    .S(_0606_));
 FA_X1 _1583_ (.A(_0607_),
    .B(_0608_),
    .CI(_0609_),
    .CO(_0605_),
    .S(_0610_));
 FA_X1 _1584_ (.A(_0611_),
    .B(_0612_),
    .CI(_0613_),
    .CO(_0614_),
    .S(_0615_));
 FA_X1 _1585_ (.A(_0606_),
    .B(_0616_),
    .CI(_0617_),
    .CO(_0618_),
    .S(_0619_));
 FA_X1 _1586_ (.A(_0610_),
    .B(_0620_),
    .CI(_0621_),
    .CO(_0616_),
    .S(_0622_));
 FA_X1 _1587_ (.A(_0623_),
    .B(_0624_),
    .CI(_0625_),
    .CO(_0626_),
    .S(_0627_));
 FA_X1 _1588_ (.A(_0628_),
    .B(_0629_),
    .CI(_0630_),
    .CO(_0624_),
    .S(_0631_));
 FA_X1 _1589_ (.A(_0632_),
    .B(_0633_),
    .CI(_0634_),
    .CO(_0635_),
    .S(_0636_));
 FA_X1 _1590_ (.A(_0637_),
    .B(_0638_),
    .CI(_0635_),
    .CO(_0639_),
    .S(_0640_));
 FA_X1 _1591_ (.A(_0642_),
    .B(_0643_),
    .CI(_0636_),
    .CO(_0641_),
    .S(_0644_));
 FA_X1 _1592_ (.A(_0645_),
    .B(_0646_),
    .CI(_0647_),
    .CO(_0643_),
    .S(_0648_));
 FA_X1 _1593_ (.A(_0649_),
    .B(_0651_),
    .CI(_0650_),
    .CO(_0646_),
    .S(_0652_));
 FA_X1 _1594_ (.A(_0655_),
    .B(_0654_),
    .CI(_0653_),
    .CO(_0656_),
    .S(_0657_));
 FA_X1 _1595_ (.A(_0656_),
    .B(_0658_),
    .CI(_0659_),
    .CO(_0660_),
    .S(_0661_));
 FA_X1 _1596_ (.A(_0644_),
    .B(_0662_),
    .CI(_0663_),
    .CO(_0664_),
    .S(_0665_));
 FA_X1 _1597_ (.A(_0661_),
    .B(_0667_),
    .CI(_0666_),
    .CO(_0668_),
    .S(_0669_));
 FA_X1 _1598_ (.A(_0657_),
    .B(_0671_),
    .CI(_0670_),
    .CO(_0667_),
    .S(_0672_));
 FA_X1 _1599_ (.A(_0673_),
    .B(_0674_),
    .CI(_0675_),
    .CO(_0671_),
    .S(_0676_));
 FA_X1 _1600_ (.A(_0677_),
    .B(_0678_),
    .CI(_0679_),
    .CO(_0680_),
    .S(_0681_));
 FA_X1 _1601_ (.A(_0680_),
    .B(_0682_),
    .CI(_0683_),
    .CO(_0684_),
    .S(_0685_));
 FA_X1 _1602_ (.A(_0687_),
    .B(_0686_),
    .CI(_0669_),
    .CO(_0688_),
    .S(_0689_));
 FA_X1 _1603_ (.A(_0685_),
    .B(_0691_),
    .CI(_0690_),
    .CO(_0692_),
    .S(_0693_));
 FA_X1 _1604_ (.A(_0694_),
    .B(_0695_),
    .CI(_0681_),
    .CO(_0691_),
    .S(_0696_));
 FA_X1 _1605_ (.A(_0697_),
    .B(_0698_),
    .CI(_0699_),
    .CO(_0695_),
    .S(_0700_));
 FA_X1 _1606_ (.A(_0701_),
    .B(_0702_),
    .CI(_0703_),
    .CO(_0704_),
    .S(_0705_));
 FA_X1 _1607_ (.A(_0706_),
    .B(_0707_),
    .CI(_0708_),
    .CO(_0709_),
    .S(_0710_));
 FA_X1 _1608_ (.A(_0711_),
    .B(_0712_),
    .CI(_0713_),
    .CO(_0707_),
    .S(_0714_));
 FA_X1 _1609_ (.A(_0705_),
    .B(_0715_),
    .CI(_0716_),
    .CO(_0712_),
    .S(_0717_));
 FA_X1 _1610_ (.A(_0718_),
    .B(_0719_),
    .CI(_0720_),
    .CO(_0715_),
    .S(_0721_));
 FA_X1 _1611_ (.A(_0722_),
    .B(_0723_),
    .CI(_0724_),
    .CO(_0725_),
    .S(_0726_));
 FA_X1 _1612_ (.A(_0727_),
    .B(_0728_),
    .CI(_0721_),
    .CO(_0729_),
    .S(_0730_));
 FA_X1 _1613_ (.A(_0731_),
    .B(_0732_),
    .CI(_0733_),
    .CO(_0728_),
    .S(_0734_));
 FA_X1 _1614_ (.A(_0735_),
    .B(_0736_),
    .CI(_0734_),
    .CO(_0737_),
    .S(_0738_));
 FA_X1 _1615_ (.A(_0739_),
    .B(_0740_),
    .CI(_0741_),
    .CO(_0742_),
    .S(_0743_));
 HA_X1 _1616_ (.A(_0744_),
    .B(_0745_),
    .CO(_0746_),
    .S(_0747_));
 HA_X1 _1617_ (.A(_0748_),
    .B(_0749_),
    .CO(_0744_),
    .S(_0593_));
 HA_X1 _1618_ (.A(_0747_),
    .B(_0750_),
    .CO(_0751_),
    .S(_0752_));
 HA_X1 _1619_ (.A(_0587_),
    .B(_0753_),
    .CO(_0594_),
    .S(_0600_));
 HA_X1 _1620_ (.A(_0754_),
    .B(_0755_),
    .CO(_0583_),
    .S(_0604_));
 HA_X1 _1621_ (.A(_0756_),
    .B(_0757_),
    .CO(_0595_),
    .S(_0609_));
 HA_X1 _1622_ (.A(_0758_),
    .B(_0602_),
    .CO(_0759_),
    .S(_0760_));
 HA_X1 _1623_ (.A(_0761_),
    .B(_0762_),
    .CO(_0608_),
    .S(_0623_));
 HA_X1 _1624_ (.A(_0763_),
    .B(_0764_),
    .CO(_0611_),
    .S(_0625_));
 HA_X1 _1625_ (.A(_0765_),
    .B(_0766_),
    .CO(_0767_),
    .S(_0647_));
 HA_X1 _1626_ (.A(_0603_),
    .B(_0768_),
    .CO(_0769_),
    .S(_0770_));
 HA_X1 _1627_ (.A(_0771_),
    .B(_0704_),
    .CO(_0706_),
    .S(_0711_));
 HA_X1 _1628_ (.A(_0772_),
    .B(_0773_),
    .CO(_0722_),
    .S(_0774_));
 HA_X1 _1629_ (.A(_0775_),
    .B(_0709_),
    .CO(_0776_),
    .S(_0777_));
 HA_X1 _1630_ (.A(_0725_),
    .B(_0778_),
    .CO(_0779_),
    .S(_0780_));
 HA_X1 _1631_ (.A(_0782_),
    .B(_0780_),
    .CO(_0783_),
    .S(_0784_));
 HA_X1 _1632_ (.A(_0785_),
    .B(_0786_),
    .CO(_0782_),
    .S(_0740_));
 HA_X1 _1633_ (.A(_0787_),
    .B(_0788_),
    .CO(_0785_),
    .S(_0789_));
 HA_X1 _1634_ (.A(_0790_),
    .B(_0791_),
    .CO(_0781_),
    .S(_0792_));
 HA_X1 _1635_ (.A(_0739_),
    .B(_0740_),
    .CO(_0793_),
    .S(_0794_));
 HA_X1 _1636_ (.A(_0795_),
    .B(_0789_),
    .CO(_0739_),
    .S(_0796_));
 HA_X1 _1637_ (.A(_0797_),
    .B(_0798_),
    .CO(_0795_),
    .S(_0799_));
 HA_X1 _1638_ (.A(_0792_),
    .B(_0800_),
    .CO(_0797_),
    .S(_0801_));
 HA_X1 _1639_ (.A(_0802_),
    .B(_0803_),
    .CO(_0804_),
    .S(_0805_));
 HA_X1 _1640_ (.A(_0806_),
    .B(_0807_),
    .CO(_0808_),
    .S(_0809_));
 HA_X1 _1641_ (.A(_0810_),
    .B(_0811_),
    .CO(_0812_),
    .S(_0813_));
 HA_X1 _1642_ (.A(_0779_),
    .B(_0814_),
    .CO(_0815_),
    .S(_0816_));
 HA_X1 _1643_ (.A(_0817_),
    .B(_0799_),
    .CO(_0818_),
    .S(_0819_));
 HA_X1 _1644_ (.A(_0820_),
    .B(_0801_),
    .CO(_0817_),
    .S(_0821_));
 HA_X1 _1645_ (.A(_0822_),
    .B(_0823_),
    .CO(_0820_),
    .S(_0824_));
 HA_X1 _1646_ (.A(\counter[8] ),
    .B(_0825_),
    .CO(_0826_),
    .S(_0827_));
 HA_X1 _1647_ (.A(_0796_),
    .B(_0818_),
    .CO(_0741_),
    .S(_0828_));
 HA_X1 _1648_ (.A(\counter[7] ),
    .B(_0829_),
    .CO(_0830_),
    .S(_0831_));
 HA_X1 _1649_ (.A(\counter[6] ),
    .B(_0832_),
    .CO(_0833_),
    .S(_0834_));
 HA_X1 _1650_ (.A(\counter[5] ),
    .B(_0835_),
    .CO(_0836_),
    .S(_0837_));
 HA_X1 _1651_ (.A(\counter[4] ),
    .B(_0838_),
    .CO(_0839_),
    .S(_0840_));
 HA_X1 _1652_ (.A(\counter[3] ),
    .B(_0841_),
    .CO(_0842_),
    .S(_0843_));
 HA_X1 _1653_ (.A(\counter[2] ),
    .B(net43),
    .CO(_0845_),
    .S(_0846_));
 HA_X1 _1654_ (.A(\counter[1] ),
    .B(_0847_),
    .CO(_0848_),
    .S(_0849_));
 HA_X1 _1655_ (.A(_0824_),
    .B(_0850_),
    .CO(_0851_),
    .S(_0852_));
 HA_X1 _1656_ (.A(_0853_),
    .B(_0854_),
    .CO(_0855_),
    .S(_0856_));
 HA_X1 _1657_ (.A(_0854_),
    .B(_0857_),
    .CO(_0858_),
    .S(_0859_));
 HA_X1 _1658_ (.A(\counter[1] ),
    .B(_0859_),
    .CO(_0860_),
    .S(_0861_));
 HA_X1 _1659_ (.A(\counter[3] ),
    .B(_0862_),
    .CO(_0863_),
    .S(_0864_));
 HA_X1 _1660_ (.A(\counter[2] ),
    .B(_0865_),
    .CO(_0866_),
    .S(_0867_));
 HA_X1 _1661_ (.A(\counter[7] ),
    .B(_0868_),
    .CO(_0869_),
    .S(_0870_));
 HA_X1 _1662_ (.A(\counter[6] ),
    .B(_0871_),
    .CO(_0872_),
    .S(_0873_));
 HA_X1 _1663_ (.A(\counter[5] ),
    .B(_0874_),
    .CO(_0875_),
    .S(_0876_));
 HA_X1 _1664_ (.A(\counter[4] ),
    .B(_0877_),
    .CO(_0878_),
    .S(_0879_));
 HA_X1 _1665_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_0880_),
    .S(_0881_));
 DFFR_X2 \clk_out$_DFF_PN0_  (.D(_0000_),
    .RN(net7),
    .CK(clknet_1_1__leaf_clk_in),
    .Q(net8),
    .QN(_0581_));
 DFFR_X2 \counter[0]$_DFF_PN0_  (.D(_0001_),
    .RN(net7),
    .CK(clknet_1_1__leaf_clk_in),
    .Q(\counter[0] ),
    .QN(_0853_));
 DFFR_X2 \counter[1]$_DFF_PN0_  (.D(_0002_),
    .RN(net7),
    .CK(clknet_1_1__leaf_clk_in),
    .Q(\counter[1] ),
    .QN(_0582_));
 DFFR_X2 \counter[2]$_DFF_PN0_  (.D(_0003_),
    .RN(net7),
    .CK(clknet_1_1__leaf_clk_in),
    .Q(\counter[2] ),
    .QN(_0013_));
 DFFR_X2 \counter[3]$_DFF_PN0_  (.D(_0004_),
    .RN(net7),
    .CK(clknet_1_1__leaf_clk_in),
    .Q(\counter[3] ),
    .QN(_0012_));
 DFFR_X2 \counter[4]$_DFF_PN0_  (.D(_0005_),
    .RN(net7),
    .CK(clknet_1_0__leaf_clk_in),
    .Q(\counter[4] ),
    .QN(_0014_));
 DFFR_X2 \counter[5]$_DFF_PN0_  (.D(_0006_),
    .RN(net7),
    .CK(clknet_1_0__leaf_clk_in),
    .Q(\counter[5] ),
    .QN(_0011_));
 DFFR_X2 \counter[6]$_DFF_PN0_  (.D(_0007_),
    .RN(net7),
    .CK(clknet_1_0__leaf_clk_in),
    .Q(\counter[6] ),
    .QN(_0010_));
 DFFR_X2 \counter[7]$_DFF_PN0_  (.D(_0008_),
    .RN(net7),
    .CK(clknet_1_0__leaf_clk_in),
    .Q(\counter[7] ),
    .QN(_0016_));
 DFFR_X1 \counter[8]$_DFF_PN0_  (.D(_0009_),
    .RN(net7),
    .CK(clknet_1_0__leaf_clk_in),
    .Q(\counter[8] ),
    .QN(_0015_));
 BUF_X2 clone1 (.A(net23),
    .Z(net1));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Right_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Right_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Right_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Right_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Right_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Left_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Left_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Left_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Left_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Left_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Left_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Left_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Left_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Left_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Left_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Left_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Left_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Left_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Left_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Left_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Left_659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_1002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_1005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_1008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_1011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_1014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_1017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_1020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_1023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_1026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_1029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_1032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_1035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_1038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_1041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_1044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_1047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_1050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_1053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_1056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_1059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_1062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_1065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_1068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_1071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_1074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_1077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_1080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_1083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_1092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_1095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_1098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_1101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_1104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_1107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_1110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_1113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_1116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_1119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_1122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_1125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_1128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_1131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_1134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_1137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_1140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_1143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_1146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_1149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_1152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1157 ();
 BUF_X1 input1 (.A(div_ratio[2]),
    .Z(net3));
 BUF_X1 input2 (.A(div_ratio[3]),
    .Z(net4));
 BUF_X4 input3 (.A(div_ratio[6]),
    .Z(net5));
 BUF_X2 input4 (.A(div_ratio[7]),
    .Z(net6));
 BUF_X4 input5 (.A(net81),
    .Z(net7));
 BUF_X1 output6 (.A(net8),
    .Z(clk_out));
 BUF_X4 max_cap7 (.A(net11),
    .Z(net9));
 CLKBUF_X2 wire8 (.A(_0284_),
    .Z(net10));
 CLKBUF_X3 clkbuf_0_clk_in (.A(clk_in),
    .Z(clknet_0_clk_in));
 CLKBUF_X3 clkbuf_1_0__f_clk_in (.A(clknet_0_clk_in),
    .Z(clknet_1_0__leaf_clk_in));
 CLKBUF_X3 clkbuf_1_1__f_clk_in (.A(clknet_0_clk_in),
    .Z(clknet_1_1__leaf_clk_in));
 CLKBUF_X1 clkload0 (.A(clknet_1_1__leaf_clk_in));
 BUF_X2 rebuffer1 (.A(_0297_),
    .Z(net11));
 BUF_X8 rebuffer2 (.A(net52),
    .Z(net12));
 BUF_X1 rebuffer3 (.A(net12),
    .Z(net13));
 BUF_X4 rebuffer4 (.A(_0138_),
    .Z(net14));
 BUF_X1 rebuffer5 (.A(net14),
    .Z(net15));
 BUF_X2 rebuffer6 (.A(net14),
    .Z(net16));
 BUF_X1 rebuffer7 (.A(net16),
    .Z(net17));
 BUF_X1 rebuffer8 (.A(net17),
    .Z(net18));
 BUF_X1 rebuffer9 (.A(net14),
    .Z(net19));
 BUF_X2 rebuffer10 (.A(_0442_),
    .Z(net20));
 BUF_X1 rebuffer11 (.A(net53),
    .Z(net21));
 BUF_X1 rebuffer12 (.A(_0190_),
    .Z(net22));
 BUF_X2 rebuffer13 (.A(_0129_),
    .Z(net23));
 BUF_X1 rebuffer14 (.A(net32),
    .Z(net24));
 BUF_X2 rebuffer15 (.A(net32),
    .Z(net25));
 BUF_X1 rebuffer16 (.A(_0241_),
    .Z(net26));
 BUF_X1 rebuffer17 (.A(_0269_),
    .Z(net27));
 BUF_X1 rebuffer18 (.A(_0269_),
    .Z(net28));
 BUF_X1 rebuffer19 (.A(_0269_),
    .Z(net29));
 BUF_X2 clone20 (.A(net31),
    .Z(net30));
 BUF_X1 rebuffer21 (.A(_0118_),
    .Z(net31));
 BUF_X2 rebuffer22 (.A(net51),
    .Z(net32));
 BUF_X1 rebuffer23 (.A(_0141_),
    .Z(net33));
 BUF_X4 rebuffer24 (.A(_0076_),
    .Z(net34));
 BUF_X4 rebuffer25 (.A(_0073_),
    .Z(net35));
 BUF_X1 rebuffer26 (.A(_0192_),
    .Z(net36));
 BUF_X1 rebuffer27 (.A(net36),
    .Z(net37));
 BUF_X1 rebuffer28 (.A(_0494_),
    .Z(net38));
 BUF_X1 rebuffer29 (.A(_0242_),
    .Z(net39));
 BUF_X1 rebuffer30 (.A(_0432_),
    .Z(net40));
 BUF_X1 rebuffer31 (.A(_0432_),
    .Z(net41));
 BUF_X2 rebuffer32 (.A(_0844_),
    .Z(net42));
 BUF_X1 rebuffer33 (.A(net42),
    .Z(net43));
 BUF_X4 rebuffer34 (.A(_0303_),
    .Z(net44));
 BUF_X1 rebuffer35 (.A(net67),
    .Z(net45));
 BUF_X4 rebuffer36 (.A(net66),
    .Z(net46));
 BUF_X1 rebuffer37 (.A(_0303_),
    .Z(net47));
 BUF_X1 rebuffer38 (.A(_0398_),
    .Z(net48));
 BUF_X1 rebuffer39 (.A(_0398_),
    .Z(net49));
 BUF_X1 rebuffer40 (.A(_0241_),
    .Z(net50));
 BUF_X2 rebuffer41 (.A(_0241_),
    .Z(net51));
 BUF_X2 rebuffer42 (.A(_0141_),
    .Z(net52));
 BUF_X1 rebuffer43 (.A(net54),
    .Z(net53));
 BUF_X1 rebuffer44 (.A(net55),
    .Z(net54));
 BUF_X1 rebuffer45 (.A(net56),
    .Z(net55));
 BUF_X1 rebuffer46 (.A(net57),
    .Z(net56));
 BUF_X1 rebuffer47 (.A(net58),
    .Z(net57));
 BUF_X1 rebuffer48 (.A(net59),
    .Z(net58));
 BUF_X1 rebuffer49 (.A(net60),
    .Z(net59));
 BUF_X1 rebuffer50 (.A(_0397_),
    .Z(net60));
 BUF_X4 rebuffer51 (.A(_0100_),
    .Z(net61));
 BUF_X2 rebuffer52 (.A(net61),
    .Z(net62));
 BUF_X1 rebuffer53 (.A(_0160_),
    .Z(net63));
 BUF_X1 rebuffer54 (.A(_0269_),
    .Z(net64));
 BUF_X1 rebuffer55 (.A(_0477_),
    .Z(net65));
 BUF_X4 rebuffer56 (.A(_0303_),
    .Z(net66));
 BUF_X1 rebuffer57 (.A(net66),
    .Z(net67));
 BUF_X4 rebuffer58 (.A(_0131_),
    .Z(net68));
 BUF_X2 rebuffer59 (.A(net68),
    .Z(net69));
 BUF_X4 rebuffer60 (.A(_0399_),
    .Z(net70));
 BUF_X2 rebuffer61 (.A(_0400_),
    .Z(net71));
 BUF_X1 rebuffer62 (.A(net71),
    .Z(net72));
 BUF_X1 rebuffer63 (.A(net71),
    .Z(net73));
 BUF_X1 rebuffer64 (.A(net11),
    .Z(net74));
 BUF_X2 rebuffer65 (.A(_0303_),
    .Z(net75));
 BUF_X1 rebuffer20 (.A(_0850_),
    .Z(net76));
 BUF_X1 rebuffer66 (.A(net76),
    .Z(net77));
 BUF_X4 rebuffer67 (.A(_0240_),
    .Z(net78));
 BUF_X4 rebuffer68 (.A(_0223_),
    .Z(net79));
 BUF_X1 rebuffer69 (.A(net79),
    .Z(net80));
 BUF_X1 rebuffer70 (.A(_0221_),
    .Z(net82));
 BUF_X4 rebuffer72 (.A(_0815_),
    .Z(net84));
 BUF_X4 rebuffer73 (.A(_0398_),
    .Z(net85));
 BUF_X2 rebuffer74 (.A(_0148_),
    .Z(net86));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X32 FILLER_0_952 ();
 FILLCELL_X32 FILLER_0_984 ();
 FILLCELL_X32 FILLER_0_1016 ();
 FILLCELL_X32 FILLER_0_1048 ();
 FILLCELL_X32 FILLER_0_1080 ();
 FILLCELL_X32 FILLER_0_1112 ();
 FILLCELL_X32 FILLER_0_1144 ();
 FILLCELL_X32 FILLER_0_1176 ();
 FILLCELL_X32 FILLER_0_1208 ();
 FILLCELL_X16 FILLER_0_1240 ();
 FILLCELL_X4 FILLER_0_1256 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X32 FILLER_0_1775 ();
 FILLCELL_X32 FILLER_0_1807 ();
 FILLCELL_X32 FILLER_0_1839 ();
 FILLCELL_X16 FILLER_0_1871 ();
 FILLCELL_X4 FILLER_0_1887 ();
 FILLCELL_X2 FILLER_0_1891 ();
 FILLCELL_X32 FILLER_0_1894 ();
 FILLCELL_X32 FILLER_0_1926 ();
 FILLCELL_X32 FILLER_0_1958 ();
 FILLCELL_X32 FILLER_0_1990 ();
 FILLCELL_X32 FILLER_0_2022 ();
 FILLCELL_X32 FILLER_0_2054 ();
 FILLCELL_X32 FILLER_0_2086 ();
 FILLCELL_X32 FILLER_0_2118 ();
 FILLCELL_X32 FILLER_0_2150 ();
 FILLCELL_X32 FILLER_0_2182 ();
 FILLCELL_X32 FILLER_0_2214 ();
 FILLCELL_X32 FILLER_0_2246 ();
 FILLCELL_X32 FILLER_0_2278 ();
 FILLCELL_X32 FILLER_0_2310 ();
 FILLCELL_X32 FILLER_0_2342 ();
 FILLCELL_X32 FILLER_0_2374 ();
 FILLCELL_X16 FILLER_0_2406 ();
 FILLCELL_X8 FILLER_0_2422 ();
 FILLCELL_X4 FILLER_0_2430 ();
 FILLCELL_X2 FILLER_0_2434 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X32 FILLER_1_833 ();
 FILLCELL_X32 FILLER_1_865 ();
 FILLCELL_X32 FILLER_1_897 ();
 FILLCELL_X32 FILLER_1_929 ();
 FILLCELL_X32 FILLER_1_961 ();
 FILLCELL_X32 FILLER_1_993 ();
 FILLCELL_X32 FILLER_1_1025 ();
 FILLCELL_X32 FILLER_1_1057 ();
 FILLCELL_X32 FILLER_1_1089 ();
 FILLCELL_X32 FILLER_1_1121 ();
 FILLCELL_X32 FILLER_1_1153 ();
 FILLCELL_X32 FILLER_1_1185 ();
 FILLCELL_X32 FILLER_1_1217 ();
 FILLCELL_X8 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X32 FILLER_1_1776 ();
 FILLCELL_X32 FILLER_1_1808 ();
 FILLCELL_X32 FILLER_1_1840 ();
 FILLCELL_X32 FILLER_1_1872 ();
 FILLCELL_X32 FILLER_1_1904 ();
 FILLCELL_X32 FILLER_1_1936 ();
 FILLCELL_X32 FILLER_1_1968 ();
 FILLCELL_X32 FILLER_1_2000 ();
 FILLCELL_X32 FILLER_1_2032 ();
 FILLCELL_X32 FILLER_1_2064 ();
 FILLCELL_X32 FILLER_1_2096 ();
 FILLCELL_X32 FILLER_1_2128 ();
 FILLCELL_X32 FILLER_1_2160 ();
 FILLCELL_X32 FILLER_1_2192 ();
 FILLCELL_X32 FILLER_1_2224 ();
 FILLCELL_X32 FILLER_1_2256 ();
 FILLCELL_X32 FILLER_1_2288 ();
 FILLCELL_X32 FILLER_1_2320 ();
 FILLCELL_X32 FILLER_1_2352 ();
 FILLCELL_X32 FILLER_1_2384 ();
 FILLCELL_X16 FILLER_1_2416 ();
 FILLCELL_X4 FILLER_1_2432 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X32 FILLER_2_1592 ();
 FILLCELL_X32 FILLER_2_1624 ();
 FILLCELL_X32 FILLER_2_1656 ();
 FILLCELL_X32 FILLER_2_1688 ();
 FILLCELL_X32 FILLER_2_1720 ();
 FILLCELL_X32 FILLER_2_1752 ();
 FILLCELL_X32 FILLER_2_1784 ();
 FILLCELL_X32 FILLER_2_1816 ();
 FILLCELL_X32 FILLER_2_1848 ();
 FILLCELL_X8 FILLER_2_1880 ();
 FILLCELL_X4 FILLER_2_1888 ();
 FILLCELL_X2 FILLER_2_1892 ();
 FILLCELL_X32 FILLER_2_1895 ();
 FILLCELL_X32 FILLER_2_1927 ();
 FILLCELL_X32 FILLER_2_1959 ();
 FILLCELL_X32 FILLER_2_1991 ();
 FILLCELL_X32 FILLER_2_2023 ();
 FILLCELL_X32 FILLER_2_2055 ();
 FILLCELL_X32 FILLER_2_2087 ();
 FILLCELL_X32 FILLER_2_2119 ();
 FILLCELL_X32 FILLER_2_2151 ();
 FILLCELL_X32 FILLER_2_2183 ();
 FILLCELL_X32 FILLER_2_2215 ();
 FILLCELL_X32 FILLER_2_2247 ();
 FILLCELL_X32 FILLER_2_2279 ();
 FILLCELL_X32 FILLER_2_2311 ();
 FILLCELL_X32 FILLER_2_2343 ();
 FILLCELL_X32 FILLER_2_2375 ();
 FILLCELL_X16 FILLER_2_2407 ();
 FILLCELL_X8 FILLER_2_2423 ();
 FILLCELL_X4 FILLER_2_2431 ();
 FILLCELL_X1 FILLER_2_2435 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X32 FILLER_3_1776 ();
 FILLCELL_X32 FILLER_3_1808 ();
 FILLCELL_X32 FILLER_3_1840 ();
 FILLCELL_X32 FILLER_3_1872 ();
 FILLCELL_X32 FILLER_3_1904 ();
 FILLCELL_X32 FILLER_3_1936 ();
 FILLCELL_X32 FILLER_3_1968 ();
 FILLCELL_X32 FILLER_3_2000 ();
 FILLCELL_X32 FILLER_3_2032 ();
 FILLCELL_X32 FILLER_3_2064 ();
 FILLCELL_X32 FILLER_3_2096 ();
 FILLCELL_X32 FILLER_3_2128 ();
 FILLCELL_X32 FILLER_3_2160 ();
 FILLCELL_X32 FILLER_3_2192 ();
 FILLCELL_X32 FILLER_3_2224 ();
 FILLCELL_X32 FILLER_3_2256 ();
 FILLCELL_X32 FILLER_3_2288 ();
 FILLCELL_X32 FILLER_3_2320 ();
 FILLCELL_X32 FILLER_3_2352 ();
 FILLCELL_X32 FILLER_3_2384 ();
 FILLCELL_X16 FILLER_3_2416 ();
 FILLCELL_X4 FILLER_3_2432 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X32 FILLER_4_1592 ();
 FILLCELL_X32 FILLER_4_1624 ();
 FILLCELL_X32 FILLER_4_1656 ();
 FILLCELL_X32 FILLER_4_1688 ();
 FILLCELL_X32 FILLER_4_1720 ();
 FILLCELL_X32 FILLER_4_1752 ();
 FILLCELL_X32 FILLER_4_1784 ();
 FILLCELL_X32 FILLER_4_1816 ();
 FILLCELL_X32 FILLER_4_1848 ();
 FILLCELL_X8 FILLER_4_1880 ();
 FILLCELL_X4 FILLER_4_1888 ();
 FILLCELL_X2 FILLER_4_1892 ();
 FILLCELL_X32 FILLER_4_1895 ();
 FILLCELL_X32 FILLER_4_1927 ();
 FILLCELL_X32 FILLER_4_1959 ();
 FILLCELL_X32 FILLER_4_1991 ();
 FILLCELL_X32 FILLER_4_2023 ();
 FILLCELL_X32 FILLER_4_2055 ();
 FILLCELL_X32 FILLER_4_2087 ();
 FILLCELL_X32 FILLER_4_2119 ();
 FILLCELL_X32 FILLER_4_2151 ();
 FILLCELL_X32 FILLER_4_2183 ();
 FILLCELL_X32 FILLER_4_2215 ();
 FILLCELL_X32 FILLER_4_2247 ();
 FILLCELL_X32 FILLER_4_2279 ();
 FILLCELL_X32 FILLER_4_2311 ();
 FILLCELL_X32 FILLER_4_2343 ();
 FILLCELL_X32 FILLER_4_2375 ();
 FILLCELL_X16 FILLER_4_2407 ();
 FILLCELL_X8 FILLER_4_2423 ();
 FILLCELL_X4 FILLER_4_2431 ();
 FILLCELL_X1 FILLER_4_2435 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X32 FILLER_5_1776 ();
 FILLCELL_X32 FILLER_5_1808 ();
 FILLCELL_X32 FILLER_5_1840 ();
 FILLCELL_X32 FILLER_5_1872 ();
 FILLCELL_X32 FILLER_5_1904 ();
 FILLCELL_X32 FILLER_5_1936 ();
 FILLCELL_X32 FILLER_5_1968 ();
 FILLCELL_X32 FILLER_5_2000 ();
 FILLCELL_X32 FILLER_5_2032 ();
 FILLCELL_X32 FILLER_5_2064 ();
 FILLCELL_X32 FILLER_5_2096 ();
 FILLCELL_X32 FILLER_5_2128 ();
 FILLCELL_X32 FILLER_5_2160 ();
 FILLCELL_X32 FILLER_5_2192 ();
 FILLCELL_X32 FILLER_5_2224 ();
 FILLCELL_X32 FILLER_5_2256 ();
 FILLCELL_X32 FILLER_5_2288 ();
 FILLCELL_X32 FILLER_5_2320 ();
 FILLCELL_X32 FILLER_5_2352 ();
 FILLCELL_X32 FILLER_5_2384 ();
 FILLCELL_X16 FILLER_5_2416 ();
 FILLCELL_X4 FILLER_5_2432 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X32 FILLER_6_1592 ();
 FILLCELL_X32 FILLER_6_1624 ();
 FILLCELL_X32 FILLER_6_1656 ();
 FILLCELL_X32 FILLER_6_1688 ();
 FILLCELL_X32 FILLER_6_1720 ();
 FILLCELL_X32 FILLER_6_1752 ();
 FILLCELL_X32 FILLER_6_1784 ();
 FILLCELL_X32 FILLER_6_1816 ();
 FILLCELL_X32 FILLER_6_1848 ();
 FILLCELL_X8 FILLER_6_1880 ();
 FILLCELL_X4 FILLER_6_1888 ();
 FILLCELL_X2 FILLER_6_1892 ();
 FILLCELL_X32 FILLER_6_1895 ();
 FILLCELL_X32 FILLER_6_1927 ();
 FILLCELL_X32 FILLER_6_1959 ();
 FILLCELL_X32 FILLER_6_1991 ();
 FILLCELL_X32 FILLER_6_2023 ();
 FILLCELL_X32 FILLER_6_2055 ();
 FILLCELL_X32 FILLER_6_2087 ();
 FILLCELL_X32 FILLER_6_2119 ();
 FILLCELL_X32 FILLER_6_2151 ();
 FILLCELL_X32 FILLER_6_2183 ();
 FILLCELL_X32 FILLER_6_2215 ();
 FILLCELL_X32 FILLER_6_2247 ();
 FILLCELL_X32 FILLER_6_2279 ();
 FILLCELL_X32 FILLER_6_2311 ();
 FILLCELL_X32 FILLER_6_2343 ();
 FILLCELL_X32 FILLER_6_2375 ();
 FILLCELL_X16 FILLER_6_2407 ();
 FILLCELL_X8 FILLER_6_2423 ();
 FILLCELL_X4 FILLER_6_2431 ();
 FILLCELL_X1 FILLER_6_2435 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X32 FILLER_7_1776 ();
 FILLCELL_X32 FILLER_7_1808 ();
 FILLCELL_X32 FILLER_7_1840 ();
 FILLCELL_X32 FILLER_7_1872 ();
 FILLCELL_X32 FILLER_7_1904 ();
 FILLCELL_X32 FILLER_7_1936 ();
 FILLCELL_X32 FILLER_7_1968 ();
 FILLCELL_X32 FILLER_7_2000 ();
 FILLCELL_X32 FILLER_7_2032 ();
 FILLCELL_X32 FILLER_7_2064 ();
 FILLCELL_X32 FILLER_7_2096 ();
 FILLCELL_X32 FILLER_7_2128 ();
 FILLCELL_X32 FILLER_7_2160 ();
 FILLCELL_X32 FILLER_7_2192 ();
 FILLCELL_X32 FILLER_7_2224 ();
 FILLCELL_X32 FILLER_7_2256 ();
 FILLCELL_X32 FILLER_7_2288 ();
 FILLCELL_X32 FILLER_7_2320 ();
 FILLCELL_X32 FILLER_7_2352 ();
 FILLCELL_X32 FILLER_7_2384 ();
 FILLCELL_X16 FILLER_7_2416 ();
 FILLCELL_X4 FILLER_7_2432 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X32 FILLER_8_1592 ();
 FILLCELL_X32 FILLER_8_1624 ();
 FILLCELL_X32 FILLER_8_1656 ();
 FILLCELL_X32 FILLER_8_1688 ();
 FILLCELL_X32 FILLER_8_1720 ();
 FILLCELL_X32 FILLER_8_1752 ();
 FILLCELL_X32 FILLER_8_1784 ();
 FILLCELL_X32 FILLER_8_1816 ();
 FILLCELL_X32 FILLER_8_1848 ();
 FILLCELL_X8 FILLER_8_1880 ();
 FILLCELL_X4 FILLER_8_1888 ();
 FILLCELL_X2 FILLER_8_1892 ();
 FILLCELL_X32 FILLER_8_1895 ();
 FILLCELL_X32 FILLER_8_1927 ();
 FILLCELL_X32 FILLER_8_1959 ();
 FILLCELL_X32 FILLER_8_1991 ();
 FILLCELL_X32 FILLER_8_2023 ();
 FILLCELL_X32 FILLER_8_2055 ();
 FILLCELL_X32 FILLER_8_2087 ();
 FILLCELL_X32 FILLER_8_2119 ();
 FILLCELL_X32 FILLER_8_2151 ();
 FILLCELL_X32 FILLER_8_2183 ();
 FILLCELL_X32 FILLER_8_2215 ();
 FILLCELL_X32 FILLER_8_2247 ();
 FILLCELL_X32 FILLER_8_2279 ();
 FILLCELL_X32 FILLER_8_2311 ();
 FILLCELL_X32 FILLER_8_2343 ();
 FILLCELL_X32 FILLER_8_2375 ();
 FILLCELL_X16 FILLER_8_2407 ();
 FILLCELL_X8 FILLER_8_2423 ();
 FILLCELL_X4 FILLER_8_2431 ();
 FILLCELL_X1 FILLER_8_2435 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X32 FILLER_9_1776 ();
 FILLCELL_X32 FILLER_9_1808 ();
 FILLCELL_X32 FILLER_9_1840 ();
 FILLCELL_X32 FILLER_9_1872 ();
 FILLCELL_X32 FILLER_9_1904 ();
 FILLCELL_X32 FILLER_9_1936 ();
 FILLCELL_X32 FILLER_9_1968 ();
 FILLCELL_X32 FILLER_9_2000 ();
 FILLCELL_X32 FILLER_9_2032 ();
 FILLCELL_X32 FILLER_9_2064 ();
 FILLCELL_X32 FILLER_9_2096 ();
 FILLCELL_X32 FILLER_9_2128 ();
 FILLCELL_X32 FILLER_9_2160 ();
 FILLCELL_X32 FILLER_9_2192 ();
 FILLCELL_X32 FILLER_9_2224 ();
 FILLCELL_X32 FILLER_9_2256 ();
 FILLCELL_X32 FILLER_9_2288 ();
 FILLCELL_X32 FILLER_9_2320 ();
 FILLCELL_X32 FILLER_9_2352 ();
 FILLCELL_X32 FILLER_9_2384 ();
 FILLCELL_X16 FILLER_9_2416 ();
 FILLCELL_X4 FILLER_9_2432 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X32 FILLER_10_1592 ();
 FILLCELL_X32 FILLER_10_1624 ();
 FILLCELL_X32 FILLER_10_1656 ();
 FILLCELL_X32 FILLER_10_1688 ();
 FILLCELL_X32 FILLER_10_1720 ();
 FILLCELL_X32 FILLER_10_1752 ();
 FILLCELL_X32 FILLER_10_1784 ();
 FILLCELL_X32 FILLER_10_1816 ();
 FILLCELL_X32 FILLER_10_1848 ();
 FILLCELL_X8 FILLER_10_1880 ();
 FILLCELL_X4 FILLER_10_1888 ();
 FILLCELL_X2 FILLER_10_1892 ();
 FILLCELL_X32 FILLER_10_1895 ();
 FILLCELL_X32 FILLER_10_1927 ();
 FILLCELL_X32 FILLER_10_1959 ();
 FILLCELL_X32 FILLER_10_1991 ();
 FILLCELL_X32 FILLER_10_2023 ();
 FILLCELL_X32 FILLER_10_2055 ();
 FILLCELL_X32 FILLER_10_2087 ();
 FILLCELL_X32 FILLER_10_2119 ();
 FILLCELL_X32 FILLER_10_2151 ();
 FILLCELL_X32 FILLER_10_2183 ();
 FILLCELL_X32 FILLER_10_2215 ();
 FILLCELL_X32 FILLER_10_2247 ();
 FILLCELL_X32 FILLER_10_2279 ();
 FILLCELL_X32 FILLER_10_2311 ();
 FILLCELL_X32 FILLER_10_2343 ();
 FILLCELL_X32 FILLER_10_2375 ();
 FILLCELL_X16 FILLER_10_2407 ();
 FILLCELL_X8 FILLER_10_2423 ();
 FILLCELL_X4 FILLER_10_2431 ();
 FILLCELL_X1 FILLER_10_2435 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X32 FILLER_11_1776 ();
 FILLCELL_X32 FILLER_11_1808 ();
 FILLCELL_X32 FILLER_11_1840 ();
 FILLCELL_X32 FILLER_11_1872 ();
 FILLCELL_X32 FILLER_11_1904 ();
 FILLCELL_X32 FILLER_11_1936 ();
 FILLCELL_X32 FILLER_11_1968 ();
 FILLCELL_X32 FILLER_11_2000 ();
 FILLCELL_X32 FILLER_11_2032 ();
 FILLCELL_X32 FILLER_11_2064 ();
 FILLCELL_X32 FILLER_11_2096 ();
 FILLCELL_X32 FILLER_11_2128 ();
 FILLCELL_X32 FILLER_11_2160 ();
 FILLCELL_X32 FILLER_11_2192 ();
 FILLCELL_X32 FILLER_11_2224 ();
 FILLCELL_X32 FILLER_11_2256 ();
 FILLCELL_X32 FILLER_11_2288 ();
 FILLCELL_X32 FILLER_11_2320 ();
 FILLCELL_X32 FILLER_11_2352 ();
 FILLCELL_X32 FILLER_11_2384 ();
 FILLCELL_X16 FILLER_11_2416 ();
 FILLCELL_X4 FILLER_11_2432 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X32 FILLER_12_1784 ();
 FILLCELL_X32 FILLER_12_1816 ();
 FILLCELL_X32 FILLER_12_1848 ();
 FILLCELL_X8 FILLER_12_1880 ();
 FILLCELL_X4 FILLER_12_1888 ();
 FILLCELL_X2 FILLER_12_1892 ();
 FILLCELL_X32 FILLER_12_1895 ();
 FILLCELL_X32 FILLER_12_1927 ();
 FILLCELL_X32 FILLER_12_1959 ();
 FILLCELL_X32 FILLER_12_1991 ();
 FILLCELL_X32 FILLER_12_2023 ();
 FILLCELL_X32 FILLER_12_2055 ();
 FILLCELL_X32 FILLER_12_2087 ();
 FILLCELL_X32 FILLER_12_2119 ();
 FILLCELL_X32 FILLER_12_2151 ();
 FILLCELL_X32 FILLER_12_2183 ();
 FILLCELL_X32 FILLER_12_2215 ();
 FILLCELL_X32 FILLER_12_2247 ();
 FILLCELL_X32 FILLER_12_2279 ();
 FILLCELL_X32 FILLER_12_2311 ();
 FILLCELL_X32 FILLER_12_2343 ();
 FILLCELL_X32 FILLER_12_2375 ();
 FILLCELL_X16 FILLER_12_2407 ();
 FILLCELL_X8 FILLER_12_2423 ();
 FILLCELL_X4 FILLER_12_2431 ();
 FILLCELL_X1 FILLER_12_2435 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X32 FILLER_13_1776 ();
 FILLCELL_X32 FILLER_13_1808 ();
 FILLCELL_X32 FILLER_13_1840 ();
 FILLCELL_X32 FILLER_13_1872 ();
 FILLCELL_X32 FILLER_13_1904 ();
 FILLCELL_X32 FILLER_13_1936 ();
 FILLCELL_X32 FILLER_13_1968 ();
 FILLCELL_X32 FILLER_13_2000 ();
 FILLCELL_X32 FILLER_13_2032 ();
 FILLCELL_X32 FILLER_13_2064 ();
 FILLCELL_X32 FILLER_13_2096 ();
 FILLCELL_X32 FILLER_13_2128 ();
 FILLCELL_X32 FILLER_13_2160 ();
 FILLCELL_X32 FILLER_13_2192 ();
 FILLCELL_X32 FILLER_13_2224 ();
 FILLCELL_X32 FILLER_13_2256 ();
 FILLCELL_X32 FILLER_13_2288 ();
 FILLCELL_X32 FILLER_13_2320 ();
 FILLCELL_X32 FILLER_13_2352 ();
 FILLCELL_X32 FILLER_13_2384 ();
 FILLCELL_X16 FILLER_13_2416 ();
 FILLCELL_X4 FILLER_13_2432 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X32 FILLER_14_1784 ();
 FILLCELL_X32 FILLER_14_1816 ();
 FILLCELL_X32 FILLER_14_1848 ();
 FILLCELL_X8 FILLER_14_1880 ();
 FILLCELL_X4 FILLER_14_1888 ();
 FILLCELL_X2 FILLER_14_1892 ();
 FILLCELL_X32 FILLER_14_1895 ();
 FILLCELL_X32 FILLER_14_1927 ();
 FILLCELL_X32 FILLER_14_1959 ();
 FILLCELL_X32 FILLER_14_1991 ();
 FILLCELL_X32 FILLER_14_2023 ();
 FILLCELL_X32 FILLER_14_2055 ();
 FILLCELL_X32 FILLER_14_2087 ();
 FILLCELL_X32 FILLER_14_2119 ();
 FILLCELL_X32 FILLER_14_2151 ();
 FILLCELL_X32 FILLER_14_2183 ();
 FILLCELL_X32 FILLER_14_2215 ();
 FILLCELL_X32 FILLER_14_2247 ();
 FILLCELL_X32 FILLER_14_2279 ();
 FILLCELL_X32 FILLER_14_2311 ();
 FILLCELL_X32 FILLER_14_2343 ();
 FILLCELL_X32 FILLER_14_2375 ();
 FILLCELL_X16 FILLER_14_2407 ();
 FILLCELL_X8 FILLER_14_2423 ();
 FILLCELL_X4 FILLER_14_2431 ();
 FILLCELL_X1 FILLER_14_2435 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X32 FILLER_15_1776 ();
 FILLCELL_X32 FILLER_15_1808 ();
 FILLCELL_X32 FILLER_15_1840 ();
 FILLCELL_X32 FILLER_15_1872 ();
 FILLCELL_X32 FILLER_15_1904 ();
 FILLCELL_X32 FILLER_15_1936 ();
 FILLCELL_X32 FILLER_15_1968 ();
 FILLCELL_X32 FILLER_15_2000 ();
 FILLCELL_X32 FILLER_15_2032 ();
 FILLCELL_X32 FILLER_15_2064 ();
 FILLCELL_X32 FILLER_15_2096 ();
 FILLCELL_X32 FILLER_15_2128 ();
 FILLCELL_X32 FILLER_15_2160 ();
 FILLCELL_X32 FILLER_15_2192 ();
 FILLCELL_X32 FILLER_15_2224 ();
 FILLCELL_X32 FILLER_15_2256 ();
 FILLCELL_X32 FILLER_15_2288 ();
 FILLCELL_X32 FILLER_15_2320 ();
 FILLCELL_X32 FILLER_15_2352 ();
 FILLCELL_X32 FILLER_15_2384 ();
 FILLCELL_X16 FILLER_15_2416 ();
 FILLCELL_X4 FILLER_15_2432 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X32 FILLER_16_1784 ();
 FILLCELL_X32 FILLER_16_1816 ();
 FILLCELL_X32 FILLER_16_1848 ();
 FILLCELL_X8 FILLER_16_1880 ();
 FILLCELL_X4 FILLER_16_1888 ();
 FILLCELL_X2 FILLER_16_1892 ();
 FILLCELL_X32 FILLER_16_1895 ();
 FILLCELL_X32 FILLER_16_1927 ();
 FILLCELL_X32 FILLER_16_1959 ();
 FILLCELL_X32 FILLER_16_1991 ();
 FILLCELL_X32 FILLER_16_2023 ();
 FILLCELL_X32 FILLER_16_2055 ();
 FILLCELL_X32 FILLER_16_2087 ();
 FILLCELL_X32 FILLER_16_2119 ();
 FILLCELL_X32 FILLER_16_2151 ();
 FILLCELL_X32 FILLER_16_2183 ();
 FILLCELL_X32 FILLER_16_2215 ();
 FILLCELL_X32 FILLER_16_2247 ();
 FILLCELL_X32 FILLER_16_2279 ();
 FILLCELL_X32 FILLER_16_2311 ();
 FILLCELL_X32 FILLER_16_2343 ();
 FILLCELL_X32 FILLER_16_2375 ();
 FILLCELL_X16 FILLER_16_2407 ();
 FILLCELL_X8 FILLER_16_2423 ();
 FILLCELL_X4 FILLER_16_2431 ();
 FILLCELL_X1 FILLER_16_2435 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X32 FILLER_17_1776 ();
 FILLCELL_X32 FILLER_17_1808 ();
 FILLCELL_X32 FILLER_17_1840 ();
 FILLCELL_X32 FILLER_17_1872 ();
 FILLCELL_X32 FILLER_17_1904 ();
 FILLCELL_X32 FILLER_17_1936 ();
 FILLCELL_X32 FILLER_17_1968 ();
 FILLCELL_X32 FILLER_17_2000 ();
 FILLCELL_X32 FILLER_17_2032 ();
 FILLCELL_X32 FILLER_17_2064 ();
 FILLCELL_X32 FILLER_17_2096 ();
 FILLCELL_X32 FILLER_17_2128 ();
 FILLCELL_X32 FILLER_17_2160 ();
 FILLCELL_X32 FILLER_17_2192 ();
 FILLCELL_X32 FILLER_17_2224 ();
 FILLCELL_X32 FILLER_17_2256 ();
 FILLCELL_X32 FILLER_17_2288 ();
 FILLCELL_X32 FILLER_17_2320 ();
 FILLCELL_X32 FILLER_17_2352 ();
 FILLCELL_X32 FILLER_17_2384 ();
 FILLCELL_X16 FILLER_17_2416 ();
 FILLCELL_X4 FILLER_17_2432 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X32 FILLER_18_1784 ();
 FILLCELL_X32 FILLER_18_1816 ();
 FILLCELL_X32 FILLER_18_1848 ();
 FILLCELL_X8 FILLER_18_1880 ();
 FILLCELL_X4 FILLER_18_1888 ();
 FILLCELL_X2 FILLER_18_1892 ();
 FILLCELL_X32 FILLER_18_1895 ();
 FILLCELL_X32 FILLER_18_1927 ();
 FILLCELL_X32 FILLER_18_1959 ();
 FILLCELL_X32 FILLER_18_1991 ();
 FILLCELL_X32 FILLER_18_2023 ();
 FILLCELL_X32 FILLER_18_2055 ();
 FILLCELL_X32 FILLER_18_2087 ();
 FILLCELL_X32 FILLER_18_2119 ();
 FILLCELL_X32 FILLER_18_2151 ();
 FILLCELL_X32 FILLER_18_2183 ();
 FILLCELL_X32 FILLER_18_2215 ();
 FILLCELL_X32 FILLER_18_2247 ();
 FILLCELL_X32 FILLER_18_2279 ();
 FILLCELL_X32 FILLER_18_2311 ();
 FILLCELL_X32 FILLER_18_2343 ();
 FILLCELL_X32 FILLER_18_2375 ();
 FILLCELL_X16 FILLER_18_2407 ();
 FILLCELL_X8 FILLER_18_2423 ();
 FILLCELL_X4 FILLER_18_2431 ();
 FILLCELL_X1 FILLER_18_2435 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X32 FILLER_19_1776 ();
 FILLCELL_X32 FILLER_19_1808 ();
 FILLCELL_X32 FILLER_19_1840 ();
 FILLCELL_X32 FILLER_19_1872 ();
 FILLCELL_X32 FILLER_19_1904 ();
 FILLCELL_X32 FILLER_19_1936 ();
 FILLCELL_X32 FILLER_19_1968 ();
 FILLCELL_X32 FILLER_19_2000 ();
 FILLCELL_X32 FILLER_19_2032 ();
 FILLCELL_X32 FILLER_19_2064 ();
 FILLCELL_X32 FILLER_19_2096 ();
 FILLCELL_X32 FILLER_19_2128 ();
 FILLCELL_X32 FILLER_19_2160 ();
 FILLCELL_X32 FILLER_19_2192 ();
 FILLCELL_X32 FILLER_19_2224 ();
 FILLCELL_X32 FILLER_19_2256 ();
 FILLCELL_X32 FILLER_19_2288 ();
 FILLCELL_X32 FILLER_19_2320 ();
 FILLCELL_X32 FILLER_19_2352 ();
 FILLCELL_X32 FILLER_19_2384 ();
 FILLCELL_X16 FILLER_19_2416 ();
 FILLCELL_X4 FILLER_19_2432 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X32 FILLER_20_1784 ();
 FILLCELL_X32 FILLER_20_1816 ();
 FILLCELL_X32 FILLER_20_1848 ();
 FILLCELL_X8 FILLER_20_1880 ();
 FILLCELL_X4 FILLER_20_1888 ();
 FILLCELL_X2 FILLER_20_1892 ();
 FILLCELL_X32 FILLER_20_1895 ();
 FILLCELL_X32 FILLER_20_1927 ();
 FILLCELL_X32 FILLER_20_1959 ();
 FILLCELL_X32 FILLER_20_1991 ();
 FILLCELL_X32 FILLER_20_2023 ();
 FILLCELL_X32 FILLER_20_2055 ();
 FILLCELL_X32 FILLER_20_2087 ();
 FILLCELL_X32 FILLER_20_2119 ();
 FILLCELL_X32 FILLER_20_2151 ();
 FILLCELL_X32 FILLER_20_2183 ();
 FILLCELL_X32 FILLER_20_2215 ();
 FILLCELL_X32 FILLER_20_2247 ();
 FILLCELL_X32 FILLER_20_2279 ();
 FILLCELL_X32 FILLER_20_2311 ();
 FILLCELL_X32 FILLER_20_2343 ();
 FILLCELL_X32 FILLER_20_2375 ();
 FILLCELL_X16 FILLER_20_2407 ();
 FILLCELL_X8 FILLER_20_2423 ();
 FILLCELL_X4 FILLER_20_2431 ();
 FILLCELL_X1 FILLER_20_2435 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X32 FILLER_21_1776 ();
 FILLCELL_X32 FILLER_21_1808 ();
 FILLCELL_X32 FILLER_21_1840 ();
 FILLCELL_X32 FILLER_21_1872 ();
 FILLCELL_X32 FILLER_21_1904 ();
 FILLCELL_X32 FILLER_21_1936 ();
 FILLCELL_X32 FILLER_21_1968 ();
 FILLCELL_X32 FILLER_21_2000 ();
 FILLCELL_X32 FILLER_21_2032 ();
 FILLCELL_X32 FILLER_21_2064 ();
 FILLCELL_X32 FILLER_21_2096 ();
 FILLCELL_X32 FILLER_21_2128 ();
 FILLCELL_X32 FILLER_21_2160 ();
 FILLCELL_X32 FILLER_21_2192 ();
 FILLCELL_X32 FILLER_21_2224 ();
 FILLCELL_X32 FILLER_21_2256 ();
 FILLCELL_X32 FILLER_21_2288 ();
 FILLCELL_X32 FILLER_21_2320 ();
 FILLCELL_X32 FILLER_21_2352 ();
 FILLCELL_X32 FILLER_21_2384 ();
 FILLCELL_X16 FILLER_21_2416 ();
 FILLCELL_X4 FILLER_21_2432 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X32 FILLER_22_1784 ();
 FILLCELL_X32 FILLER_22_1816 ();
 FILLCELL_X32 FILLER_22_1848 ();
 FILLCELL_X8 FILLER_22_1880 ();
 FILLCELL_X4 FILLER_22_1888 ();
 FILLCELL_X2 FILLER_22_1892 ();
 FILLCELL_X32 FILLER_22_1895 ();
 FILLCELL_X32 FILLER_22_1927 ();
 FILLCELL_X32 FILLER_22_1959 ();
 FILLCELL_X32 FILLER_22_1991 ();
 FILLCELL_X32 FILLER_22_2023 ();
 FILLCELL_X32 FILLER_22_2055 ();
 FILLCELL_X32 FILLER_22_2087 ();
 FILLCELL_X32 FILLER_22_2119 ();
 FILLCELL_X32 FILLER_22_2151 ();
 FILLCELL_X32 FILLER_22_2183 ();
 FILLCELL_X32 FILLER_22_2215 ();
 FILLCELL_X32 FILLER_22_2247 ();
 FILLCELL_X32 FILLER_22_2279 ();
 FILLCELL_X32 FILLER_22_2311 ();
 FILLCELL_X32 FILLER_22_2343 ();
 FILLCELL_X32 FILLER_22_2375 ();
 FILLCELL_X16 FILLER_22_2407 ();
 FILLCELL_X8 FILLER_22_2423 ();
 FILLCELL_X4 FILLER_22_2431 ();
 FILLCELL_X1 FILLER_22_2435 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X32 FILLER_23_1776 ();
 FILLCELL_X32 FILLER_23_1808 ();
 FILLCELL_X32 FILLER_23_1840 ();
 FILLCELL_X32 FILLER_23_1872 ();
 FILLCELL_X32 FILLER_23_1904 ();
 FILLCELL_X32 FILLER_23_1936 ();
 FILLCELL_X32 FILLER_23_1968 ();
 FILLCELL_X32 FILLER_23_2000 ();
 FILLCELL_X32 FILLER_23_2032 ();
 FILLCELL_X32 FILLER_23_2064 ();
 FILLCELL_X32 FILLER_23_2096 ();
 FILLCELL_X32 FILLER_23_2128 ();
 FILLCELL_X32 FILLER_23_2160 ();
 FILLCELL_X32 FILLER_23_2192 ();
 FILLCELL_X32 FILLER_23_2224 ();
 FILLCELL_X32 FILLER_23_2256 ();
 FILLCELL_X32 FILLER_23_2288 ();
 FILLCELL_X32 FILLER_23_2320 ();
 FILLCELL_X32 FILLER_23_2352 ();
 FILLCELL_X32 FILLER_23_2384 ();
 FILLCELL_X16 FILLER_23_2416 ();
 FILLCELL_X4 FILLER_23_2432 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X32 FILLER_24_1784 ();
 FILLCELL_X32 FILLER_24_1816 ();
 FILLCELL_X32 FILLER_24_1848 ();
 FILLCELL_X8 FILLER_24_1880 ();
 FILLCELL_X4 FILLER_24_1888 ();
 FILLCELL_X2 FILLER_24_1892 ();
 FILLCELL_X32 FILLER_24_1895 ();
 FILLCELL_X32 FILLER_24_1927 ();
 FILLCELL_X32 FILLER_24_1959 ();
 FILLCELL_X32 FILLER_24_1991 ();
 FILLCELL_X32 FILLER_24_2023 ();
 FILLCELL_X32 FILLER_24_2055 ();
 FILLCELL_X32 FILLER_24_2087 ();
 FILLCELL_X32 FILLER_24_2119 ();
 FILLCELL_X32 FILLER_24_2151 ();
 FILLCELL_X32 FILLER_24_2183 ();
 FILLCELL_X32 FILLER_24_2215 ();
 FILLCELL_X32 FILLER_24_2247 ();
 FILLCELL_X32 FILLER_24_2279 ();
 FILLCELL_X32 FILLER_24_2311 ();
 FILLCELL_X32 FILLER_24_2343 ();
 FILLCELL_X32 FILLER_24_2375 ();
 FILLCELL_X16 FILLER_24_2407 ();
 FILLCELL_X8 FILLER_24_2423 ();
 FILLCELL_X4 FILLER_24_2431 ();
 FILLCELL_X1 FILLER_24_2435 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X32 FILLER_25_1776 ();
 FILLCELL_X32 FILLER_25_1808 ();
 FILLCELL_X32 FILLER_25_1840 ();
 FILLCELL_X32 FILLER_25_1872 ();
 FILLCELL_X32 FILLER_25_1904 ();
 FILLCELL_X32 FILLER_25_1936 ();
 FILLCELL_X32 FILLER_25_1968 ();
 FILLCELL_X32 FILLER_25_2000 ();
 FILLCELL_X32 FILLER_25_2032 ();
 FILLCELL_X32 FILLER_25_2064 ();
 FILLCELL_X32 FILLER_25_2096 ();
 FILLCELL_X32 FILLER_25_2128 ();
 FILLCELL_X32 FILLER_25_2160 ();
 FILLCELL_X32 FILLER_25_2192 ();
 FILLCELL_X32 FILLER_25_2224 ();
 FILLCELL_X32 FILLER_25_2256 ();
 FILLCELL_X32 FILLER_25_2288 ();
 FILLCELL_X32 FILLER_25_2320 ();
 FILLCELL_X32 FILLER_25_2352 ();
 FILLCELL_X32 FILLER_25_2384 ();
 FILLCELL_X16 FILLER_25_2416 ();
 FILLCELL_X4 FILLER_25_2432 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X32 FILLER_26_1784 ();
 FILLCELL_X32 FILLER_26_1816 ();
 FILLCELL_X32 FILLER_26_1848 ();
 FILLCELL_X8 FILLER_26_1880 ();
 FILLCELL_X4 FILLER_26_1888 ();
 FILLCELL_X2 FILLER_26_1892 ();
 FILLCELL_X32 FILLER_26_1895 ();
 FILLCELL_X32 FILLER_26_1927 ();
 FILLCELL_X32 FILLER_26_1959 ();
 FILLCELL_X32 FILLER_26_1991 ();
 FILLCELL_X32 FILLER_26_2023 ();
 FILLCELL_X32 FILLER_26_2055 ();
 FILLCELL_X32 FILLER_26_2087 ();
 FILLCELL_X32 FILLER_26_2119 ();
 FILLCELL_X32 FILLER_26_2151 ();
 FILLCELL_X32 FILLER_26_2183 ();
 FILLCELL_X32 FILLER_26_2215 ();
 FILLCELL_X32 FILLER_26_2247 ();
 FILLCELL_X32 FILLER_26_2279 ();
 FILLCELL_X32 FILLER_26_2311 ();
 FILLCELL_X32 FILLER_26_2343 ();
 FILLCELL_X32 FILLER_26_2375 ();
 FILLCELL_X16 FILLER_26_2407 ();
 FILLCELL_X8 FILLER_26_2423 ();
 FILLCELL_X4 FILLER_26_2431 ();
 FILLCELL_X1 FILLER_26_2435 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X32 FILLER_27_1776 ();
 FILLCELL_X32 FILLER_27_1808 ();
 FILLCELL_X32 FILLER_27_1840 ();
 FILLCELL_X32 FILLER_27_1872 ();
 FILLCELL_X32 FILLER_27_1904 ();
 FILLCELL_X32 FILLER_27_1936 ();
 FILLCELL_X32 FILLER_27_1968 ();
 FILLCELL_X32 FILLER_27_2000 ();
 FILLCELL_X32 FILLER_27_2032 ();
 FILLCELL_X32 FILLER_27_2064 ();
 FILLCELL_X32 FILLER_27_2096 ();
 FILLCELL_X32 FILLER_27_2128 ();
 FILLCELL_X32 FILLER_27_2160 ();
 FILLCELL_X32 FILLER_27_2192 ();
 FILLCELL_X32 FILLER_27_2224 ();
 FILLCELL_X32 FILLER_27_2256 ();
 FILLCELL_X32 FILLER_27_2288 ();
 FILLCELL_X32 FILLER_27_2320 ();
 FILLCELL_X32 FILLER_27_2352 ();
 FILLCELL_X32 FILLER_27_2384 ();
 FILLCELL_X16 FILLER_27_2416 ();
 FILLCELL_X4 FILLER_27_2432 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X32 FILLER_28_1784 ();
 FILLCELL_X32 FILLER_28_1816 ();
 FILLCELL_X32 FILLER_28_1848 ();
 FILLCELL_X8 FILLER_28_1880 ();
 FILLCELL_X4 FILLER_28_1888 ();
 FILLCELL_X2 FILLER_28_1892 ();
 FILLCELL_X32 FILLER_28_1895 ();
 FILLCELL_X32 FILLER_28_1927 ();
 FILLCELL_X32 FILLER_28_1959 ();
 FILLCELL_X32 FILLER_28_1991 ();
 FILLCELL_X32 FILLER_28_2023 ();
 FILLCELL_X32 FILLER_28_2055 ();
 FILLCELL_X32 FILLER_28_2087 ();
 FILLCELL_X32 FILLER_28_2119 ();
 FILLCELL_X32 FILLER_28_2151 ();
 FILLCELL_X32 FILLER_28_2183 ();
 FILLCELL_X32 FILLER_28_2215 ();
 FILLCELL_X32 FILLER_28_2247 ();
 FILLCELL_X32 FILLER_28_2279 ();
 FILLCELL_X32 FILLER_28_2311 ();
 FILLCELL_X32 FILLER_28_2343 ();
 FILLCELL_X32 FILLER_28_2375 ();
 FILLCELL_X16 FILLER_28_2407 ();
 FILLCELL_X8 FILLER_28_2423 ();
 FILLCELL_X4 FILLER_28_2431 ();
 FILLCELL_X1 FILLER_28_2435 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X32 FILLER_29_1776 ();
 FILLCELL_X32 FILLER_29_1808 ();
 FILLCELL_X32 FILLER_29_1840 ();
 FILLCELL_X32 FILLER_29_1872 ();
 FILLCELL_X32 FILLER_29_1904 ();
 FILLCELL_X32 FILLER_29_1936 ();
 FILLCELL_X32 FILLER_29_1968 ();
 FILLCELL_X32 FILLER_29_2000 ();
 FILLCELL_X32 FILLER_29_2032 ();
 FILLCELL_X32 FILLER_29_2064 ();
 FILLCELL_X32 FILLER_29_2096 ();
 FILLCELL_X32 FILLER_29_2128 ();
 FILLCELL_X32 FILLER_29_2160 ();
 FILLCELL_X32 FILLER_29_2192 ();
 FILLCELL_X32 FILLER_29_2224 ();
 FILLCELL_X32 FILLER_29_2256 ();
 FILLCELL_X32 FILLER_29_2288 ();
 FILLCELL_X32 FILLER_29_2320 ();
 FILLCELL_X32 FILLER_29_2352 ();
 FILLCELL_X32 FILLER_29_2384 ();
 FILLCELL_X16 FILLER_29_2416 ();
 FILLCELL_X4 FILLER_29_2432 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X32 FILLER_30_1784 ();
 FILLCELL_X32 FILLER_30_1816 ();
 FILLCELL_X32 FILLER_30_1848 ();
 FILLCELL_X8 FILLER_30_1880 ();
 FILLCELL_X4 FILLER_30_1888 ();
 FILLCELL_X2 FILLER_30_1892 ();
 FILLCELL_X32 FILLER_30_1895 ();
 FILLCELL_X32 FILLER_30_1927 ();
 FILLCELL_X32 FILLER_30_1959 ();
 FILLCELL_X32 FILLER_30_1991 ();
 FILLCELL_X32 FILLER_30_2023 ();
 FILLCELL_X32 FILLER_30_2055 ();
 FILLCELL_X32 FILLER_30_2087 ();
 FILLCELL_X32 FILLER_30_2119 ();
 FILLCELL_X32 FILLER_30_2151 ();
 FILLCELL_X32 FILLER_30_2183 ();
 FILLCELL_X32 FILLER_30_2215 ();
 FILLCELL_X32 FILLER_30_2247 ();
 FILLCELL_X32 FILLER_30_2279 ();
 FILLCELL_X32 FILLER_30_2311 ();
 FILLCELL_X32 FILLER_30_2343 ();
 FILLCELL_X32 FILLER_30_2375 ();
 FILLCELL_X16 FILLER_30_2407 ();
 FILLCELL_X8 FILLER_30_2423 ();
 FILLCELL_X4 FILLER_30_2431 ();
 FILLCELL_X1 FILLER_30_2435 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X32 FILLER_31_1776 ();
 FILLCELL_X32 FILLER_31_1808 ();
 FILLCELL_X32 FILLER_31_1840 ();
 FILLCELL_X32 FILLER_31_1872 ();
 FILLCELL_X32 FILLER_31_1904 ();
 FILLCELL_X32 FILLER_31_1936 ();
 FILLCELL_X32 FILLER_31_1968 ();
 FILLCELL_X32 FILLER_31_2000 ();
 FILLCELL_X32 FILLER_31_2032 ();
 FILLCELL_X32 FILLER_31_2064 ();
 FILLCELL_X32 FILLER_31_2096 ();
 FILLCELL_X32 FILLER_31_2128 ();
 FILLCELL_X32 FILLER_31_2160 ();
 FILLCELL_X32 FILLER_31_2192 ();
 FILLCELL_X32 FILLER_31_2224 ();
 FILLCELL_X32 FILLER_31_2256 ();
 FILLCELL_X32 FILLER_31_2288 ();
 FILLCELL_X32 FILLER_31_2320 ();
 FILLCELL_X32 FILLER_31_2352 ();
 FILLCELL_X32 FILLER_31_2384 ();
 FILLCELL_X16 FILLER_31_2416 ();
 FILLCELL_X4 FILLER_31_2432 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X32 FILLER_32_1784 ();
 FILLCELL_X32 FILLER_32_1816 ();
 FILLCELL_X32 FILLER_32_1848 ();
 FILLCELL_X8 FILLER_32_1880 ();
 FILLCELL_X4 FILLER_32_1888 ();
 FILLCELL_X2 FILLER_32_1892 ();
 FILLCELL_X32 FILLER_32_1895 ();
 FILLCELL_X32 FILLER_32_1927 ();
 FILLCELL_X32 FILLER_32_1959 ();
 FILLCELL_X32 FILLER_32_1991 ();
 FILLCELL_X32 FILLER_32_2023 ();
 FILLCELL_X32 FILLER_32_2055 ();
 FILLCELL_X32 FILLER_32_2087 ();
 FILLCELL_X32 FILLER_32_2119 ();
 FILLCELL_X32 FILLER_32_2151 ();
 FILLCELL_X32 FILLER_32_2183 ();
 FILLCELL_X32 FILLER_32_2215 ();
 FILLCELL_X32 FILLER_32_2247 ();
 FILLCELL_X32 FILLER_32_2279 ();
 FILLCELL_X32 FILLER_32_2311 ();
 FILLCELL_X32 FILLER_32_2343 ();
 FILLCELL_X32 FILLER_32_2375 ();
 FILLCELL_X16 FILLER_32_2407 ();
 FILLCELL_X8 FILLER_32_2423 ();
 FILLCELL_X4 FILLER_32_2431 ();
 FILLCELL_X1 FILLER_32_2435 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X32 FILLER_33_1776 ();
 FILLCELL_X32 FILLER_33_1808 ();
 FILLCELL_X32 FILLER_33_1840 ();
 FILLCELL_X32 FILLER_33_1872 ();
 FILLCELL_X32 FILLER_33_1904 ();
 FILLCELL_X32 FILLER_33_1936 ();
 FILLCELL_X32 FILLER_33_1968 ();
 FILLCELL_X32 FILLER_33_2000 ();
 FILLCELL_X32 FILLER_33_2032 ();
 FILLCELL_X32 FILLER_33_2064 ();
 FILLCELL_X32 FILLER_33_2096 ();
 FILLCELL_X32 FILLER_33_2128 ();
 FILLCELL_X32 FILLER_33_2160 ();
 FILLCELL_X32 FILLER_33_2192 ();
 FILLCELL_X32 FILLER_33_2224 ();
 FILLCELL_X32 FILLER_33_2256 ();
 FILLCELL_X32 FILLER_33_2288 ();
 FILLCELL_X32 FILLER_33_2320 ();
 FILLCELL_X32 FILLER_33_2352 ();
 FILLCELL_X32 FILLER_33_2384 ();
 FILLCELL_X16 FILLER_33_2416 ();
 FILLCELL_X4 FILLER_33_2432 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X32 FILLER_34_1784 ();
 FILLCELL_X32 FILLER_34_1816 ();
 FILLCELL_X32 FILLER_34_1848 ();
 FILLCELL_X8 FILLER_34_1880 ();
 FILLCELL_X4 FILLER_34_1888 ();
 FILLCELL_X2 FILLER_34_1892 ();
 FILLCELL_X32 FILLER_34_1895 ();
 FILLCELL_X32 FILLER_34_1927 ();
 FILLCELL_X32 FILLER_34_1959 ();
 FILLCELL_X32 FILLER_34_1991 ();
 FILLCELL_X32 FILLER_34_2023 ();
 FILLCELL_X32 FILLER_34_2055 ();
 FILLCELL_X32 FILLER_34_2087 ();
 FILLCELL_X32 FILLER_34_2119 ();
 FILLCELL_X32 FILLER_34_2151 ();
 FILLCELL_X32 FILLER_34_2183 ();
 FILLCELL_X32 FILLER_34_2215 ();
 FILLCELL_X32 FILLER_34_2247 ();
 FILLCELL_X32 FILLER_34_2279 ();
 FILLCELL_X32 FILLER_34_2311 ();
 FILLCELL_X32 FILLER_34_2343 ();
 FILLCELL_X32 FILLER_34_2375 ();
 FILLCELL_X16 FILLER_34_2407 ();
 FILLCELL_X8 FILLER_34_2423 ();
 FILLCELL_X4 FILLER_34_2431 ();
 FILLCELL_X1 FILLER_34_2435 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X32 FILLER_35_1776 ();
 FILLCELL_X32 FILLER_35_1808 ();
 FILLCELL_X32 FILLER_35_1840 ();
 FILLCELL_X32 FILLER_35_1872 ();
 FILLCELL_X32 FILLER_35_1904 ();
 FILLCELL_X32 FILLER_35_1936 ();
 FILLCELL_X32 FILLER_35_1968 ();
 FILLCELL_X32 FILLER_35_2000 ();
 FILLCELL_X32 FILLER_35_2032 ();
 FILLCELL_X32 FILLER_35_2064 ();
 FILLCELL_X32 FILLER_35_2096 ();
 FILLCELL_X32 FILLER_35_2128 ();
 FILLCELL_X32 FILLER_35_2160 ();
 FILLCELL_X32 FILLER_35_2192 ();
 FILLCELL_X32 FILLER_35_2224 ();
 FILLCELL_X32 FILLER_35_2256 ();
 FILLCELL_X32 FILLER_35_2288 ();
 FILLCELL_X32 FILLER_35_2320 ();
 FILLCELL_X32 FILLER_35_2352 ();
 FILLCELL_X32 FILLER_35_2384 ();
 FILLCELL_X16 FILLER_35_2416 ();
 FILLCELL_X4 FILLER_35_2432 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X32 FILLER_36_1784 ();
 FILLCELL_X32 FILLER_36_1816 ();
 FILLCELL_X32 FILLER_36_1848 ();
 FILLCELL_X8 FILLER_36_1880 ();
 FILLCELL_X4 FILLER_36_1888 ();
 FILLCELL_X2 FILLER_36_1892 ();
 FILLCELL_X32 FILLER_36_1895 ();
 FILLCELL_X32 FILLER_36_1927 ();
 FILLCELL_X32 FILLER_36_1959 ();
 FILLCELL_X32 FILLER_36_1991 ();
 FILLCELL_X32 FILLER_36_2023 ();
 FILLCELL_X32 FILLER_36_2055 ();
 FILLCELL_X32 FILLER_36_2087 ();
 FILLCELL_X32 FILLER_36_2119 ();
 FILLCELL_X32 FILLER_36_2151 ();
 FILLCELL_X32 FILLER_36_2183 ();
 FILLCELL_X32 FILLER_36_2215 ();
 FILLCELL_X32 FILLER_36_2247 ();
 FILLCELL_X32 FILLER_36_2279 ();
 FILLCELL_X32 FILLER_36_2311 ();
 FILLCELL_X32 FILLER_36_2343 ();
 FILLCELL_X32 FILLER_36_2375 ();
 FILLCELL_X16 FILLER_36_2407 ();
 FILLCELL_X8 FILLER_36_2423 ();
 FILLCELL_X4 FILLER_36_2431 ();
 FILLCELL_X1 FILLER_36_2435 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X32 FILLER_37_1776 ();
 FILLCELL_X32 FILLER_37_1808 ();
 FILLCELL_X32 FILLER_37_1840 ();
 FILLCELL_X32 FILLER_37_1872 ();
 FILLCELL_X32 FILLER_37_1904 ();
 FILLCELL_X32 FILLER_37_1936 ();
 FILLCELL_X32 FILLER_37_1968 ();
 FILLCELL_X32 FILLER_37_2000 ();
 FILLCELL_X32 FILLER_37_2032 ();
 FILLCELL_X32 FILLER_37_2064 ();
 FILLCELL_X32 FILLER_37_2096 ();
 FILLCELL_X32 FILLER_37_2128 ();
 FILLCELL_X32 FILLER_37_2160 ();
 FILLCELL_X32 FILLER_37_2192 ();
 FILLCELL_X32 FILLER_37_2224 ();
 FILLCELL_X32 FILLER_37_2256 ();
 FILLCELL_X32 FILLER_37_2288 ();
 FILLCELL_X32 FILLER_37_2320 ();
 FILLCELL_X32 FILLER_37_2352 ();
 FILLCELL_X32 FILLER_37_2384 ();
 FILLCELL_X16 FILLER_37_2416 ();
 FILLCELL_X4 FILLER_37_2432 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X32 FILLER_38_1784 ();
 FILLCELL_X32 FILLER_38_1816 ();
 FILLCELL_X32 FILLER_38_1848 ();
 FILLCELL_X8 FILLER_38_1880 ();
 FILLCELL_X4 FILLER_38_1888 ();
 FILLCELL_X2 FILLER_38_1892 ();
 FILLCELL_X32 FILLER_38_1895 ();
 FILLCELL_X32 FILLER_38_1927 ();
 FILLCELL_X32 FILLER_38_1959 ();
 FILLCELL_X32 FILLER_38_1991 ();
 FILLCELL_X32 FILLER_38_2023 ();
 FILLCELL_X32 FILLER_38_2055 ();
 FILLCELL_X32 FILLER_38_2087 ();
 FILLCELL_X32 FILLER_38_2119 ();
 FILLCELL_X32 FILLER_38_2151 ();
 FILLCELL_X32 FILLER_38_2183 ();
 FILLCELL_X32 FILLER_38_2215 ();
 FILLCELL_X32 FILLER_38_2247 ();
 FILLCELL_X32 FILLER_38_2279 ();
 FILLCELL_X32 FILLER_38_2311 ();
 FILLCELL_X32 FILLER_38_2343 ();
 FILLCELL_X32 FILLER_38_2375 ();
 FILLCELL_X16 FILLER_38_2407 ();
 FILLCELL_X8 FILLER_38_2423 ();
 FILLCELL_X4 FILLER_38_2431 ();
 FILLCELL_X1 FILLER_38_2435 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X32 FILLER_39_1776 ();
 FILLCELL_X32 FILLER_39_1808 ();
 FILLCELL_X32 FILLER_39_1840 ();
 FILLCELL_X32 FILLER_39_1872 ();
 FILLCELL_X32 FILLER_39_1904 ();
 FILLCELL_X32 FILLER_39_1936 ();
 FILLCELL_X32 FILLER_39_1968 ();
 FILLCELL_X32 FILLER_39_2000 ();
 FILLCELL_X32 FILLER_39_2032 ();
 FILLCELL_X32 FILLER_39_2064 ();
 FILLCELL_X32 FILLER_39_2096 ();
 FILLCELL_X32 FILLER_39_2128 ();
 FILLCELL_X32 FILLER_39_2160 ();
 FILLCELL_X32 FILLER_39_2192 ();
 FILLCELL_X32 FILLER_39_2224 ();
 FILLCELL_X32 FILLER_39_2256 ();
 FILLCELL_X32 FILLER_39_2288 ();
 FILLCELL_X32 FILLER_39_2320 ();
 FILLCELL_X32 FILLER_39_2352 ();
 FILLCELL_X32 FILLER_39_2384 ();
 FILLCELL_X16 FILLER_39_2416 ();
 FILLCELL_X4 FILLER_39_2432 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X32 FILLER_40_1784 ();
 FILLCELL_X32 FILLER_40_1816 ();
 FILLCELL_X32 FILLER_40_1848 ();
 FILLCELL_X8 FILLER_40_1880 ();
 FILLCELL_X4 FILLER_40_1888 ();
 FILLCELL_X2 FILLER_40_1892 ();
 FILLCELL_X32 FILLER_40_1895 ();
 FILLCELL_X32 FILLER_40_1927 ();
 FILLCELL_X32 FILLER_40_1959 ();
 FILLCELL_X32 FILLER_40_1991 ();
 FILLCELL_X32 FILLER_40_2023 ();
 FILLCELL_X32 FILLER_40_2055 ();
 FILLCELL_X32 FILLER_40_2087 ();
 FILLCELL_X32 FILLER_40_2119 ();
 FILLCELL_X32 FILLER_40_2151 ();
 FILLCELL_X32 FILLER_40_2183 ();
 FILLCELL_X32 FILLER_40_2215 ();
 FILLCELL_X32 FILLER_40_2247 ();
 FILLCELL_X32 FILLER_40_2279 ();
 FILLCELL_X32 FILLER_40_2311 ();
 FILLCELL_X32 FILLER_40_2343 ();
 FILLCELL_X32 FILLER_40_2375 ();
 FILLCELL_X16 FILLER_40_2407 ();
 FILLCELL_X8 FILLER_40_2423 ();
 FILLCELL_X4 FILLER_40_2431 ();
 FILLCELL_X1 FILLER_40_2435 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X32 FILLER_41_1776 ();
 FILLCELL_X32 FILLER_41_1808 ();
 FILLCELL_X32 FILLER_41_1840 ();
 FILLCELL_X32 FILLER_41_1872 ();
 FILLCELL_X32 FILLER_41_1904 ();
 FILLCELL_X32 FILLER_41_1936 ();
 FILLCELL_X32 FILLER_41_1968 ();
 FILLCELL_X32 FILLER_41_2000 ();
 FILLCELL_X32 FILLER_41_2032 ();
 FILLCELL_X32 FILLER_41_2064 ();
 FILLCELL_X32 FILLER_41_2096 ();
 FILLCELL_X32 FILLER_41_2128 ();
 FILLCELL_X32 FILLER_41_2160 ();
 FILLCELL_X32 FILLER_41_2192 ();
 FILLCELL_X32 FILLER_41_2224 ();
 FILLCELL_X32 FILLER_41_2256 ();
 FILLCELL_X32 FILLER_41_2288 ();
 FILLCELL_X32 FILLER_41_2320 ();
 FILLCELL_X32 FILLER_41_2352 ();
 FILLCELL_X32 FILLER_41_2384 ();
 FILLCELL_X16 FILLER_41_2416 ();
 FILLCELL_X4 FILLER_41_2432 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X32 FILLER_42_1784 ();
 FILLCELL_X32 FILLER_42_1816 ();
 FILLCELL_X32 FILLER_42_1848 ();
 FILLCELL_X8 FILLER_42_1880 ();
 FILLCELL_X4 FILLER_42_1888 ();
 FILLCELL_X2 FILLER_42_1892 ();
 FILLCELL_X32 FILLER_42_1895 ();
 FILLCELL_X32 FILLER_42_1927 ();
 FILLCELL_X32 FILLER_42_1959 ();
 FILLCELL_X32 FILLER_42_1991 ();
 FILLCELL_X32 FILLER_42_2023 ();
 FILLCELL_X32 FILLER_42_2055 ();
 FILLCELL_X32 FILLER_42_2087 ();
 FILLCELL_X32 FILLER_42_2119 ();
 FILLCELL_X32 FILLER_42_2151 ();
 FILLCELL_X32 FILLER_42_2183 ();
 FILLCELL_X32 FILLER_42_2215 ();
 FILLCELL_X32 FILLER_42_2247 ();
 FILLCELL_X32 FILLER_42_2279 ();
 FILLCELL_X32 FILLER_42_2311 ();
 FILLCELL_X32 FILLER_42_2343 ();
 FILLCELL_X32 FILLER_42_2375 ();
 FILLCELL_X16 FILLER_42_2407 ();
 FILLCELL_X8 FILLER_42_2423 ();
 FILLCELL_X4 FILLER_42_2431 ();
 FILLCELL_X1 FILLER_42_2435 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X32 FILLER_43_1776 ();
 FILLCELL_X32 FILLER_43_1808 ();
 FILLCELL_X32 FILLER_43_1840 ();
 FILLCELL_X32 FILLER_43_1872 ();
 FILLCELL_X32 FILLER_43_1904 ();
 FILLCELL_X32 FILLER_43_1936 ();
 FILLCELL_X32 FILLER_43_1968 ();
 FILLCELL_X32 FILLER_43_2000 ();
 FILLCELL_X32 FILLER_43_2032 ();
 FILLCELL_X32 FILLER_43_2064 ();
 FILLCELL_X32 FILLER_43_2096 ();
 FILLCELL_X32 FILLER_43_2128 ();
 FILLCELL_X32 FILLER_43_2160 ();
 FILLCELL_X32 FILLER_43_2192 ();
 FILLCELL_X32 FILLER_43_2224 ();
 FILLCELL_X32 FILLER_43_2256 ();
 FILLCELL_X32 FILLER_43_2288 ();
 FILLCELL_X32 FILLER_43_2320 ();
 FILLCELL_X32 FILLER_43_2352 ();
 FILLCELL_X32 FILLER_43_2384 ();
 FILLCELL_X16 FILLER_43_2416 ();
 FILLCELL_X4 FILLER_43_2432 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X32 FILLER_44_1784 ();
 FILLCELL_X32 FILLER_44_1816 ();
 FILLCELL_X32 FILLER_44_1848 ();
 FILLCELL_X8 FILLER_44_1880 ();
 FILLCELL_X4 FILLER_44_1888 ();
 FILLCELL_X2 FILLER_44_1892 ();
 FILLCELL_X32 FILLER_44_1895 ();
 FILLCELL_X32 FILLER_44_1927 ();
 FILLCELL_X32 FILLER_44_1959 ();
 FILLCELL_X32 FILLER_44_1991 ();
 FILLCELL_X32 FILLER_44_2023 ();
 FILLCELL_X32 FILLER_44_2055 ();
 FILLCELL_X32 FILLER_44_2087 ();
 FILLCELL_X32 FILLER_44_2119 ();
 FILLCELL_X32 FILLER_44_2151 ();
 FILLCELL_X32 FILLER_44_2183 ();
 FILLCELL_X32 FILLER_44_2215 ();
 FILLCELL_X32 FILLER_44_2247 ();
 FILLCELL_X32 FILLER_44_2279 ();
 FILLCELL_X32 FILLER_44_2311 ();
 FILLCELL_X32 FILLER_44_2343 ();
 FILLCELL_X32 FILLER_44_2375 ();
 FILLCELL_X16 FILLER_44_2407 ();
 FILLCELL_X8 FILLER_44_2423 ();
 FILLCELL_X4 FILLER_44_2431 ();
 FILLCELL_X1 FILLER_44_2435 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X32 FILLER_45_1776 ();
 FILLCELL_X32 FILLER_45_1808 ();
 FILLCELL_X32 FILLER_45_1840 ();
 FILLCELL_X32 FILLER_45_1872 ();
 FILLCELL_X32 FILLER_45_1904 ();
 FILLCELL_X32 FILLER_45_1936 ();
 FILLCELL_X32 FILLER_45_1968 ();
 FILLCELL_X32 FILLER_45_2000 ();
 FILLCELL_X32 FILLER_45_2032 ();
 FILLCELL_X32 FILLER_45_2064 ();
 FILLCELL_X32 FILLER_45_2096 ();
 FILLCELL_X32 FILLER_45_2128 ();
 FILLCELL_X32 FILLER_45_2160 ();
 FILLCELL_X32 FILLER_45_2192 ();
 FILLCELL_X32 FILLER_45_2224 ();
 FILLCELL_X32 FILLER_45_2256 ();
 FILLCELL_X32 FILLER_45_2288 ();
 FILLCELL_X32 FILLER_45_2320 ();
 FILLCELL_X32 FILLER_45_2352 ();
 FILLCELL_X32 FILLER_45_2384 ();
 FILLCELL_X16 FILLER_45_2416 ();
 FILLCELL_X4 FILLER_45_2432 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X32 FILLER_46_1784 ();
 FILLCELL_X32 FILLER_46_1816 ();
 FILLCELL_X32 FILLER_46_1848 ();
 FILLCELL_X8 FILLER_46_1880 ();
 FILLCELL_X4 FILLER_46_1888 ();
 FILLCELL_X2 FILLER_46_1892 ();
 FILLCELL_X32 FILLER_46_1895 ();
 FILLCELL_X32 FILLER_46_1927 ();
 FILLCELL_X32 FILLER_46_1959 ();
 FILLCELL_X32 FILLER_46_1991 ();
 FILLCELL_X32 FILLER_46_2023 ();
 FILLCELL_X32 FILLER_46_2055 ();
 FILLCELL_X32 FILLER_46_2087 ();
 FILLCELL_X32 FILLER_46_2119 ();
 FILLCELL_X32 FILLER_46_2151 ();
 FILLCELL_X32 FILLER_46_2183 ();
 FILLCELL_X32 FILLER_46_2215 ();
 FILLCELL_X32 FILLER_46_2247 ();
 FILLCELL_X32 FILLER_46_2279 ();
 FILLCELL_X32 FILLER_46_2311 ();
 FILLCELL_X32 FILLER_46_2343 ();
 FILLCELL_X32 FILLER_46_2375 ();
 FILLCELL_X16 FILLER_46_2407 ();
 FILLCELL_X8 FILLER_46_2423 ();
 FILLCELL_X4 FILLER_46_2431 ();
 FILLCELL_X1 FILLER_46_2435 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X32 FILLER_47_1776 ();
 FILLCELL_X32 FILLER_47_1808 ();
 FILLCELL_X32 FILLER_47_1840 ();
 FILLCELL_X32 FILLER_47_1872 ();
 FILLCELL_X32 FILLER_47_1904 ();
 FILLCELL_X32 FILLER_47_1936 ();
 FILLCELL_X32 FILLER_47_1968 ();
 FILLCELL_X32 FILLER_47_2000 ();
 FILLCELL_X32 FILLER_47_2032 ();
 FILLCELL_X32 FILLER_47_2064 ();
 FILLCELL_X32 FILLER_47_2096 ();
 FILLCELL_X32 FILLER_47_2128 ();
 FILLCELL_X32 FILLER_47_2160 ();
 FILLCELL_X32 FILLER_47_2192 ();
 FILLCELL_X32 FILLER_47_2224 ();
 FILLCELL_X32 FILLER_47_2256 ();
 FILLCELL_X32 FILLER_47_2288 ();
 FILLCELL_X32 FILLER_47_2320 ();
 FILLCELL_X32 FILLER_47_2352 ();
 FILLCELL_X32 FILLER_47_2384 ();
 FILLCELL_X16 FILLER_47_2416 ();
 FILLCELL_X4 FILLER_47_2432 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X32 FILLER_48_1784 ();
 FILLCELL_X32 FILLER_48_1816 ();
 FILLCELL_X32 FILLER_48_1848 ();
 FILLCELL_X8 FILLER_48_1880 ();
 FILLCELL_X4 FILLER_48_1888 ();
 FILLCELL_X2 FILLER_48_1892 ();
 FILLCELL_X32 FILLER_48_1895 ();
 FILLCELL_X32 FILLER_48_1927 ();
 FILLCELL_X32 FILLER_48_1959 ();
 FILLCELL_X32 FILLER_48_1991 ();
 FILLCELL_X32 FILLER_48_2023 ();
 FILLCELL_X32 FILLER_48_2055 ();
 FILLCELL_X32 FILLER_48_2087 ();
 FILLCELL_X32 FILLER_48_2119 ();
 FILLCELL_X32 FILLER_48_2151 ();
 FILLCELL_X32 FILLER_48_2183 ();
 FILLCELL_X32 FILLER_48_2215 ();
 FILLCELL_X32 FILLER_48_2247 ();
 FILLCELL_X32 FILLER_48_2279 ();
 FILLCELL_X32 FILLER_48_2311 ();
 FILLCELL_X32 FILLER_48_2343 ();
 FILLCELL_X32 FILLER_48_2375 ();
 FILLCELL_X16 FILLER_48_2407 ();
 FILLCELL_X8 FILLER_48_2423 ();
 FILLCELL_X4 FILLER_48_2431 ();
 FILLCELL_X1 FILLER_48_2435 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X32 FILLER_49_1776 ();
 FILLCELL_X32 FILLER_49_1808 ();
 FILLCELL_X32 FILLER_49_1840 ();
 FILLCELL_X32 FILLER_49_1872 ();
 FILLCELL_X32 FILLER_49_1904 ();
 FILLCELL_X32 FILLER_49_1936 ();
 FILLCELL_X32 FILLER_49_1968 ();
 FILLCELL_X32 FILLER_49_2000 ();
 FILLCELL_X32 FILLER_49_2032 ();
 FILLCELL_X32 FILLER_49_2064 ();
 FILLCELL_X32 FILLER_49_2096 ();
 FILLCELL_X32 FILLER_49_2128 ();
 FILLCELL_X32 FILLER_49_2160 ();
 FILLCELL_X32 FILLER_49_2192 ();
 FILLCELL_X32 FILLER_49_2224 ();
 FILLCELL_X32 FILLER_49_2256 ();
 FILLCELL_X32 FILLER_49_2288 ();
 FILLCELL_X32 FILLER_49_2320 ();
 FILLCELL_X32 FILLER_49_2352 ();
 FILLCELL_X32 FILLER_49_2384 ();
 FILLCELL_X16 FILLER_49_2416 ();
 FILLCELL_X4 FILLER_49_2432 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X32 FILLER_50_1784 ();
 FILLCELL_X32 FILLER_50_1816 ();
 FILLCELL_X32 FILLER_50_1848 ();
 FILLCELL_X8 FILLER_50_1880 ();
 FILLCELL_X4 FILLER_50_1888 ();
 FILLCELL_X2 FILLER_50_1892 ();
 FILLCELL_X32 FILLER_50_1895 ();
 FILLCELL_X32 FILLER_50_1927 ();
 FILLCELL_X32 FILLER_50_1959 ();
 FILLCELL_X32 FILLER_50_1991 ();
 FILLCELL_X32 FILLER_50_2023 ();
 FILLCELL_X32 FILLER_50_2055 ();
 FILLCELL_X32 FILLER_50_2087 ();
 FILLCELL_X32 FILLER_50_2119 ();
 FILLCELL_X32 FILLER_50_2151 ();
 FILLCELL_X32 FILLER_50_2183 ();
 FILLCELL_X32 FILLER_50_2215 ();
 FILLCELL_X32 FILLER_50_2247 ();
 FILLCELL_X32 FILLER_50_2279 ();
 FILLCELL_X32 FILLER_50_2311 ();
 FILLCELL_X32 FILLER_50_2343 ();
 FILLCELL_X32 FILLER_50_2375 ();
 FILLCELL_X16 FILLER_50_2407 ();
 FILLCELL_X8 FILLER_50_2423 ();
 FILLCELL_X4 FILLER_50_2431 ();
 FILLCELL_X1 FILLER_50_2435 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X32 FILLER_51_1776 ();
 FILLCELL_X32 FILLER_51_1808 ();
 FILLCELL_X32 FILLER_51_1840 ();
 FILLCELL_X32 FILLER_51_1872 ();
 FILLCELL_X32 FILLER_51_1904 ();
 FILLCELL_X32 FILLER_51_1936 ();
 FILLCELL_X32 FILLER_51_1968 ();
 FILLCELL_X32 FILLER_51_2000 ();
 FILLCELL_X32 FILLER_51_2032 ();
 FILLCELL_X32 FILLER_51_2064 ();
 FILLCELL_X32 FILLER_51_2096 ();
 FILLCELL_X32 FILLER_51_2128 ();
 FILLCELL_X32 FILLER_51_2160 ();
 FILLCELL_X32 FILLER_51_2192 ();
 FILLCELL_X32 FILLER_51_2224 ();
 FILLCELL_X32 FILLER_51_2256 ();
 FILLCELL_X32 FILLER_51_2288 ();
 FILLCELL_X32 FILLER_51_2320 ();
 FILLCELL_X32 FILLER_51_2352 ();
 FILLCELL_X32 FILLER_51_2384 ();
 FILLCELL_X16 FILLER_51_2416 ();
 FILLCELL_X4 FILLER_51_2432 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X32 FILLER_52_1784 ();
 FILLCELL_X32 FILLER_52_1816 ();
 FILLCELL_X32 FILLER_52_1848 ();
 FILLCELL_X8 FILLER_52_1880 ();
 FILLCELL_X4 FILLER_52_1888 ();
 FILLCELL_X2 FILLER_52_1892 ();
 FILLCELL_X32 FILLER_52_1895 ();
 FILLCELL_X32 FILLER_52_1927 ();
 FILLCELL_X32 FILLER_52_1959 ();
 FILLCELL_X32 FILLER_52_1991 ();
 FILLCELL_X32 FILLER_52_2023 ();
 FILLCELL_X32 FILLER_52_2055 ();
 FILLCELL_X32 FILLER_52_2087 ();
 FILLCELL_X32 FILLER_52_2119 ();
 FILLCELL_X32 FILLER_52_2151 ();
 FILLCELL_X32 FILLER_52_2183 ();
 FILLCELL_X32 FILLER_52_2215 ();
 FILLCELL_X32 FILLER_52_2247 ();
 FILLCELL_X32 FILLER_52_2279 ();
 FILLCELL_X32 FILLER_52_2311 ();
 FILLCELL_X32 FILLER_52_2343 ();
 FILLCELL_X32 FILLER_52_2375 ();
 FILLCELL_X16 FILLER_52_2407 ();
 FILLCELL_X8 FILLER_52_2423 ();
 FILLCELL_X4 FILLER_52_2431 ();
 FILLCELL_X1 FILLER_52_2435 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X32 FILLER_53_1776 ();
 FILLCELL_X32 FILLER_53_1808 ();
 FILLCELL_X32 FILLER_53_1840 ();
 FILLCELL_X32 FILLER_53_1872 ();
 FILLCELL_X32 FILLER_53_1904 ();
 FILLCELL_X32 FILLER_53_1936 ();
 FILLCELL_X32 FILLER_53_1968 ();
 FILLCELL_X32 FILLER_53_2000 ();
 FILLCELL_X32 FILLER_53_2032 ();
 FILLCELL_X32 FILLER_53_2064 ();
 FILLCELL_X32 FILLER_53_2096 ();
 FILLCELL_X32 FILLER_53_2128 ();
 FILLCELL_X32 FILLER_53_2160 ();
 FILLCELL_X32 FILLER_53_2192 ();
 FILLCELL_X32 FILLER_53_2224 ();
 FILLCELL_X32 FILLER_53_2256 ();
 FILLCELL_X32 FILLER_53_2288 ();
 FILLCELL_X32 FILLER_53_2320 ();
 FILLCELL_X32 FILLER_53_2352 ();
 FILLCELL_X32 FILLER_53_2384 ();
 FILLCELL_X16 FILLER_53_2416 ();
 FILLCELL_X4 FILLER_53_2432 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X32 FILLER_54_1784 ();
 FILLCELL_X32 FILLER_54_1816 ();
 FILLCELL_X32 FILLER_54_1848 ();
 FILLCELL_X8 FILLER_54_1880 ();
 FILLCELL_X4 FILLER_54_1888 ();
 FILLCELL_X2 FILLER_54_1892 ();
 FILLCELL_X32 FILLER_54_1895 ();
 FILLCELL_X32 FILLER_54_1927 ();
 FILLCELL_X32 FILLER_54_1959 ();
 FILLCELL_X32 FILLER_54_1991 ();
 FILLCELL_X32 FILLER_54_2023 ();
 FILLCELL_X32 FILLER_54_2055 ();
 FILLCELL_X32 FILLER_54_2087 ();
 FILLCELL_X32 FILLER_54_2119 ();
 FILLCELL_X32 FILLER_54_2151 ();
 FILLCELL_X32 FILLER_54_2183 ();
 FILLCELL_X32 FILLER_54_2215 ();
 FILLCELL_X32 FILLER_54_2247 ();
 FILLCELL_X32 FILLER_54_2279 ();
 FILLCELL_X32 FILLER_54_2311 ();
 FILLCELL_X32 FILLER_54_2343 ();
 FILLCELL_X32 FILLER_54_2375 ();
 FILLCELL_X16 FILLER_54_2407 ();
 FILLCELL_X8 FILLER_54_2423 ();
 FILLCELL_X4 FILLER_54_2431 ();
 FILLCELL_X1 FILLER_54_2435 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X32 FILLER_55_1776 ();
 FILLCELL_X32 FILLER_55_1808 ();
 FILLCELL_X32 FILLER_55_1840 ();
 FILLCELL_X32 FILLER_55_1872 ();
 FILLCELL_X32 FILLER_55_1904 ();
 FILLCELL_X32 FILLER_55_1936 ();
 FILLCELL_X32 FILLER_55_1968 ();
 FILLCELL_X32 FILLER_55_2000 ();
 FILLCELL_X32 FILLER_55_2032 ();
 FILLCELL_X32 FILLER_55_2064 ();
 FILLCELL_X32 FILLER_55_2096 ();
 FILLCELL_X32 FILLER_55_2128 ();
 FILLCELL_X32 FILLER_55_2160 ();
 FILLCELL_X32 FILLER_55_2192 ();
 FILLCELL_X32 FILLER_55_2224 ();
 FILLCELL_X32 FILLER_55_2256 ();
 FILLCELL_X32 FILLER_55_2288 ();
 FILLCELL_X32 FILLER_55_2320 ();
 FILLCELL_X32 FILLER_55_2352 ();
 FILLCELL_X32 FILLER_55_2384 ();
 FILLCELL_X16 FILLER_55_2416 ();
 FILLCELL_X4 FILLER_55_2432 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X32 FILLER_56_1784 ();
 FILLCELL_X32 FILLER_56_1816 ();
 FILLCELL_X32 FILLER_56_1848 ();
 FILLCELL_X8 FILLER_56_1880 ();
 FILLCELL_X4 FILLER_56_1888 ();
 FILLCELL_X2 FILLER_56_1892 ();
 FILLCELL_X32 FILLER_56_1895 ();
 FILLCELL_X32 FILLER_56_1927 ();
 FILLCELL_X32 FILLER_56_1959 ();
 FILLCELL_X32 FILLER_56_1991 ();
 FILLCELL_X32 FILLER_56_2023 ();
 FILLCELL_X32 FILLER_56_2055 ();
 FILLCELL_X32 FILLER_56_2087 ();
 FILLCELL_X32 FILLER_56_2119 ();
 FILLCELL_X32 FILLER_56_2151 ();
 FILLCELL_X32 FILLER_56_2183 ();
 FILLCELL_X32 FILLER_56_2215 ();
 FILLCELL_X32 FILLER_56_2247 ();
 FILLCELL_X32 FILLER_56_2279 ();
 FILLCELL_X32 FILLER_56_2311 ();
 FILLCELL_X32 FILLER_56_2343 ();
 FILLCELL_X32 FILLER_56_2375 ();
 FILLCELL_X16 FILLER_56_2407 ();
 FILLCELL_X8 FILLER_56_2423 ();
 FILLCELL_X4 FILLER_56_2431 ();
 FILLCELL_X1 FILLER_56_2435 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X32 FILLER_57_1776 ();
 FILLCELL_X32 FILLER_57_1808 ();
 FILLCELL_X32 FILLER_57_1840 ();
 FILLCELL_X32 FILLER_57_1872 ();
 FILLCELL_X32 FILLER_57_1904 ();
 FILLCELL_X32 FILLER_57_1936 ();
 FILLCELL_X32 FILLER_57_1968 ();
 FILLCELL_X32 FILLER_57_2000 ();
 FILLCELL_X32 FILLER_57_2032 ();
 FILLCELL_X32 FILLER_57_2064 ();
 FILLCELL_X32 FILLER_57_2096 ();
 FILLCELL_X32 FILLER_57_2128 ();
 FILLCELL_X32 FILLER_57_2160 ();
 FILLCELL_X32 FILLER_57_2192 ();
 FILLCELL_X32 FILLER_57_2224 ();
 FILLCELL_X32 FILLER_57_2256 ();
 FILLCELL_X32 FILLER_57_2288 ();
 FILLCELL_X32 FILLER_57_2320 ();
 FILLCELL_X32 FILLER_57_2352 ();
 FILLCELL_X32 FILLER_57_2384 ();
 FILLCELL_X16 FILLER_57_2416 ();
 FILLCELL_X4 FILLER_57_2432 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X32 FILLER_58_1784 ();
 FILLCELL_X32 FILLER_58_1816 ();
 FILLCELL_X32 FILLER_58_1848 ();
 FILLCELL_X8 FILLER_58_1880 ();
 FILLCELL_X4 FILLER_58_1888 ();
 FILLCELL_X2 FILLER_58_1892 ();
 FILLCELL_X32 FILLER_58_1895 ();
 FILLCELL_X32 FILLER_58_1927 ();
 FILLCELL_X32 FILLER_58_1959 ();
 FILLCELL_X32 FILLER_58_1991 ();
 FILLCELL_X32 FILLER_58_2023 ();
 FILLCELL_X32 FILLER_58_2055 ();
 FILLCELL_X32 FILLER_58_2087 ();
 FILLCELL_X32 FILLER_58_2119 ();
 FILLCELL_X32 FILLER_58_2151 ();
 FILLCELL_X32 FILLER_58_2183 ();
 FILLCELL_X32 FILLER_58_2215 ();
 FILLCELL_X32 FILLER_58_2247 ();
 FILLCELL_X32 FILLER_58_2279 ();
 FILLCELL_X32 FILLER_58_2311 ();
 FILLCELL_X32 FILLER_58_2343 ();
 FILLCELL_X32 FILLER_58_2375 ();
 FILLCELL_X16 FILLER_58_2407 ();
 FILLCELL_X8 FILLER_58_2423 ();
 FILLCELL_X4 FILLER_58_2431 ();
 FILLCELL_X1 FILLER_58_2435 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X32 FILLER_59_1776 ();
 FILLCELL_X32 FILLER_59_1808 ();
 FILLCELL_X32 FILLER_59_1840 ();
 FILLCELL_X32 FILLER_59_1872 ();
 FILLCELL_X32 FILLER_59_1904 ();
 FILLCELL_X32 FILLER_59_1936 ();
 FILLCELL_X32 FILLER_59_1968 ();
 FILLCELL_X32 FILLER_59_2000 ();
 FILLCELL_X32 FILLER_59_2032 ();
 FILLCELL_X32 FILLER_59_2064 ();
 FILLCELL_X32 FILLER_59_2096 ();
 FILLCELL_X32 FILLER_59_2128 ();
 FILLCELL_X32 FILLER_59_2160 ();
 FILLCELL_X32 FILLER_59_2192 ();
 FILLCELL_X32 FILLER_59_2224 ();
 FILLCELL_X32 FILLER_59_2256 ();
 FILLCELL_X32 FILLER_59_2288 ();
 FILLCELL_X32 FILLER_59_2320 ();
 FILLCELL_X32 FILLER_59_2352 ();
 FILLCELL_X32 FILLER_59_2384 ();
 FILLCELL_X16 FILLER_59_2416 ();
 FILLCELL_X4 FILLER_59_2432 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X32 FILLER_60_1784 ();
 FILLCELL_X32 FILLER_60_1816 ();
 FILLCELL_X32 FILLER_60_1848 ();
 FILLCELL_X8 FILLER_60_1880 ();
 FILLCELL_X4 FILLER_60_1888 ();
 FILLCELL_X2 FILLER_60_1892 ();
 FILLCELL_X32 FILLER_60_1895 ();
 FILLCELL_X32 FILLER_60_1927 ();
 FILLCELL_X32 FILLER_60_1959 ();
 FILLCELL_X32 FILLER_60_1991 ();
 FILLCELL_X32 FILLER_60_2023 ();
 FILLCELL_X32 FILLER_60_2055 ();
 FILLCELL_X32 FILLER_60_2087 ();
 FILLCELL_X32 FILLER_60_2119 ();
 FILLCELL_X32 FILLER_60_2151 ();
 FILLCELL_X32 FILLER_60_2183 ();
 FILLCELL_X32 FILLER_60_2215 ();
 FILLCELL_X32 FILLER_60_2247 ();
 FILLCELL_X32 FILLER_60_2279 ();
 FILLCELL_X32 FILLER_60_2311 ();
 FILLCELL_X32 FILLER_60_2343 ();
 FILLCELL_X32 FILLER_60_2375 ();
 FILLCELL_X16 FILLER_60_2407 ();
 FILLCELL_X8 FILLER_60_2423 ();
 FILLCELL_X4 FILLER_60_2431 ();
 FILLCELL_X1 FILLER_60_2435 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X32 FILLER_61_1776 ();
 FILLCELL_X32 FILLER_61_1808 ();
 FILLCELL_X32 FILLER_61_1840 ();
 FILLCELL_X32 FILLER_61_1872 ();
 FILLCELL_X32 FILLER_61_1904 ();
 FILLCELL_X32 FILLER_61_1936 ();
 FILLCELL_X32 FILLER_61_1968 ();
 FILLCELL_X32 FILLER_61_2000 ();
 FILLCELL_X32 FILLER_61_2032 ();
 FILLCELL_X32 FILLER_61_2064 ();
 FILLCELL_X32 FILLER_61_2096 ();
 FILLCELL_X32 FILLER_61_2128 ();
 FILLCELL_X32 FILLER_61_2160 ();
 FILLCELL_X32 FILLER_61_2192 ();
 FILLCELL_X32 FILLER_61_2224 ();
 FILLCELL_X32 FILLER_61_2256 ();
 FILLCELL_X32 FILLER_61_2288 ();
 FILLCELL_X32 FILLER_61_2320 ();
 FILLCELL_X32 FILLER_61_2352 ();
 FILLCELL_X32 FILLER_61_2384 ();
 FILLCELL_X16 FILLER_61_2416 ();
 FILLCELL_X4 FILLER_61_2432 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X32 FILLER_62_1784 ();
 FILLCELL_X32 FILLER_62_1816 ();
 FILLCELL_X32 FILLER_62_1848 ();
 FILLCELL_X8 FILLER_62_1880 ();
 FILLCELL_X4 FILLER_62_1888 ();
 FILLCELL_X2 FILLER_62_1892 ();
 FILLCELL_X32 FILLER_62_1895 ();
 FILLCELL_X32 FILLER_62_1927 ();
 FILLCELL_X32 FILLER_62_1959 ();
 FILLCELL_X32 FILLER_62_1991 ();
 FILLCELL_X32 FILLER_62_2023 ();
 FILLCELL_X32 FILLER_62_2055 ();
 FILLCELL_X32 FILLER_62_2087 ();
 FILLCELL_X32 FILLER_62_2119 ();
 FILLCELL_X32 FILLER_62_2151 ();
 FILLCELL_X32 FILLER_62_2183 ();
 FILLCELL_X32 FILLER_62_2215 ();
 FILLCELL_X32 FILLER_62_2247 ();
 FILLCELL_X32 FILLER_62_2279 ();
 FILLCELL_X32 FILLER_62_2311 ();
 FILLCELL_X32 FILLER_62_2343 ();
 FILLCELL_X32 FILLER_62_2375 ();
 FILLCELL_X16 FILLER_62_2407 ();
 FILLCELL_X8 FILLER_62_2423 ();
 FILLCELL_X4 FILLER_62_2431 ();
 FILLCELL_X1 FILLER_62_2435 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X32 FILLER_63_1776 ();
 FILLCELL_X32 FILLER_63_1808 ();
 FILLCELL_X32 FILLER_63_1840 ();
 FILLCELL_X32 FILLER_63_1872 ();
 FILLCELL_X32 FILLER_63_1904 ();
 FILLCELL_X32 FILLER_63_1936 ();
 FILLCELL_X32 FILLER_63_1968 ();
 FILLCELL_X32 FILLER_63_2000 ();
 FILLCELL_X32 FILLER_63_2032 ();
 FILLCELL_X32 FILLER_63_2064 ();
 FILLCELL_X32 FILLER_63_2096 ();
 FILLCELL_X32 FILLER_63_2128 ();
 FILLCELL_X32 FILLER_63_2160 ();
 FILLCELL_X32 FILLER_63_2192 ();
 FILLCELL_X32 FILLER_63_2224 ();
 FILLCELL_X32 FILLER_63_2256 ();
 FILLCELL_X32 FILLER_63_2288 ();
 FILLCELL_X32 FILLER_63_2320 ();
 FILLCELL_X32 FILLER_63_2352 ();
 FILLCELL_X32 FILLER_63_2384 ();
 FILLCELL_X16 FILLER_63_2416 ();
 FILLCELL_X4 FILLER_63_2432 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X32 FILLER_64_1784 ();
 FILLCELL_X32 FILLER_64_1816 ();
 FILLCELL_X32 FILLER_64_1848 ();
 FILLCELL_X8 FILLER_64_1880 ();
 FILLCELL_X4 FILLER_64_1888 ();
 FILLCELL_X2 FILLER_64_1892 ();
 FILLCELL_X32 FILLER_64_1895 ();
 FILLCELL_X32 FILLER_64_1927 ();
 FILLCELL_X32 FILLER_64_1959 ();
 FILLCELL_X32 FILLER_64_1991 ();
 FILLCELL_X32 FILLER_64_2023 ();
 FILLCELL_X32 FILLER_64_2055 ();
 FILLCELL_X32 FILLER_64_2087 ();
 FILLCELL_X32 FILLER_64_2119 ();
 FILLCELL_X32 FILLER_64_2151 ();
 FILLCELL_X32 FILLER_64_2183 ();
 FILLCELL_X32 FILLER_64_2215 ();
 FILLCELL_X32 FILLER_64_2247 ();
 FILLCELL_X32 FILLER_64_2279 ();
 FILLCELL_X32 FILLER_64_2311 ();
 FILLCELL_X32 FILLER_64_2343 ();
 FILLCELL_X32 FILLER_64_2375 ();
 FILLCELL_X16 FILLER_64_2407 ();
 FILLCELL_X8 FILLER_64_2423 ();
 FILLCELL_X4 FILLER_64_2431 ();
 FILLCELL_X1 FILLER_64_2435 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X32 FILLER_65_1776 ();
 FILLCELL_X32 FILLER_65_1808 ();
 FILLCELL_X32 FILLER_65_1840 ();
 FILLCELL_X32 FILLER_65_1872 ();
 FILLCELL_X32 FILLER_65_1904 ();
 FILLCELL_X32 FILLER_65_1936 ();
 FILLCELL_X32 FILLER_65_1968 ();
 FILLCELL_X32 FILLER_65_2000 ();
 FILLCELL_X32 FILLER_65_2032 ();
 FILLCELL_X32 FILLER_65_2064 ();
 FILLCELL_X32 FILLER_65_2096 ();
 FILLCELL_X32 FILLER_65_2128 ();
 FILLCELL_X32 FILLER_65_2160 ();
 FILLCELL_X32 FILLER_65_2192 ();
 FILLCELL_X32 FILLER_65_2224 ();
 FILLCELL_X32 FILLER_65_2256 ();
 FILLCELL_X32 FILLER_65_2288 ();
 FILLCELL_X32 FILLER_65_2320 ();
 FILLCELL_X32 FILLER_65_2352 ();
 FILLCELL_X32 FILLER_65_2384 ();
 FILLCELL_X16 FILLER_65_2416 ();
 FILLCELL_X4 FILLER_65_2432 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X32 FILLER_66_1784 ();
 FILLCELL_X32 FILLER_66_1816 ();
 FILLCELL_X32 FILLER_66_1848 ();
 FILLCELL_X8 FILLER_66_1880 ();
 FILLCELL_X4 FILLER_66_1888 ();
 FILLCELL_X2 FILLER_66_1892 ();
 FILLCELL_X32 FILLER_66_1895 ();
 FILLCELL_X32 FILLER_66_1927 ();
 FILLCELL_X32 FILLER_66_1959 ();
 FILLCELL_X32 FILLER_66_1991 ();
 FILLCELL_X32 FILLER_66_2023 ();
 FILLCELL_X32 FILLER_66_2055 ();
 FILLCELL_X32 FILLER_66_2087 ();
 FILLCELL_X32 FILLER_66_2119 ();
 FILLCELL_X32 FILLER_66_2151 ();
 FILLCELL_X32 FILLER_66_2183 ();
 FILLCELL_X32 FILLER_66_2215 ();
 FILLCELL_X32 FILLER_66_2247 ();
 FILLCELL_X32 FILLER_66_2279 ();
 FILLCELL_X32 FILLER_66_2311 ();
 FILLCELL_X32 FILLER_66_2343 ();
 FILLCELL_X32 FILLER_66_2375 ();
 FILLCELL_X16 FILLER_66_2407 ();
 FILLCELL_X8 FILLER_66_2423 ();
 FILLCELL_X4 FILLER_66_2431 ();
 FILLCELL_X1 FILLER_66_2435 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X32 FILLER_67_1776 ();
 FILLCELL_X32 FILLER_67_1808 ();
 FILLCELL_X32 FILLER_67_1840 ();
 FILLCELL_X32 FILLER_67_1872 ();
 FILLCELL_X32 FILLER_67_1904 ();
 FILLCELL_X32 FILLER_67_1936 ();
 FILLCELL_X32 FILLER_67_1968 ();
 FILLCELL_X32 FILLER_67_2000 ();
 FILLCELL_X32 FILLER_67_2032 ();
 FILLCELL_X32 FILLER_67_2064 ();
 FILLCELL_X32 FILLER_67_2096 ();
 FILLCELL_X32 FILLER_67_2128 ();
 FILLCELL_X32 FILLER_67_2160 ();
 FILLCELL_X32 FILLER_67_2192 ();
 FILLCELL_X32 FILLER_67_2224 ();
 FILLCELL_X32 FILLER_67_2256 ();
 FILLCELL_X32 FILLER_67_2288 ();
 FILLCELL_X32 FILLER_67_2320 ();
 FILLCELL_X32 FILLER_67_2352 ();
 FILLCELL_X32 FILLER_67_2384 ();
 FILLCELL_X16 FILLER_67_2416 ();
 FILLCELL_X4 FILLER_67_2432 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X32 FILLER_68_1592 ();
 FILLCELL_X32 FILLER_68_1624 ();
 FILLCELL_X32 FILLER_68_1656 ();
 FILLCELL_X32 FILLER_68_1688 ();
 FILLCELL_X32 FILLER_68_1720 ();
 FILLCELL_X32 FILLER_68_1752 ();
 FILLCELL_X32 FILLER_68_1784 ();
 FILLCELL_X32 FILLER_68_1816 ();
 FILLCELL_X32 FILLER_68_1848 ();
 FILLCELL_X8 FILLER_68_1880 ();
 FILLCELL_X4 FILLER_68_1888 ();
 FILLCELL_X2 FILLER_68_1892 ();
 FILLCELL_X32 FILLER_68_1895 ();
 FILLCELL_X32 FILLER_68_1927 ();
 FILLCELL_X32 FILLER_68_1959 ();
 FILLCELL_X32 FILLER_68_1991 ();
 FILLCELL_X32 FILLER_68_2023 ();
 FILLCELL_X32 FILLER_68_2055 ();
 FILLCELL_X32 FILLER_68_2087 ();
 FILLCELL_X32 FILLER_68_2119 ();
 FILLCELL_X32 FILLER_68_2151 ();
 FILLCELL_X32 FILLER_68_2183 ();
 FILLCELL_X32 FILLER_68_2215 ();
 FILLCELL_X32 FILLER_68_2247 ();
 FILLCELL_X32 FILLER_68_2279 ();
 FILLCELL_X32 FILLER_68_2311 ();
 FILLCELL_X32 FILLER_68_2343 ();
 FILLCELL_X32 FILLER_68_2375 ();
 FILLCELL_X16 FILLER_68_2407 ();
 FILLCELL_X8 FILLER_68_2423 ();
 FILLCELL_X4 FILLER_68_2431 ();
 FILLCELL_X1 FILLER_68_2435 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X32 FILLER_69_1776 ();
 FILLCELL_X32 FILLER_69_1808 ();
 FILLCELL_X32 FILLER_69_1840 ();
 FILLCELL_X32 FILLER_69_1872 ();
 FILLCELL_X32 FILLER_69_1904 ();
 FILLCELL_X32 FILLER_69_1936 ();
 FILLCELL_X32 FILLER_69_1968 ();
 FILLCELL_X32 FILLER_69_2000 ();
 FILLCELL_X32 FILLER_69_2032 ();
 FILLCELL_X32 FILLER_69_2064 ();
 FILLCELL_X32 FILLER_69_2096 ();
 FILLCELL_X32 FILLER_69_2128 ();
 FILLCELL_X32 FILLER_69_2160 ();
 FILLCELL_X32 FILLER_69_2192 ();
 FILLCELL_X32 FILLER_69_2224 ();
 FILLCELL_X32 FILLER_69_2256 ();
 FILLCELL_X32 FILLER_69_2288 ();
 FILLCELL_X32 FILLER_69_2320 ();
 FILLCELL_X32 FILLER_69_2352 ();
 FILLCELL_X32 FILLER_69_2384 ();
 FILLCELL_X16 FILLER_69_2416 ();
 FILLCELL_X4 FILLER_69_2432 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X32 FILLER_70_1784 ();
 FILLCELL_X32 FILLER_70_1816 ();
 FILLCELL_X32 FILLER_70_1848 ();
 FILLCELL_X8 FILLER_70_1880 ();
 FILLCELL_X4 FILLER_70_1888 ();
 FILLCELL_X2 FILLER_70_1892 ();
 FILLCELL_X32 FILLER_70_1895 ();
 FILLCELL_X32 FILLER_70_1927 ();
 FILLCELL_X32 FILLER_70_1959 ();
 FILLCELL_X32 FILLER_70_1991 ();
 FILLCELL_X32 FILLER_70_2023 ();
 FILLCELL_X32 FILLER_70_2055 ();
 FILLCELL_X32 FILLER_70_2087 ();
 FILLCELL_X32 FILLER_70_2119 ();
 FILLCELL_X32 FILLER_70_2151 ();
 FILLCELL_X32 FILLER_70_2183 ();
 FILLCELL_X32 FILLER_70_2215 ();
 FILLCELL_X32 FILLER_70_2247 ();
 FILLCELL_X32 FILLER_70_2279 ();
 FILLCELL_X32 FILLER_70_2311 ();
 FILLCELL_X32 FILLER_70_2343 ();
 FILLCELL_X32 FILLER_70_2375 ();
 FILLCELL_X16 FILLER_70_2407 ();
 FILLCELL_X8 FILLER_70_2423 ();
 FILLCELL_X4 FILLER_70_2431 ();
 FILLCELL_X1 FILLER_70_2435 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X32 FILLER_71_1776 ();
 FILLCELL_X32 FILLER_71_1808 ();
 FILLCELL_X32 FILLER_71_1840 ();
 FILLCELL_X32 FILLER_71_1872 ();
 FILLCELL_X32 FILLER_71_1904 ();
 FILLCELL_X32 FILLER_71_1936 ();
 FILLCELL_X32 FILLER_71_1968 ();
 FILLCELL_X32 FILLER_71_2000 ();
 FILLCELL_X32 FILLER_71_2032 ();
 FILLCELL_X32 FILLER_71_2064 ();
 FILLCELL_X32 FILLER_71_2096 ();
 FILLCELL_X32 FILLER_71_2128 ();
 FILLCELL_X32 FILLER_71_2160 ();
 FILLCELL_X32 FILLER_71_2192 ();
 FILLCELL_X32 FILLER_71_2224 ();
 FILLCELL_X32 FILLER_71_2256 ();
 FILLCELL_X32 FILLER_71_2288 ();
 FILLCELL_X32 FILLER_71_2320 ();
 FILLCELL_X32 FILLER_71_2352 ();
 FILLCELL_X32 FILLER_71_2384 ();
 FILLCELL_X16 FILLER_71_2416 ();
 FILLCELL_X4 FILLER_71_2432 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X32 FILLER_72_1784 ();
 FILLCELL_X32 FILLER_72_1816 ();
 FILLCELL_X32 FILLER_72_1848 ();
 FILLCELL_X8 FILLER_72_1880 ();
 FILLCELL_X4 FILLER_72_1888 ();
 FILLCELL_X2 FILLER_72_1892 ();
 FILLCELL_X32 FILLER_72_1895 ();
 FILLCELL_X32 FILLER_72_1927 ();
 FILLCELL_X32 FILLER_72_1959 ();
 FILLCELL_X32 FILLER_72_1991 ();
 FILLCELL_X32 FILLER_72_2023 ();
 FILLCELL_X32 FILLER_72_2055 ();
 FILLCELL_X32 FILLER_72_2087 ();
 FILLCELL_X32 FILLER_72_2119 ();
 FILLCELL_X32 FILLER_72_2151 ();
 FILLCELL_X32 FILLER_72_2183 ();
 FILLCELL_X32 FILLER_72_2215 ();
 FILLCELL_X32 FILLER_72_2247 ();
 FILLCELL_X32 FILLER_72_2279 ();
 FILLCELL_X32 FILLER_72_2311 ();
 FILLCELL_X32 FILLER_72_2343 ();
 FILLCELL_X32 FILLER_72_2375 ();
 FILLCELL_X16 FILLER_72_2407 ();
 FILLCELL_X8 FILLER_72_2423 ();
 FILLCELL_X4 FILLER_72_2431 ();
 FILLCELL_X1 FILLER_72_2435 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X32 FILLER_73_1776 ();
 FILLCELL_X32 FILLER_73_1808 ();
 FILLCELL_X32 FILLER_73_1840 ();
 FILLCELL_X32 FILLER_73_1872 ();
 FILLCELL_X32 FILLER_73_1904 ();
 FILLCELL_X32 FILLER_73_1936 ();
 FILLCELL_X32 FILLER_73_1968 ();
 FILLCELL_X32 FILLER_73_2000 ();
 FILLCELL_X32 FILLER_73_2032 ();
 FILLCELL_X32 FILLER_73_2064 ();
 FILLCELL_X32 FILLER_73_2096 ();
 FILLCELL_X32 FILLER_73_2128 ();
 FILLCELL_X32 FILLER_73_2160 ();
 FILLCELL_X32 FILLER_73_2192 ();
 FILLCELL_X32 FILLER_73_2224 ();
 FILLCELL_X32 FILLER_73_2256 ();
 FILLCELL_X32 FILLER_73_2288 ();
 FILLCELL_X32 FILLER_73_2320 ();
 FILLCELL_X32 FILLER_73_2352 ();
 FILLCELL_X32 FILLER_73_2384 ();
 FILLCELL_X16 FILLER_73_2416 ();
 FILLCELL_X4 FILLER_73_2432 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X32 FILLER_74_1784 ();
 FILLCELL_X32 FILLER_74_1816 ();
 FILLCELL_X32 FILLER_74_1848 ();
 FILLCELL_X8 FILLER_74_1880 ();
 FILLCELL_X4 FILLER_74_1888 ();
 FILLCELL_X2 FILLER_74_1892 ();
 FILLCELL_X32 FILLER_74_1895 ();
 FILLCELL_X32 FILLER_74_1927 ();
 FILLCELL_X32 FILLER_74_1959 ();
 FILLCELL_X32 FILLER_74_1991 ();
 FILLCELL_X32 FILLER_74_2023 ();
 FILLCELL_X32 FILLER_74_2055 ();
 FILLCELL_X32 FILLER_74_2087 ();
 FILLCELL_X32 FILLER_74_2119 ();
 FILLCELL_X32 FILLER_74_2151 ();
 FILLCELL_X32 FILLER_74_2183 ();
 FILLCELL_X32 FILLER_74_2215 ();
 FILLCELL_X32 FILLER_74_2247 ();
 FILLCELL_X32 FILLER_74_2279 ();
 FILLCELL_X32 FILLER_74_2311 ();
 FILLCELL_X32 FILLER_74_2343 ();
 FILLCELL_X32 FILLER_74_2375 ();
 FILLCELL_X16 FILLER_74_2407 ();
 FILLCELL_X8 FILLER_74_2423 ();
 FILLCELL_X4 FILLER_74_2431 ();
 FILLCELL_X1 FILLER_74_2435 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X32 FILLER_75_1776 ();
 FILLCELL_X32 FILLER_75_1808 ();
 FILLCELL_X32 FILLER_75_1840 ();
 FILLCELL_X32 FILLER_75_1872 ();
 FILLCELL_X32 FILLER_75_1904 ();
 FILLCELL_X32 FILLER_75_1936 ();
 FILLCELL_X32 FILLER_75_1968 ();
 FILLCELL_X32 FILLER_75_2000 ();
 FILLCELL_X32 FILLER_75_2032 ();
 FILLCELL_X32 FILLER_75_2064 ();
 FILLCELL_X32 FILLER_75_2096 ();
 FILLCELL_X32 FILLER_75_2128 ();
 FILLCELL_X32 FILLER_75_2160 ();
 FILLCELL_X32 FILLER_75_2192 ();
 FILLCELL_X32 FILLER_75_2224 ();
 FILLCELL_X32 FILLER_75_2256 ();
 FILLCELL_X32 FILLER_75_2288 ();
 FILLCELL_X32 FILLER_75_2320 ();
 FILLCELL_X32 FILLER_75_2352 ();
 FILLCELL_X32 FILLER_75_2384 ();
 FILLCELL_X16 FILLER_75_2416 ();
 FILLCELL_X4 FILLER_75_2432 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X32 FILLER_76_1592 ();
 FILLCELL_X32 FILLER_76_1624 ();
 FILLCELL_X32 FILLER_76_1656 ();
 FILLCELL_X32 FILLER_76_1688 ();
 FILLCELL_X32 FILLER_76_1720 ();
 FILLCELL_X32 FILLER_76_1752 ();
 FILLCELL_X32 FILLER_76_1784 ();
 FILLCELL_X32 FILLER_76_1816 ();
 FILLCELL_X32 FILLER_76_1848 ();
 FILLCELL_X8 FILLER_76_1880 ();
 FILLCELL_X4 FILLER_76_1888 ();
 FILLCELL_X2 FILLER_76_1892 ();
 FILLCELL_X32 FILLER_76_1895 ();
 FILLCELL_X32 FILLER_76_1927 ();
 FILLCELL_X32 FILLER_76_1959 ();
 FILLCELL_X32 FILLER_76_1991 ();
 FILLCELL_X32 FILLER_76_2023 ();
 FILLCELL_X32 FILLER_76_2055 ();
 FILLCELL_X32 FILLER_76_2087 ();
 FILLCELL_X32 FILLER_76_2119 ();
 FILLCELL_X32 FILLER_76_2151 ();
 FILLCELL_X32 FILLER_76_2183 ();
 FILLCELL_X32 FILLER_76_2215 ();
 FILLCELL_X32 FILLER_76_2247 ();
 FILLCELL_X32 FILLER_76_2279 ();
 FILLCELL_X32 FILLER_76_2311 ();
 FILLCELL_X32 FILLER_76_2343 ();
 FILLCELL_X32 FILLER_76_2375 ();
 FILLCELL_X16 FILLER_76_2407 ();
 FILLCELL_X8 FILLER_76_2423 ();
 FILLCELL_X4 FILLER_76_2431 ();
 FILLCELL_X1 FILLER_76_2435 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X32 FILLER_77_1776 ();
 FILLCELL_X32 FILLER_77_1808 ();
 FILLCELL_X32 FILLER_77_1840 ();
 FILLCELL_X32 FILLER_77_1872 ();
 FILLCELL_X32 FILLER_77_1904 ();
 FILLCELL_X32 FILLER_77_1936 ();
 FILLCELL_X32 FILLER_77_1968 ();
 FILLCELL_X32 FILLER_77_2000 ();
 FILLCELL_X32 FILLER_77_2032 ();
 FILLCELL_X32 FILLER_77_2064 ();
 FILLCELL_X32 FILLER_77_2096 ();
 FILLCELL_X32 FILLER_77_2128 ();
 FILLCELL_X32 FILLER_77_2160 ();
 FILLCELL_X32 FILLER_77_2192 ();
 FILLCELL_X32 FILLER_77_2224 ();
 FILLCELL_X32 FILLER_77_2256 ();
 FILLCELL_X32 FILLER_77_2288 ();
 FILLCELL_X32 FILLER_77_2320 ();
 FILLCELL_X32 FILLER_77_2352 ();
 FILLCELL_X32 FILLER_77_2384 ();
 FILLCELL_X16 FILLER_77_2416 ();
 FILLCELL_X4 FILLER_77_2432 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X32 FILLER_78_1592 ();
 FILLCELL_X32 FILLER_78_1624 ();
 FILLCELL_X32 FILLER_78_1656 ();
 FILLCELL_X32 FILLER_78_1688 ();
 FILLCELL_X32 FILLER_78_1720 ();
 FILLCELL_X32 FILLER_78_1752 ();
 FILLCELL_X32 FILLER_78_1784 ();
 FILLCELL_X32 FILLER_78_1816 ();
 FILLCELL_X32 FILLER_78_1848 ();
 FILLCELL_X8 FILLER_78_1880 ();
 FILLCELL_X4 FILLER_78_1888 ();
 FILLCELL_X2 FILLER_78_1892 ();
 FILLCELL_X32 FILLER_78_1895 ();
 FILLCELL_X32 FILLER_78_1927 ();
 FILLCELL_X32 FILLER_78_1959 ();
 FILLCELL_X32 FILLER_78_1991 ();
 FILLCELL_X32 FILLER_78_2023 ();
 FILLCELL_X32 FILLER_78_2055 ();
 FILLCELL_X32 FILLER_78_2087 ();
 FILLCELL_X32 FILLER_78_2119 ();
 FILLCELL_X32 FILLER_78_2151 ();
 FILLCELL_X32 FILLER_78_2183 ();
 FILLCELL_X32 FILLER_78_2215 ();
 FILLCELL_X32 FILLER_78_2247 ();
 FILLCELL_X32 FILLER_78_2279 ();
 FILLCELL_X32 FILLER_78_2311 ();
 FILLCELL_X32 FILLER_78_2343 ();
 FILLCELL_X32 FILLER_78_2375 ();
 FILLCELL_X16 FILLER_78_2407 ();
 FILLCELL_X8 FILLER_78_2423 ();
 FILLCELL_X4 FILLER_78_2431 ();
 FILLCELL_X1 FILLER_78_2435 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X32 FILLER_79_1776 ();
 FILLCELL_X32 FILLER_79_1808 ();
 FILLCELL_X32 FILLER_79_1840 ();
 FILLCELL_X32 FILLER_79_1872 ();
 FILLCELL_X32 FILLER_79_1904 ();
 FILLCELL_X32 FILLER_79_1936 ();
 FILLCELL_X32 FILLER_79_1968 ();
 FILLCELL_X32 FILLER_79_2000 ();
 FILLCELL_X32 FILLER_79_2032 ();
 FILLCELL_X32 FILLER_79_2064 ();
 FILLCELL_X32 FILLER_79_2096 ();
 FILLCELL_X32 FILLER_79_2128 ();
 FILLCELL_X32 FILLER_79_2160 ();
 FILLCELL_X32 FILLER_79_2192 ();
 FILLCELL_X32 FILLER_79_2224 ();
 FILLCELL_X32 FILLER_79_2256 ();
 FILLCELL_X32 FILLER_79_2288 ();
 FILLCELL_X32 FILLER_79_2320 ();
 FILLCELL_X32 FILLER_79_2352 ();
 FILLCELL_X32 FILLER_79_2384 ();
 FILLCELL_X16 FILLER_79_2416 ();
 FILLCELL_X4 FILLER_79_2432 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X32 FILLER_80_1592 ();
 FILLCELL_X32 FILLER_80_1624 ();
 FILLCELL_X32 FILLER_80_1656 ();
 FILLCELL_X32 FILLER_80_1688 ();
 FILLCELL_X32 FILLER_80_1720 ();
 FILLCELL_X32 FILLER_80_1752 ();
 FILLCELL_X32 FILLER_80_1784 ();
 FILLCELL_X32 FILLER_80_1816 ();
 FILLCELL_X32 FILLER_80_1848 ();
 FILLCELL_X8 FILLER_80_1880 ();
 FILLCELL_X4 FILLER_80_1888 ();
 FILLCELL_X2 FILLER_80_1892 ();
 FILLCELL_X32 FILLER_80_1895 ();
 FILLCELL_X32 FILLER_80_1927 ();
 FILLCELL_X32 FILLER_80_1959 ();
 FILLCELL_X32 FILLER_80_1991 ();
 FILLCELL_X32 FILLER_80_2023 ();
 FILLCELL_X32 FILLER_80_2055 ();
 FILLCELL_X32 FILLER_80_2087 ();
 FILLCELL_X32 FILLER_80_2119 ();
 FILLCELL_X32 FILLER_80_2151 ();
 FILLCELL_X32 FILLER_80_2183 ();
 FILLCELL_X32 FILLER_80_2215 ();
 FILLCELL_X32 FILLER_80_2247 ();
 FILLCELL_X32 FILLER_80_2279 ();
 FILLCELL_X32 FILLER_80_2311 ();
 FILLCELL_X32 FILLER_80_2343 ();
 FILLCELL_X32 FILLER_80_2375 ();
 FILLCELL_X16 FILLER_80_2407 ();
 FILLCELL_X8 FILLER_80_2423 ();
 FILLCELL_X4 FILLER_80_2431 ();
 FILLCELL_X1 FILLER_80_2435 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X32 FILLER_81_1776 ();
 FILLCELL_X32 FILLER_81_1808 ();
 FILLCELL_X32 FILLER_81_1840 ();
 FILLCELL_X32 FILLER_81_1872 ();
 FILLCELL_X32 FILLER_81_1904 ();
 FILLCELL_X32 FILLER_81_1936 ();
 FILLCELL_X32 FILLER_81_1968 ();
 FILLCELL_X32 FILLER_81_2000 ();
 FILLCELL_X32 FILLER_81_2032 ();
 FILLCELL_X32 FILLER_81_2064 ();
 FILLCELL_X32 FILLER_81_2096 ();
 FILLCELL_X32 FILLER_81_2128 ();
 FILLCELL_X32 FILLER_81_2160 ();
 FILLCELL_X32 FILLER_81_2192 ();
 FILLCELL_X32 FILLER_81_2224 ();
 FILLCELL_X32 FILLER_81_2256 ();
 FILLCELL_X32 FILLER_81_2288 ();
 FILLCELL_X32 FILLER_81_2320 ();
 FILLCELL_X32 FILLER_81_2352 ();
 FILLCELL_X32 FILLER_81_2384 ();
 FILLCELL_X16 FILLER_81_2416 ();
 FILLCELL_X4 FILLER_81_2432 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X32 FILLER_82_1784 ();
 FILLCELL_X32 FILLER_82_1816 ();
 FILLCELL_X32 FILLER_82_1848 ();
 FILLCELL_X8 FILLER_82_1880 ();
 FILLCELL_X4 FILLER_82_1888 ();
 FILLCELL_X2 FILLER_82_1892 ();
 FILLCELL_X32 FILLER_82_1895 ();
 FILLCELL_X32 FILLER_82_1927 ();
 FILLCELL_X32 FILLER_82_1959 ();
 FILLCELL_X32 FILLER_82_1991 ();
 FILLCELL_X32 FILLER_82_2023 ();
 FILLCELL_X32 FILLER_82_2055 ();
 FILLCELL_X32 FILLER_82_2087 ();
 FILLCELL_X32 FILLER_82_2119 ();
 FILLCELL_X32 FILLER_82_2151 ();
 FILLCELL_X32 FILLER_82_2183 ();
 FILLCELL_X32 FILLER_82_2215 ();
 FILLCELL_X32 FILLER_82_2247 ();
 FILLCELL_X32 FILLER_82_2279 ();
 FILLCELL_X32 FILLER_82_2311 ();
 FILLCELL_X32 FILLER_82_2343 ();
 FILLCELL_X32 FILLER_82_2375 ();
 FILLCELL_X16 FILLER_82_2407 ();
 FILLCELL_X8 FILLER_82_2423 ();
 FILLCELL_X4 FILLER_82_2431 ();
 FILLCELL_X1 FILLER_82_2435 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X32 FILLER_83_1776 ();
 FILLCELL_X32 FILLER_83_1808 ();
 FILLCELL_X32 FILLER_83_1840 ();
 FILLCELL_X32 FILLER_83_1872 ();
 FILLCELL_X32 FILLER_83_1904 ();
 FILLCELL_X32 FILLER_83_1936 ();
 FILLCELL_X32 FILLER_83_1968 ();
 FILLCELL_X32 FILLER_83_2000 ();
 FILLCELL_X32 FILLER_83_2032 ();
 FILLCELL_X32 FILLER_83_2064 ();
 FILLCELL_X32 FILLER_83_2096 ();
 FILLCELL_X32 FILLER_83_2128 ();
 FILLCELL_X32 FILLER_83_2160 ();
 FILLCELL_X32 FILLER_83_2192 ();
 FILLCELL_X32 FILLER_83_2224 ();
 FILLCELL_X32 FILLER_83_2256 ();
 FILLCELL_X32 FILLER_83_2288 ();
 FILLCELL_X32 FILLER_83_2320 ();
 FILLCELL_X32 FILLER_83_2352 ();
 FILLCELL_X32 FILLER_83_2384 ();
 FILLCELL_X16 FILLER_83_2416 ();
 FILLCELL_X4 FILLER_83_2432 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X32 FILLER_84_1784 ();
 FILLCELL_X32 FILLER_84_1816 ();
 FILLCELL_X32 FILLER_84_1848 ();
 FILLCELL_X8 FILLER_84_1880 ();
 FILLCELL_X4 FILLER_84_1888 ();
 FILLCELL_X2 FILLER_84_1892 ();
 FILLCELL_X32 FILLER_84_1895 ();
 FILLCELL_X32 FILLER_84_1927 ();
 FILLCELL_X32 FILLER_84_1959 ();
 FILLCELL_X32 FILLER_84_1991 ();
 FILLCELL_X32 FILLER_84_2023 ();
 FILLCELL_X32 FILLER_84_2055 ();
 FILLCELL_X32 FILLER_84_2087 ();
 FILLCELL_X32 FILLER_84_2119 ();
 FILLCELL_X32 FILLER_84_2151 ();
 FILLCELL_X32 FILLER_84_2183 ();
 FILLCELL_X32 FILLER_84_2215 ();
 FILLCELL_X32 FILLER_84_2247 ();
 FILLCELL_X32 FILLER_84_2279 ();
 FILLCELL_X32 FILLER_84_2311 ();
 FILLCELL_X32 FILLER_84_2343 ();
 FILLCELL_X32 FILLER_84_2375 ();
 FILLCELL_X16 FILLER_84_2407 ();
 FILLCELL_X8 FILLER_84_2423 ();
 FILLCELL_X4 FILLER_84_2431 ();
 FILLCELL_X1 FILLER_84_2435 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X32 FILLER_85_1776 ();
 FILLCELL_X32 FILLER_85_1808 ();
 FILLCELL_X32 FILLER_85_1840 ();
 FILLCELL_X32 FILLER_85_1872 ();
 FILLCELL_X32 FILLER_85_1904 ();
 FILLCELL_X32 FILLER_85_1936 ();
 FILLCELL_X32 FILLER_85_1968 ();
 FILLCELL_X32 FILLER_85_2000 ();
 FILLCELL_X32 FILLER_85_2032 ();
 FILLCELL_X32 FILLER_85_2064 ();
 FILLCELL_X32 FILLER_85_2096 ();
 FILLCELL_X32 FILLER_85_2128 ();
 FILLCELL_X32 FILLER_85_2160 ();
 FILLCELL_X32 FILLER_85_2192 ();
 FILLCELL_X32 FILLER_85_2224 ();
 FILLCELL_X32 FILLER_85_2256 ();
 FILLCELL_X32 FILLER_85_2288 ();
 FILLCELL_X32 FILLER_85_2320 ();
 FILLCELL_X32 FILLER_85_2352 ();
 FILLCELL_X32 FILLER_85_2384 ();
 FILLCELL_X16 FILLER_85_2416 ();
 FILLCELL_X4 FILLER_85_2432 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X32 FILLER_86_1784 ();
 FILLCELL_X32 FILLER_86_1816 ();
 FILLCELL_X32 FILLER_86_1848 ();
 FILLCELL_X8 FILLER_86_1880 ();
 FILLCELL_X4 FILLER_86_1888 ();
 FILLCELL_X2 FILLER_86_1892 ();
 FILLCELL_X32 FILLER_86_1895 ();
 FILLCELL_X32 FILLER_86_1927 ();
 FILLCELL_X32 FILLER_86_1959 ();
 FILLCELL_X32 FILLER_86_1991 ();
 FILLCELL_X32 FILLER_86_2023 ();
 FILLCELL_X32 FILLER_86_2055 ();
 FILLCELL_X32 FILLER_86_2087 ();
 FILLCELL_X32 FILLER_86_2119 ();
 FILLCELL_X32 FILLER_86_2151 ();
 FILLCELL_X32 FILLER_86_2183 ();
 FILLCELL_X32 FILLER_86_2215 ();
 FILLCELL_X32 FILLER_86_2247 ();
 FILLCELL_X32 FILLER_86_2279 ();
 FILLCELL_X32 FILLER_86_2311 ();
 FILLCELL_X32 FILLER_86_2343 ();
 FILLCELL_X32 FILLER_86_2375 ();
 FILLCELL_X16 FILLER_86_2407 ();
 FILLCELL_X8 FILLER_86_2423 ();
 FILLCELL_X4 FILLER_86_2431 ();
 FILLCELL_X1 FILLER_86_2435 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X32 FILLER_87_1776 ();
 FILLCELL_X32 FILLER_87_1808 ();
 FILLCELL_X32 FILLER_87_1840 ();
 FILLCELL_X32 FILLER_87_1872 ();
 FILLCELL_X32 FILLER_87_1904 ();
 FILLCELL_X32 FILLER_87_1936 ();
 FILLCELL_X32 FILLER_87_1968 ();
 FILLCELL_X32 FILLER_87_2000 ();
 FILLCELL_X32 FILLER_87_2032 ();
 FILLCELL_X32 FILLER_87_2064 ();
 FILLCELL_X32 FILLER_87_2096 ();
 FILLCELL_X32 FILLER_87_2128 ();
 FILLCELL_X32 FILLER_87_2160 ();
 FILLCELL_X32 FILLER_87_2192 ();
 FILLCELL_X32 FILLER_87_2224 ();
 FILLCELL_X32 FILLER_87_2256 ();
 FILLCELL_X32 FILLER_87_2288 ();
 FILLCELL_X32 FILLER_87_2320 ();
 FILLCELL_X32 FILLER_87_2352 ();
 FILLCELL_X32 FILLER_87_2384 ();
 FILLCELL_X16 FILLER_87_2416 ();
 FILLCELL_X4 FILLER_87_2432 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X32 FILLER_88_1784 ();
 FILLCELL_X32 FILLER_88_1816 ();
 FILLCELL_X32 FILLER_88_1848 ();
 FILLCELL_X8 FILLER_88_1880 ();
 FILLCELL_X4 FILLER_88_1888 ();
 FILLCELL_X2 FILLER_88_1892 ();
 FILLCELL_X32 FILLER_88_1895 ();
 FILLCELL_X32 FILLER_88_1927 ();
 FILLCELL_X32 FILLER_88_1959 ();
 FILLCELL_X32 FILLER_88_1991 ();
 FILLCELL_X32 FILLER_88_2023 ();
 FILLCELL_X32 FILLER_88_2055 ();
 FILLCELL_X32 FILLER_88_2087 ();
 FILLCELL_X32 FILLER_88_2119 ();
 FILLCELL_X32 FILLER_88_2151 ();
 FILLCELL_X32 FILLER_88_2183 ();
 FILLCELL_X32 FILLER_88_2215 ();
 FILLCELL_X32 FILLER_88_2247 ();
 FILLCELL_X32 FILLER_88_2279 ();
 FILLCELL_X32 FILLER_88_2311 ();
 FILLCELL_X32 FILLER_88_2343 ();
 FILLCELL_X32 FILLER_88_2375 ();
 FILLCELL_X16 FILLER_88_2407 ();
 FILLCELL_X8 FILLER_88_2423 ();
 FILLCELL_X4 FILLER_88_2431 ();
 FILLCELL_X1 FILLER_88_2435 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X32 FILLER_89_1776 ();
 FILLCELL_X32 FILLER_89_1808 ();
 FILLCELL_X32 FILLER_89_1840 ();
 FILLCELL_X32 FILLER_89_1872 ();
 FILLCELL_X32 FILLER_89_1904 ();
 FILLCELL_X32 FILLER_89_1936 ();
 FILLCELL_X32 FILLER_89_1968 ();
 FILLCELL_X32 FILLER_89_2000 ();
 FILLCELL_X32 FILLER_89_2032 ();
 FILLCELL_X32 FILLER_89_2064 ();
 FILLCELL_X32 FILLER_89_2096 ();
 FILLCELL_X32 FILLER_89_2128 ();
 FILLCELL_X32 FILLER_89_2160 ();
 FILLCELL_X32 FILLER_89_2192 ();
 FILLCELL_X32 FILLER_89_2224 ();
 FILLCELL_X32 FILLER_89_2256 ();
 FILLCELL_X32 FILLER_89_2288 ();
 FILLCELL_X32 FILLER_89_2320 ();
 FILLCELL_X32 FILLER_89_2352 ();
 FILLCELL_X32 FILLER_89_2384 ();
 FILLCELL_X16 FILLER_89_2416 ();
 FILLCELL_X4 FILLER_89_2432 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X32 FILLER_90_1784 ();
 FILLCELL_X32 FILLER_90_1816 ();
 FILLCELL_X32 FILLER_90_1848 ();
 FILLCELL_X8 FILLER_90_1880 ();
 FILLCELL_X4 FILLER_90_1888 ();
 FILLCELL_X2 FILLER_90_1892 ();
 FILLCELL_X32 FILLER_90_1895 ();
 FILLCELL_X32 FILLER_90_1927 ();
 FILLCELL_X32 FILLER_90_1959 ();
 FILLCELL_X32 FILLER_90_1991 ();
 FILLCELL_X32 FILLER_90_2023 ();
 FILLCELL_X32 FILLER_90_2055 ();
 FILLCELL_X32 FILLER_90_2087 ();
 FILLCELL_X32 FILLER_90_2119 ();
 FILLCELL_X32 FILLER_90_2151 ();
 FILLCELL_X32 FILLER_90_2183 ();
 FILLCELL_X32 FILLER_90_2215 ();
 FILLCELL_X32 FILLER_90_2247 ();
 FILLCELL_X32 FILLER_90_2279 ();
 FILLCELL_X32 FILLER_90_2311 ();
 FILLCELL_X32 FILLER_90_2343 ();
 FILLCELL_X32 FILLER_90_2375 ();
 FILLCELL_X16 FILLER_90_2407 ();
 FILLCELL_X8 FILLER_90_2423 ();
 FILLCELL_X4 FILLER_90_2431 ();
 FILLCELL_X1 FILLER_90_2435 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X32 FILLER_91_1776 ();
 FILLCELL_X32 FILLER_91_1808 ();
 FILLCELL_X32 FILLER_91_1840 ();
 FILLCELL_X32 FILLER_91_1872 ();
 FILLCELL_X32 FILLER_91_1904 ();
 FILLCELL_X32 FILLER_91_1936 ();
 FILLCELL_X32 FILLER_91_1968 ();
 FILLCELL_X32 FILLER_91_2000 ();
 FILLCELL_X32 FILLER_91_2032 ();
 FILLCELL_X32 FILLER_91_2064 ();
 FILLCELL_X32 FILLER_91_2096 ();
 FILLCELL_X32 FILLER_91_2128 ();
 FILLCELL_X32 FILLER_91_2160 ();
 FILLCELL_X32 FILLER_91_2192 ();
 FILLCELL_X32 FILLER_91_2224 ();
 FILLCELL_X32 FILLER_91_2256 ();
 FILLCELL_X32 FILLER_91_2288 ();
 FILLCELL_X32 FILLER_91_2320 ();
 FILLCELL_X32 FILLER_91_2352 ();
 FILLCELL_X32 FILLER_91_2384 ();
 FILLCELL_X16 FILLER_91_2416 ();
 FILLCELL_X4 FILLER_91_2432 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X32 FILLER_92_1784 ();
 FILLCELL_X32 FILLER_92_1816 ();
 FILLCELL_X32 FILLER_92_1848 ();
 FILLCELL_X8 FILLER_92_1880 ();
 FILLCELL_X4 FILLER_92_1888 ();
 FILLCELL_X2 FILLER_92_1892 ();
 FILLCELL_X32 FILLER_92_1895 ();
 FILLCELL_X32 FILLER_92_1927 ();
 FILLCELL_X32 FILLER_92_1959 ();
 FILLCELL_X32 FILLER_92_1991 ();
 FILLCELL_X32 FILLER_92_2023 ();
 FILLCELL_X32 FILLER_92_2055 ();
 FILLCELL_X32 FILLER_92_2087 ();
 FILLCELL_X32 FILLER_92_2119 ();
 FILLCELL_X32 FILLER_92_2151 ();
 FILLCELL_X32 FILLER_92_2183 ();
 FILLCELL_X32 FILLER_92_2215 ();
 FILLCELL_X32 FILLER_92_2247 ();
 FILLCELL_X32 FILLER_92_2279 ();
 FILLCELL_X32 FILLER_92_2311 ();
 FILLCELL_X32 FILLER_92_2343 ();
 FILLCELL_X32 FILLER_92_2375 ();
 FILLCELL_X16 FILLER_92_2407 ();
 FILLCELL_X8 FILLER_92_2423 ();
 FILLCELL_X4 FILLER_92_2431 ();
 FILLCELL_X1 FILLER_92_2435 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X32 FILLER_93_1776 ();
 FILLCELL_X32 FILLER_93_1808 ();
 FILLCELL_X32 FILLER_93_1840 ();
 FILLCELL_X32 FILLER_93_1872 ();
 FILLCELL_X32 FILLER_93_1904 ();
 FILLCELL_X32 FILLER_93_1936 ();
 FILLCELL_X32 FILLER_93_1968 ();
 FILLCELL_X32 FILLER_93_2000 ();
 FILLCELL_X32 FILLER_93_2032 ();
 FILLCELL_X32 FILLER_93_2064 ();
 FILLCELL_X32 FILLER_93_2096 ();
 FILLCELL_X32 FILLER_93_2128 ();
 FILLCELL_X32 FILLER_93_2160 ();
 FILLCELL_X32 FILLER_93_2192 ();
 FILLCELL_X32 FILLER_93_2224 ();
 FILLCELL_X32 FILLER_93_2256 ();
 FILLCELL_X32 FILLER_93_2288 ();
 FILLCELL_X32 FILLER_93_2320 ();
 FILLCELL_X32 FILLER_93_2352 ();
 FILLCELL_X32 FILLER_93_2384 ();
 FILLCELL_X16 FILLER_93_2416 ();
 FILLCELL_X4 FILLER_93_2432 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X32 FILLER_94_1784 ();
 FILLCELL_X32 FILLER_94_1816 ();
 FILLCELL_X32 FILLER_94_1848 ();
 FILLCELL_X8 FILLER_94_1880 ();
 FILLCELL_X4 FILLER_94_1888 ();
 FILLCELL_X2 FILLER_94_1892 ();
 FILLCELL_X32 FILLER_94_1895 ();
 FILLCELL_X32 FILLER_94_1927 ();
 FILLCELL_X32 FILLER_94_1959 ();
 FILLCELL_X32 FILLER_94_1991 ();
 FILLCELL_X32 FILLER_94_2023 ();
 FILLCELL_X32 FILLER_94_2055 ();
 FILLCELL_X32 FILLER_94_2087 ();
 FILLCELL_X32 FILLER_94_2119 ();
 FILLCELL_X32 FILLER_94_2151 ();
 FILLCELL_X32 FILLER_94_2183 ();
 FILLCELL_X32 FILLER_94_2215 ();
 FILLCELL_X32 FILLER_94_2247 ();
 FILLCELL_X32 FILLER_94_2279 ();
 FILLCELL_X32 FILLER_94_2311 ();
 FILLCELL_X32 FILLER_94_2343 ();
 FILLCELL_X32 FILLER_94_2375 ();
 FILLCELL_X16 FILLER_94_2407 ();
 FILLCELL_X8 FILLER_94_2423 ();
 FILLCELL_X4 FILLER_94_2431 ();
 FILLCELL_X1 FILLER_94_2435 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X32 FILLER_95_1776 ();
 FILLCELL_X32 FILLER_95_1808 ();
 FILLCELL_X32 FILLER_95_1840 ();
 FILLCELL_X32 FILLER_95_1872 ();
 FILLCELL_X32 FILLER_95_1904 ();
 FILLCELL_X32 FILLER_95_1936 ();
 FILLCELL_X32 FILLER_95_1968 ();
 FILLCELL_X32 FILLER_95_2000 ();
 FILLCELL_X32 FILLER_95_2032 ();
 FILLCELL_X32 FILLER_95_2064 ();
 FILLCELL_X32 FILLER_95_2096 ();
 FILLCELL_X32 FILLER_95_2128 ();
 FILLCELL_X32 FILLER_95_2160 ();
 FILLCELL_X32 FILLER_95_2192 ();
 FILLCELL_X32 FILLER_95_2224 ();
 FILLCELL_X32 FILLER_95_2256 ();
 FILLCELL_X32 FILLER_95_2288 ();
 FILLCELL_X32 FILLER_95_2320 ();
 FILLCELL_X32 FILLER_95_2352 ();
 FILLCELL_X32 FILLER_95_2384 ();
 FILLCELL_X16 FILLER_95_2416 ();
 FILLCELL_X4 FILLER_95_2432 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X32 FILLER_96_1784 ();
 FILLCELL_X32 FILLER_96_1816 ();
 FILLCELL_X32 FILLER_96_1848 ();
 FILLCELL_X8 FILLER_96_1880 ();
 FILLCELL_X4 FILLER_96_1888 ();
 FILLCELL_X2 FILLER_96_1892 ();
 FILLCELL_X32 FILLER_96_1895 ();
 FILLCELL_X32 FILLER_96_1927 ();
 FILLCELL_X32 FILLER_96_1959 ();
 FILLCELL_X32 FILLER_96_1991 ();
 FILLCELL_X32 FILLER_96_2023 ();
 FILLCELL_X32 FILLER_96_2055 ();
 FILLCELL_X32 FILLER_96_2087 ();
 FILLCELL_X32 FILLER_96_2119 ();
 FILLCELL_X32 FILLER_96_2151 ();
 FILLCELL_X32 FILLER_96_2183 ();
 FILLCELL_X32 FILLER_96_2215 ();
 FILLCELL_X32 FILLER_96_2247 ();
 FILLCELL_X32 FILLER_96_2279 ();
 FILLCELL_X32 FILLER_96_2311 ();
 FILLCELL_X32 FILLER_96_2343 ();
 FILLCELL_X32 FILLER_96_2375 ();
 FILLCELL_X16 FILLER_96_2407 ();
 FILLCELL_X8 FILLER_96_2423 ();
 FILLCELL_X4 FILLER_96_2431 ();
 FILLCELL_X1 FILLER_96_2435 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X32 FILLER_97_1776 ();
 FILLCELL_X32 FILLER_97_1808 ();
 FILLCELL_X32 FILLER_97_1840 ();
 FILLCELL_X32 FILLER_97_1872 ();
 FILLCELL_X32 FILLER_97_1904 ();
 FILLCELL_X32 FILLER_97_1936 ();
 FILLCELL_X32 FILLER_97_1968 ();
 FILLCELL_X32 FILLER_97_2000 ();
 FILLCELL_X32 FILLER_97_2032 ();
 FILLCELL_X32 FILLER_97_2064 ();
 FILLCELL_X32 FILLER_97_2096 ();
 FILLCELL_X32 FILLER_97_2128 ();
 FILLCELL_X32 FILLER_97_2160 ();
 FILLCELL_X32 FILLER_97_2192 ();
 FILLCELL_X32 FILLER_97_2224 ();
 FILLCELL_X32 FILLER_97_2256 ();
 FILLCELL_X32 FILLER_97_2288 ();
 FILLCELL_X32 FILLER_97_2320 ();
 FILLCELL_X32 FILLER_97_2352 ();
 FILLCELL_X32 FILLER_97_2384 ();
 FILLCELL_X16 FILLER_97_2416 ();
 FILLCELL_X4 FILLER_97_2432 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X32 FILLER_98_1784 ();
 FILLCELL_X32 FILLER_98_1816 ();
 FILLCELL_X32 FILLER_98_1848 ();
 FILLCELL_X8 FILLER_98_1880 ();
 FILLCELL_X4 FILLER_98_1888 ();
 FILLCELL_X2 FILLER_98_1892 ();
 FILLCELL_X32 FILLER_98_1895 ();
 FILLCELL_X32 FILLER_98_1927 ();
 FILLCELL_X32 FILLER_98_1959 ();
 FILLCELL_X32 FILLER_98_1991 ();
 FILLCELL_X32 FILLER_98_2023 ();
 FILLCELL_X32 FILLER_98_2055 ();
 FILLCELL_X32 FILLER_98_2087 ();
 FILLCELL_X32 FILLER_98_2119 ();
 FILLCELL_X32 FILLER_98_2151 ();
 FILLCELL_X32 FILLER_98_2183 ();
 FILLCELL_X32 FILLER_98_2215 ();
 FILLCELL_X32 FILLER_98_2247 ();
 FILLCELL_X32 FILLER_98_2279 ();
 FILLCELL_X32 FILLER_98_2311 ();
 FILLCELL_X32 FILLER_98_2343 ();
 FILLCELL_X32 FILLER_98_2375 ();
 FILLCELL_X16 FILLER_98_2407 ();
 FILLCELL_X8 FILLER_98_2423 ();
 FILLCELL_X4 FILLER_98_2431 ();
 FILLCELL_X1 FILLER_98_2435 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X32 FILLER_99_1776 ();
 FILLCELL_X32 FILLER_99_1808 ();
 FILLCELL_X32 FILLER_99_1840 ();
 FILLCELL_X32 FILLER_99_1872 ();
 FILLCELL_X32 FILLER_99_1904 ();
 FILLCELL_X32 FILLER_99_1936 ();
 FILLCELL_X32 FILLER_99_1968 ();
 FILLCELL_X32 FILLER_99_2000 ();
 FILLCELL_X32 FILLER_99_2032 ();
 FILLCELL_X32 FILLER_99_2064 ();
 FILLCELL_X32 FILLER_99_2096 ();
 FILLCELL_X32 FILLER_99_2128 ();
 FILLCELL_X32 FILLER_99_2160 ();
 FILLCELL_X32 FILLER_99_2192 ();
 FILLCELL_X32 FILLER_99_2224 ();
 FILLCELL_X32 FILLER_99_2256 ();
 FILLCELL_X32 FILLER_99_2288 ();
 FILLCELL_X32 FILLER_99_2320 ();
 FILLCELL_X32 FILLER_99_2352 ();
 FILLCELL_X32 FILLER_99_2384 ();
 FILLCELL_X16 FILLER_99_2416 ();
 FILLCELL_X4 FILLER_99_2432 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X32 FILLER_100_1784 ();
 FILLCELL_X32 FILLER_100_1816 ();
 FILLCELL_X32 FILLER_100_1848 ();
 FILLCELL_X8 FILLER_100_1880 ();
 FILLCELL_X4 FILLER_100_1888 ();
 FILLCELL_X2 FILLER_100_1892 ();
 FILLCELL_X32 FILLER_100_1895 ();
 FILLCELL_X32 FILLER_100_1927 ();
 FILLCELL_X32 FILLER_100_1959 ();
 FILLCELL_X32 FILLER_100_1991 ();
 FILLCELL_X32 FILLER_100_2023 ();
 FILLCELL_X32 FILLER_100_2055 ();
 FILLCELL_X32 FILLER_100_2087 ();
 FILLCELL_X32 FILLER_100_2119 ();
 FILLCELL_X32 FILLER_100_2151 ();
 FILLCELL_X32 FILLER_100_2183 ();
 FILLCELL_X32 FILLER_100_2215 ();
 FILLCELL_X32 FILLER_100_2247 ();
 FILLCELL_X32 FILLER_100_2279 ();
 FILLCELL_X32 FILLER_100_2311 ();
 FILLCELL_X32 FILLER_100_2343 ();
 FILLCELL_X32 FILLER_100_2375 ();
 FILLCELL_X16 FILLER_100_2407 ();
 FILLCELL_X8 FILLER_100_2423 ();
 FILLCELL_X4 FILLER_100_2431 ();
 FILLCELL_X1 FILLER_100_2435 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X32 FILLER_101_1776 ();
 FILLCELL_X32 FILLER_101_1808 ();
 FILLCELL_X32 FILLER_101_1840 ();
 FILLCELL_X32 FILLER_101_1872 ();
 FILLCELL_X32 FILLER_101_1904 ();
 FILLCELL_X32 FILLER_101_1936 ();
 FILLCELL_X32 FILLER_101_1968 ();
 FILLCELL_X32 FILLER_101_2000 ();
 FILLCELL_X32 FILLER_101_2032 ();
 FILLCELL_X32 FILLER_101_2064 ();
 FILLCELL_X32 FILLER_101_2096 ();
 FILLCELL_X32 FILLER_101_2128 ();
 FILLCELL_X32 FILLER_101_2160 ();
 FILLCELL_X32 FILLER_101_2192 ();
 FILLCELL_X32 FILLER_101_2224 ();
 FILLCELL_X32 FILLER_101_2256 ();
 FILLCELL_X32 FILLER_101_2288 ();
 FILLCELL_X32 FILLER_101_2320 ();
 FILLCELL_X32 FILLER_101_2352 ();
 FILLCELL_X32 FILLER_101_2384 ();
 FILLCELL_X16 FILLER_101_2416 ();
 FILLCELL_X4 FILLER_101_2432 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X32 FILLER_102_1784 ();
 FILLCELL_X32 FILLER_102_1816 ();
 FILLCELL_X32 FILLER_102_1848 ();
 FILLCELL_X8 FILLER_102_1880 ();
 FILLCELL_X4 FILLER_102_1888 ();
 FILLCELL_X2 FILLER_102_1892 ();
 FILLCELL_X32 FILLER_102_1895 ();
 FILLCELL_X32 FILLER_102_1927 ();
 FILLCELL_X32 FILLER_102_1959 ();
 FILLCELL_X32 FILLER_102_1991 ();
 FILLCELL_X32 FILLER_102_2023 ();
 FILLCELL_X32 FILLER_102_2055 ();
 FILLCELL_X32 FILLER_102_2087 ();
 FILLCELL_X32 FILLER_102_2119 ();
 FILLCELL_X32 FILLER_102_2151 ();
 FILLCELL_X32 FILLER_102_2183 ();
 FILLCELL_X32 FILLER_102_2215 ();
 FILLCELL_X32 FILLER_102_2247 ();
 FILLCELL_X32 FILLER_102_2279 ();
 FILLCELL_X32 FILLER_102_2311 ();
 FILLCELL_X32 FILLER_102_2343 ();
 FILLCELL_X32 FILLER_102_2375 ();
 FILLCELL_X16 FILLER_102_2407 ();
 FILLCELL_X8 FILLER_102_2423 ();
 FILLCELL_X4 FILLER_102_2431 ();
 FILLCELL_X1 FILLER_102_2435 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X32 FILLER_103_1776 ();
 FILLCELL_X32 FILLER_103_1808 ();
 FILLCELL_X32 FILLER_103_1840 ();
 FILLCELL_X32 FILLER_103_1872 ();
 FILLCELL_X32 FILLER_103_1904 ();
 FILLCELL_X32 FILLER_103_1936 ();
 FILLCELL_X32 FILLER_103_1968 ();
 FILLCELL_X32 FILLER_103_2000 ();
 FILLCELL_X32 FILLER_103_2032 ();
 FILLCELL_X32 FILLER_103_2064 ();
 FILLCELL_X32 FILLER_103_2096 ();
 FILLCELL_X32 FILLER_103_2128 ();
 FILLCELL_X32 FILLER_103_2160 ();
 FILLCELL_X32 FILLER_103_2192 ();
 FILLCELL_X32 FILLER_103_2224 ();
 FILLCELL_X32 FILLER_103_2256 ();
 FILLCELL_X32 FILLER_103_2288 ();
 FILLCELL_X32 FILLER_103_2320 ();
 FILLCELL_X32 FILLER_103_2352 ();
 FILLCELL_X32 FILLER_103_2384 ();
 FILLCELL_X16 FILLER_103_2416 ();
 FILLCELL_X4 FILLER_103_2432 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X32 FILLER_104_1784 ();
 FILLCELL_X32 FILLER_104_1816 ();
 FILLCELL_X32 FILLER_104_1848 ();
 FILLCELL_X8 FILLER_104_1880 ();
 FILLCELL_X4 FILLER_104_1888 ();
 FILLCELL_X2 FILLER_104_1892 ();
 FILLCELL_X32 FILLER_104_1895 ();
 FILLCELL_X32 FILLER_104_1927 ();
 FILLCELL_X32 FILLER_104_1959 ();
 FILLCELL_X32 FILLER_104_1991 ();
 FILLCELL_X32 FILLER_104_2023 ();
 FILLCELL_X32 FILLER_104_2055 ();
 FILLCELL_X32 FILLER_104_2087 ();
 FILLCELL_X32 FILLER_104_2119 ();
 FILLCELL_X32 FILLER_104_2151 ();
 FILLCELL_X32 FILLER_104_2183 ();
 FILLCELL_X32 FILLER_104_2215 ();
 FILLCELL_X32 FILLER_104_2247 ();
 FILLCELL_X32 FILLER_104_2279 ();
 FILLCELL_X32 FILLER_104_2311 ();
 FILLCELL_X32 FILLER_104_2343 ();
 FILLCELL_X32 FILLER_104_2375 ();
 FILLCELL_X16 FILLER_104_2407 ();
 FILLCELL_X8 FILLER_104_2423 ();
 FILLCELL_X4 FILLER_104_2431 ();
 FILLCELL_X1 FILLER_104_2435 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X32 FILLER_105_1776 ();
 FILLCELL_X32 FILLER_105_1808 ();
 FILLCELL_X32 FILLER_105_1840 ();
 FILLCELL_X32 FILLER_105_1872 ();
 FILLCELL_X32 FILLER_105_1904 ();
 FILLCELL_X32 FILLER_105_1936 ();
 FILLCELL_X32 FILLER_105_1968 ();
 FILLCELL_X32 FILLER_105_2000 ();
 FILLCELL_X32 FILLER_105_2032 ();
 FILLCELL_X32 FILLER_105_2064 ();
 FILLCELL_X32 FILLER_105_2096 ();
 FILLCELL_X32 FILLER_105_2128 ();
 FILLCELL_X32 FILLER_105_2160 ();
 FILLCELL_X32 FILLER_105_2192 ();
 FILLCELL_X32 FILLER_105_2224 ();
 FILLCELL_X32 FILLER_105_2256 ();
 FILLCELL_X32 FILLER_105_2288 ();
 FILLCELL_X32 FILLER_105_2320 ();
 FILLCELL_X32 FILLER_105_2352 ();
 FILLCELL_X32 FILLER_105_2384 ();
 FILLCELL_X16 FILLER_105_2416 ();
 FILLCELL_X4 FILLER_105_2432 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_106_1784 ();
 FILLCELL_X32 FILLER_106_1816 ();
 FILLCELL_X32 FILLER_106_1848 ();
 FILLCELL_X8 FILLER_106_1880 ();
 FILLCELL_X4 FILLER_106_1888 ();
 FILLCELL_X2 FILLER_106_1892 ();
 FILLCELL_X32 FILLER_106_1895 ();
 FILLCELL_X32 FILLER_106_1927 ();
 FILLCELL_X32 FILLER_106_1959 ();
 FILLCELL_X32 FILLER_106_1991 ();
 FILLCELL_X32 FILLER_106_2023 ();
 FILLCELL_X32 FILLER_106_2055 ();
 FILLCELL_X32 FILLER_106_2087 ();
 FILLCELL_X32 FILLER_106_2119 ();
 FILLCELL_X32 FILLER_106_2151 ();
 FILLCELL_X32 FILLER_106_2183 ();
 FILLCELL_X32 FILLER_106_2215 ();
 FILLCELL_X32 FILLER_106_2247 ();
 FILLCELL_X32 FILLER_106_2279 ();
 FILLCELL_X32 FILLER_106_2311 ();
 FILLCELL_X32 FILLER_106_2343 ();
 FILLCELL_X32 FILLER_106_2375 ();
 FILLCELL_X16 FILLER_106_2407 ();
 FILLCELL_X8 FILLER_106_2423 ();
 FILLCELL_X4 FILLER_106_2431 ();
 FILLCELL_X1 FILLER_106_2435 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X32 FILLER_107_1776 ();
 FILLCELL_X32 FILLER_107_1808 ();
 FILLCELL_X32 FILLER_107_1840 ();
 FILLCELL_X32 FILLER_107_1872 ();
 FILLCELL_X32 FILLER_107_1904 ();
 FILLCELL_X32 FILLER_107_1936 ();
 FILLCELL_X32 FILLER_107_1968 ();
 FILLCELL_X32 FILLER_107_2000 ();
 FILLCELL_X32 FILLER_107_2032 ();
 FILLCELL_X32 FILLER_107_2064 ();
 FILLCELL_X32 FILLER_107_2096 ();
 FILLCELL_X32 FILLER_107_2128 ();
 FILLCELL_X32 FILLER_107_2160 ();
 FILLCELL_X32 FILLER_107_2192 ();
 FILLCELL_X32 FILLER_107_2224 ();
 FILLCELL_X32 FILLER_107_2256 ();
 FILLCELL_X32 FILLER_107_2288 ();
 FILLCELL_X32 FILLER_107_2320 ();
 FILLCELL_X32 FILLER_107_2352 ();
 FILLCELL_X32 FILLER_107_2384 ();
 FILLCELL_X16 FILLER_107_2416 ();
 FILLCELL_X4 FILLER_107_2432 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X32 FILLER_108_952 ();
 FILLCELL_X32 FILLER_108_984 ();
 FILLCELL_X32 FILLER_108_1016 ();
 FILLCELL_X32 FILLER_108_1048 ();
 FILLCELL_X32 FILLER_108_1080 ();
 FILLCELL_X32 FILLER_108_1112 ();
 FILLCELL_X32 FILLER_108_1144 ();
 FILLCELL_X32 FILLER_108_1176 ();
 FILLCELL_X32 FILLER_108_1208 ();
 FILLCELL_X32 FILLER_108_1240 ();
 FILLCELL_X32 FILLER_108_1272 ();
 FILLCELL_X32 FILLER_108_1304 ();
 FILLCELL_X32 FILLER_108_1336 ();
 FILLCELL_X32 FILLER_108_1368 ();
 FILLCELL_X32 FILLER_108_1400 ();
 FILLCELL_X32 FILLER_108_1432 ();
 FILLCELL_X32 FILLER_108_1464 ();
 FILLCELL_X32 FILLER_108_1496 ();
 FILLCELL_X32 FILLER_108_1528 ();
 FILLCELL_X32 FILLER_108_1560 ();
 FILLCELL_X32 FILLER_108_1592 ();
 FILLCELL_X32 FILLER_108_1624 ();
 FILLCELL_X32 FILLER_108_1656 ();
 FILLCELL_X32 FILLER_108_1688 ();
 FILLCELL_X32 FILLER_108_1720 ();
 FILLCELL_X32 FILLER_108_1752 ();
 FILLCELL_X32 FILLER_108_1784 ();
 FILLCELL_X32 FILLER_108_1816 ();
 FILLCELL_X32 FILLER_108_1848 ();
 FILLCELL_X8 FILLER_108_1880 ();
 FILLCELL_X4 FILLER_108_1888 ();
 FILLCELL_X2 FILLER_108_1892 ();
 FILLCELL_X32 FILLER_108_1895 ();
 FILLCELL_X32 FILLER_108_1927 ();
 FILLCELL_X32 FILLER_108_1959 ();
 FILLCELL_X32 FILLER_108_1991 ();
 FILLCELL_X32 FILLER_108_2023 ();
 FILLCELL_X32 FILLER_108_2055 ();
 FILLCELL_X32 FILLER_108_2087 ();
 FILLCELL_X32 FILLER_108_2119 ();
 FILLCELL_X32 FILLER_108_2151 ();
 FILLCELL_X32 FILLER_108_2183 ();
 FILLCELL_X32 FILLER_108_2215 ();
 FILLCELL_X32 FILLER_108_2247 ();
 FILLCELL_X32 FILLER_108_2279 ();
 FILLCELL_X32 FILLER_108_2311 ();
 FILLCELL_X32 FILLER_108_2343 ();
 FILLCELL_X32 FILLER_108_2375 ();
 FILLCELL_X16 FILLER_108_2407 ();
 FILLCELL_X8 FILLER_108_2423 ();
 FILLCELL_X4 FILLER_108_2431 ();
 FILLCELL_X1 FILLER_108_2435 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X32 FILLER_109_1712 ();
 FILLCELL_X32 FILLER_109_1744 ();
 FILLCELL_X32 FILLER_109_1776 ();
 FILLCELL_X32 FILLER_109_1808 ();
 FILLCELL_X32 FILLER_109_1840 ();
 FILLCELL_X32 FILLER_109_1872 ();
 FILLCELL_X32 FILLER_109_1904 ();
 FILLCELL_X32 FILLER_109_1936 ();
 FILLCELL_X32 FILLER_109_1968 ();
 FILLCELL_X32 FILLER_109_2000 ();
 FILLCELL_X32 FILLER_109_2032 ();
 FILLCELL_X32 FILLER_109_2064 ();
 FILLCELL_X32 FILLER_109_2096 ();
 FILLCELL_X32 FILLER_109_2128 ();
 FILLCELL_X32 FILLER_109_2160 ();
 FILLCELL_X32 FILLER_109_2192 ();
 FILLCELL_X32 FILLER_109_2224 ();
 FILLCELL_X32 FILLER_109_2256 ();
 FILLCELL_X32 FILLER_109_2288 ();
 FILLCELL_X32 FILLER_109_2320 ();
 FILLCELL_X32 FILLER_109_2352 ();
 FILLCELL_X32 FILLER_109_2384 ();
 FILLCELL_X16 FILLER_109_2416 ();
 FILLCELL_X4 FILLER_109_2432 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X32 FILLER_110_1304 ();
 FILLCELL_X32 FILLER_110_1336 ();
 FILLCELL_X32 FILLER_110_1368 ();
 FILLCELL_X32 FILLER_110_1400 ();
 FILLCELL_X32 FILLER_110_1432 ();
 FILLCELL_X32 FILLER_110_1464 ();
 FILLCELL_X32 FILLER_110_1496 ();
 FILLCELL_X32 FILLER_110_1528 ();
 FILLCELL_X32 FILLER_110_1560 ();
 FILLCELL_X32 FILLER_110_1592 ();
 FILLCELL_X32 FILLER_110_1624 ();
 FILLCELL_X32 FILLER_110_1656 ();
 FILLCELL_X32 FILLER_110_1688 ();
 FILLCELL_X32 FILLER_110_1720 ();
 FILLCELL_X32 FILLER_110_1752 ();
 FILLCELL_X32 FILLER_110_1784 ();
 FILLCELL_X32 FILLER_110_1816 ();
 FILLCELL_X32 FILLER_110_1848 ();
 FILLCELL_X8 FILLER_110_1880 ();
 FILLCELL_X4 FILLER_110_1888 ();
 FILLCELL_X2 FILLER_110_1892 ();
 FILLCELL_X32 FILLER_110_1895 ();
 FILLCELL_X32 FILLER_110_1927 ();
 FILLCELL_X32 FILLER_110_1959 ();
 FILLCELL_X32 FILLER_110_1991 ();
 FILLCELL_X32 FILLER_110_2023 ();
 FILLCELL_X32 FILLER_110_2055 ();
 FILLCELL_X32 FILLER_110_2087 ();
 FILLCELL_X32 FILLER_110_2119 ();
 FILLCELL_X32 FILLER_110_2151 ();
 FILLCELL_X32 FILLER_110_2183 ();
 FILLCELL_X32 FILLER_110_2215 ();
 FILLCELL_X32 FILLER_110_2247 ();
 FILLCELL_X32 FILLER_110_2279 ();
 FILLCELL_X32 FILLER_110_2311 ();
 FILLCELL_X32 FILLER_110_2343 ();
 FILLCELL_X32 FILLER_110_2375 ();
 FILLCELL_X16 FILLER_110_2407 ();
 FILLCELL_X8 FILLER_110_2423 ();
 FILLCELL_X4 FILLER_110_2431 ();
 FILLCELL_X1 FILLER_110_2435 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X32 FILLER_111_1712 ();
 FILLCELL_X32 FILLER_111_1744 ();
 FILLCELL_X32 FILLER_111_1776 ();
 FILLCELL_X32 FILLER_111_1808 ();
 FILLCELL_X32 FILLER_111_1840 ();
 FILLCELL_X32 FILLER_111_1872 ();
 FILLCELL_X32 FILLER_111_1904 ();
 FILLCELL_X32 FILLER_111_1936 ();
 FILLCELL_X32 FILLER_111_1968 ();
 FILLCELL_X32 FILLER_111_2000 ();
 FILLCELL_X32 FILLER_111_2032 ();
 FILLCELL_X32 FILLER_111_2064 ();
 FILLCELL_X32 FILLER_111_2096 ();
 FILLCELL_X32 FILLER_111_2128 ();
 FILLCELL_X32 FILLER_111_2160 ();
 FILLCELL_X32 FILLER_111_2192 ();
 FILLCELL_X32 FILLER_111_2224 ();
 FILLCELL_X32 FILLER_111_2256 ();
 FILLCELL_X32 FILLER_111_2288 ();
 FILLCELL_X32 FILLER_111_2320 ();
 FILLCELL_X32 FILLER_111_2352 ();
 FILLCELL_X32 FILLER_111_2384 ();
 FILLCELL_X16 FILLER_111_2416 ();
 FILLCELL_X4 FILLER_111_2432 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X32 FILLER_112_1272 ();
 FILLCELL_X32 FILLER_112_1304 ();
 FILLCELL_X32 FILLER_112_1336 ();
 FILLCELL_X32 FILLER_112_1368 ();
 FILLCELL_X32 FILLER_112_1400 ();
 FILLCELL_X32 FILLER_112_1432 ();
 FILLCELL_X32 FILLER_112_1464 ();
 FILLCELL_X32 FILLER_112_1496 ();
 FILLCELL_X32 FILLER_112_1528 ();
 FILLCELL_X32 FILLER_112_1560 ();
 FILLCELL_X32 FILLER_112_1592 ();
 FILLCELL_X32 FILLER_112_1624 ();
 FILLCELL_X32 FILLER_112_1656 ();
 FILLCELL_X32 FILLER_112_1688 ();
 FILLCELL_X32 FILLER_112_1720 ();
 FILLCELL_X32 FILLER_112_1752 ();
 FILLCELL_X32 FILLER_112_1784 ();
 FILLCELL_X32 FILLER_112_1816 ();
 FILLCELL_X32 FILLER_112_1848 ();
 FILLCELL_X8 FILLER_112_1880 ();
 FILLCELL_X4 FILLER_112_1888 ();
 FILLCELL_X2 FILLER_112_1892 ();
 FILLCELL_X32 FILLER_112_1895 ();
 FILLCELL_X32 FILLER_112_1927 ();
 FILLCELL_X32 FILLER_112_1959 ();
 FILLCELL_X32 FILLER_112_1991 ();
 FILLCELL_X32 FILLER_112_2023 ();
 FILLCELL_X32 FILLER_112_2055 ();
 FILLCELL_X32 FILLER_112_2087 ();
 FILLCELL_X32 FILLER_112_2119 ();
 FILLCELL_X32 FILLER_112_2151 ();
 FILLCELL_X32 FILLER_112_2183 ();
 FILLCELL_X32 FILLER_112_2215 ();
 FILLCELL_X32 FILLER_112_2247 ();
 FILLCELL_X32 FILLER_112_2279 ();
 FILLCELL_X32 FILLER_112_2311 ();
 FILLCELL_X32 FILLER_112_2343 ();
 FILLCELL_X32 FILLER_112_2375 ();
 FILLCELL_X16 FILLER_112_2407 ();
 FILLCELL_X8 FILLER_112_2423 ();
 FILLCELL_X4 FILLER_112_2431 ();
 FILLCELL_X1 FILLER_112_2435 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X32 FILLER_113_865 ();
 FILLCELL_X32 FILLER_113_897 ();
 FILLCELL_X32 FILLER_113_929 ();
 FILLCELL_X32 FILLER_113_961 ();
 FILLCELL_X32 FILLER_113_993 ();
 FILLCELL_X32 FILLER_113_1025 ();
 FILLCELL_X32 FILLER_113_1057 ();
 FILLCELL_X32 FILLER_113_1089 ();
 FILLCELL_X32 FILLER_113_1121 ();
 FILLCELL_X32 FILLER_113_1153 ();
 FILLCELL_X32 FILLER_113_1185 ();
 FILLCELL_X32 FILLER_113_1217 ();
 FILLCELL_X8 FILLER_113_1249 ();
 FILLCELL_X4 FILLER_113_1257 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X32 FILLER_113_1712 ();
 FILLCELL_X32 FILLER_113_1744 ();
 FILLCELL_X32 FILLER_113_1776 ();
 FILLCELL_X32 FILLER_113_1808 ();
 FILLCELL_X32 FILLER_113_1840 ();
 FILLCELL_X32 FILLER_113_1872 ();
 FILLCELL_X32 FILLER_113_1904 ();
 FILLCELL_X32 FILLER_113_1936 ();
 FILLCELL_X32 FILLER_113_1968 ();
 FILLCELL_X32 FILLER_113_2000 ();
 FILLCELL_X32 FILLER_113_2032 ();
 FILLCELL_X32 FILLER_113_2064 ();
 FILLCELL_X32 FILLER_113_2096 ();
 FILLCELL_X32 FILLER_113_2128 ();
 FILLCELL_X32 FILLER_113_2160 ();
 FILLCELL_X32 FILLER_113_2192 ();
 FILLCELL_X32 FILLER_113_2224 ();
 FILLCELL_X32 FILLER_113_2256 ();
 FILLCELL_X32 FILLER_113_2288 ();
 FILLCELL_X32 FILLER_113_2320 ();
 FILLCELL_X32 FILLER_113_2352 ();
 FILLCELL_X32 FILLER_113_2384 ();
 FILLCELL_X16 FILLER_113_2416 ();
 FILLCELL_X4 FILLER_113_2432 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X32 FILLER_114_1176 ();
 FILLCELL_X32 FILLER_114_1208 ();
 FILLCELL_X32 FILLER_114_1240 ();
 FILLCELL_X32 FILLER_114_1272 ();
 FILLCELL_X32 FILLER_114_1304 ();
 FILLCELL_X32 FILLER_114_1336 ();
 FILLCELL_X32 FILLER_114_1368 ();
 FILLCELL_X32 FILLER_114_1400 ();
 FILLCELL_X32 FILLER_114_1432 ();
 FILLCELL_X32 FILLER_114_1464 ();
 FILLCELL_X32 FILLER_114_1496 ();
 FILLCELL_X32 FILLER_114_1528 ();
 FILLCELL_X32 FILLER_114_1560 ();
 FILLCELL_X32 FILLER_114_1592 ();
 FILLCELL_X32 FILLER_114_1624 ();
 FILLCELL_X32 FILLER_114_1656 ();
 FILLCELL_X32 FILLER_114_1688 ();
 FILLCELL_X32 FILLER_114_1720 ();
 FILLCELL_X32 FILLER_114_1752 ();
 FILLCELL_X32 FILLER_114_1784 ();
 FILLCELL_X32 FILLER_114_1816 ();
 FILLCELL_X32 FILLER_114_1848 ();
 FILLCELL_X8 FILLER_114_1880 ();
 FILLCELL_X4 FILLER_114_1888 ();
 FILLCELL_X2 FILLER_114_1892 ();
 FILLCELL_X32 FILLER_114_1895 ();
 FILLCELL_X32 FILLER_114_1927 ();
 FILLCELL_X32 FILLER_114_1959 ();
 FILLCELL_X32 FILLER_114_1991 ();
 FILLCELL_X32 FILLER_114_2023 ();
 FILLCELL_X32 FILLER_114_2055 ();
 FILLCELL_X32 FILLER_114_2087 ();
 FILLCELL_X32 FILLER_114_2119 ();
 FILLCELL_X32 FILLER_114_2151 ();
 FILLCELL_X32 FILLER_114_2183 ();
 FILLCELL_X32 FILLER_114_2215 ();
 FILLCELL_X32 FILLER_114_2247 ();
 FILLCELL_X32 FILLER_114_2279 ();
 FILLCELL_X32 FILLER_114_2311 ();
 FILLCELL_X32 FILLER_114_2343 ();
 FILLCELL_X32 FILLER_114_2375 ();
 FILLCELL_X16 FILLER_114_2407 ();
 FILLCELL_X8 FILLER_114_2423 ();
 FILLCELL_X4 FILLER_114_2431 ();
 FILLCELL_X1 FILLER_114_2435 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X32 FILLER_115_961 ();
 FILLCELL_X32 FILLER_115_993 ();
 FILLCELL_X32 FILLER_115_1025 ();
 FILLCELL_X32 FILLER_115_1057 ();
 FILLCELL_X32 FILLER_115_1089 ();
 FILLCELL_X32 FILLER_115_1121 ();
 FILLCELL_X32 FILLER_115_1153 ();
 FILLCELL_X32 FILLER_115_1185 ();
 FILLCELL_X32 FILLER_115_1217 ();
 FILLCELL_X8 FILLER_115_1249 ();
 FILLCELL_X4 FILLER_115_1257 ();
 FILLCELL_X2 FILLER_115_1261 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X32 FILLER_115_1744 ();
 FILLCELL_X32 FILLER_115_1776 ();
 FILLCELL_X32 FILLER_115_1808 ();
 FILLCELL_X32 FILLER_115_1840 ();
 FILLCELL_X32 FILLER_115_1872 ();
 FILLCELL_X32 FILLER_115_1904 ();
 FILLCELL_X32 FILLER_115_1936 ();
 FILLCELL_X32 FILLER_115_1968 ();
 FILLCELL_X32 FILLER_115_2000 ();
 FILLCELL_X32 FILLER_115_2032 ();
 FILLCELL_X32 FILLER_115_2064 ();
 FILLCELL_X32 FILLER_115_2096 ();
 FILLCELL_X32 FILLER_115_2128 ();
 FILLCELL_X32 FILLER_115_2160 ();
 FILLCELL_X32 FILLER_115_2192 ();
 FILLCELL_X32 FILLER_115_2224 ();
 FILLCELL_X32 FILLER_115_2256 ();
 FILLCELL_X32 FILLER_115_2288 ();
 FILLCELL_X32 FILLER_115_2320 ();
 FILLCELL_X32 FILLER_115_2352 ();
 FILLCELL_X32 FILLER_115_2384 ();
 FILLCELL_X16 FILLER_115_2416 ();
 FILLCELL_X4 FILLER_115_2432 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X32 FILLER_116_952 ();
 FILLCELL_X32 FILLER_116_984 ();
 FILLCELL_X32 FILLER_116_1016 ();
 FILLCELL_X32 FILLER_116_1048 ();
 FILLCELL_X32 FILLER_116_1080 ();
 FILLCELL_X32 FILLER_116_1112 ();
 FILLCELL_X32 FILLER_116_1144 ();
 FILLCELL_X32 FILLER_116_1176 ();
 FILLCELL_X32 FILLER_116_1208 ();
 FILLCELL_X32 FILLER_116_1240 ();
 FILLCELL_X32 FILLER_116_1272 ();
 FILLCELL_X32 FILLER_116_1304 ();
 FILLCELL_X32 FILLER_116_1336 ();
 FILLCELL_X32 FILLER_116_1368 ();
 FILLCELL_X32 FILLER_116_1400 ();
 FILLCELL_X32 FILLER_116_1432 ();
 FILLCELL_X32 FILLER_116_1464 ();
 FILLCELL_X32 FILLER_116_1496 ();
 FILLCELL_X32 FILLER_116_1528 ();
 FILLCELL_X32 FILLER_116_1560 ();
 FILLCELL_X32 FILLER_116_1592 ();
 FILLCELL_X32 FILLER_116_1624 ();
 FILLCELL_X32 FILLER_116_1656 ();
 FILLCELL_X32 FILLER_116_1688 ();
 FILLCELL_X32 FILLER_116_1720 ();
 FILLCELL_X32 FILLER_116_1752 ();
 FILLCELL_X32 FILLER_116_1784 ();
 FILLCELL_X32 FILLER_116_1816 ();
 FILLCELL_X32 FILLER_116_1848 ();
 FILLCELL_X8 FILLER_116_1880 ();
 FILLCELL_X4 FILLER_116_1888 ();
 FILLCELL_X2 FILLER_116_1892 ();
 FILLCELL_X32 FILLER_116_1895 ();
 FILLCELL_X32 FILLER_116_1927 ();
 FILLCELL_X32 FILLER_116_1959 ();
 FILLCELL_X32 FILLER_116_1991 ();
 FILLCELL_X32 FILLER_116_2023 ();
 FILLCELL_X32 FILLER_116_2055 ();
 FILLCELL_X32 FILLER_116_2087 ();
 FILLCELL_X32 FILLER_116_2119 ();
 FILLCELL_X32 FILLER_116_2151 ();
 FILLCELL_X32 FILLER_116_2183 ();
 FILLCELL_X32 FILLER_116_2215 ();
 FILLCELL_X32 FILLER_116_2247 ();
 FILLCELL_X32 FILLER_116_2279 ();
 FILLCELL_X32 FILLER_116_2311 ();
 FILLCELL_X32 FILLER_116_2343 ();
 FILLCELL_X32 FILLER_116_2375 ();
 FILLCELL_X16 FILLER_116_2407 ();
 FILLCELL_X8 FILLER_116_2423 ();
 FILLCELL_X4 FILLER_116_2431 ();
 FILLCELL_X1 FILLER_116_2435 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X32 FILLER_117_961 ();
 FILLCELL_X32 FILLER_117_993 ();
 FILLCELL_X32 FILLER_117_1025 ();
 FILLCELL_X32 FILLER_117_1057 ();
 FILLCELL_X32 FILLER_117_1089 ();
 FILLCELL_X32 FILLER_117_1121 ();
 FILLCELL_X32 FILLER_117_1153 ();
 FILLCELL_X32 FILLER_117_1185 ();
 FILLCELL_X32 FILLER_117_1217 ();
 FILLCELL_X8 FILLER_117_1249 ();
 FILLCELL_X4 FILLER_117_1257 ();
 FILLCELL_X2 FILLER_117_1261 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X32 FILLER_117_1744 ();
 FILLCELL_X32 FILLER_117_1776 ();
 FILLCELL_X32 FILLER_117_1808 ();
 FILLCELL_X32 FILLER_117_1840 ();
 FILLCELL_X32 FILLER_117_1872 ();
 FILLCELL_X32 FILLER_117_1904 ();
 FILLCELL_X32 FILLER_117_1936 ();
 FILLCELL_X32 FILLER_117_1968 ();
 FILLCELL_X32 FILLER_117_2000 ();
 FILLCELL_X32 FILLER_117_2032 ();
 FILLCELL_X32 FILLER_117_2064 ();
 FILLCELL_X32 FILLER_117_2096 ();
 FILLCELL_X32 FILLER_117_2128 ();
 FILLCELL_X32 FILLER_117_2160 ();
 FILLCELL_X32 FILLER_117_2192 ();
 FILLCELL_X32 FILLER_117_2224 ();
 FILLCELL_X32 FILLER_117_2256 ();
 FILLCELL_X32 FILLER_117_2288 ();
 FILLCELL_X32 FILLER_117_2320 ();
 FILLCELL_X32 FILLER_117_2352 ();
 FILLCELL_X32 FILLER_117_2384 ();
 FILLCELL_X16 FILLER_117_2416 ();
 FILLCELL_X4 FILLER_117_2432 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X32 FILLER_118_1016 ();
 FILLCELL_X32 FILLER_118_1048 ();
 FILLCELL_X32 FILLER_118_1080 ();
 FILLCELL_X32 FILLER_118_1112 ();
 FILLCELL_X32 FILLER_118_1144 ();
 FILLCELL_X32 FILLER_118_1176 ();
 FILLCELL_X32 FILLER_118_1208 ();
 FILLCELL_X32 FILLER_118_1240 ();
 FILLCELL_X32 FILLER_118_1272 ();
 FILLCELL_X32 FILLER_118_1304 ();
 FILLCELL_X32 FILLER_118_1336 ();
 FILLCELL_X32 FILLER_118_1368 ();
 FILLCELL_X32 FILLER_118_1400 ();
 FILLCELL_X32 FILLER_118_1432 ();
 FILLCELL_X32 FILLER_118_1464 ();
 FILLCELL_X32 FILLER_118_1496 ();
 FILLCELL_X32 FILLER_118_1528 ();
 FILLCELL_X32 FILLER_118_1560 ();
 FILLCELL_X32 FILLER_118_1592 ();
 FILLCELL_X32 FILLER_118_1624 ();
 FILLCELL_X32 FILLER_118_1656 ();
 FILLCELL_X32 FILLER_118_1688 ();
 FILLCELL_X32 FILLER_118_1720 ();
 FILLCELL_X32 FILLER_118_1752 ();
 FILLCELL_X32 FILLER_118_1784 ();
 FILLCELL_X32 FILLER_118_1816 ();
 FILLCELL_X32 FILLER_118_1848 ();
 FILLCELL_X8 FILLER_118_1880 ();
 FILLCELL_X4 FILLER_118_1888 ();
 FILLCELL_X2 FILLER_118_1892 ();
 FILLCELL_X32 FILLER_118_1895 ();
 FILLCELL_X32 FILLER_118_1927 ();
 FILLCELL_X32 FILLER_118_1959 ();
 FILLCELL_X32 FILLER_118_1991 ();
 FILLCELL_X32 FILLER_118_2023 ();
 FILLCELL_X32 FILLER_118_2055 ();
 FILLCELL_X32 FILLER_118_2087 ();
 FILLCELL_X32 FILLER_118_2119 ();
 FILLCELL_X32 FILLER_118_2151 ();
 FILLCELL_X32 FILLER_118_2183 ();
 FILLCELL_X32 FILLER_118_2215 ();
 FILLCELL_X32 FILLER_118_2247 ();
 FILLCELL_X32 FILLER_118_2279 ();
 FILLCELL_X32 FILLER_118_2311 ();
 FILLCELL_X32 FILLER_118_2343 ();
 FILLCELL_X32 FILLER_118_2375 ();
 FILLCELL_X16 FILLER_118_2407 ();
 FILLCELL_X8 FILLER_118_2423 ();
 FILLCELL_X4 FILLER_118_2431 ();
 FILLCELL_X1 FILLER_118_2435 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X32 FILLER_119_993 ();
 FILLCELL_X32 FILLER_119_1025 ();
 FILLCELL_X32 FILLER_119_1057 ();
 FILLCELL_X32 FILLER_119_1089 ();
 FILLCELL_X32 FILLER_119_1121 ();
 FILLCELL_X32 FILLER_119_1153 ();
 FILLCELL_X32 FILLER_119_1185 ();
 FILLCELL_X32 FILLER_119_1217 ();
 FILLCELL_X8 FILLER_119_1249 ();
 FILLCELL_X4 FILLER_119_1257 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X32 FILLER_119_1712 ();
 FILLCELL_X32 FILLER_119_1744 ();
 FILLCELL_X32 FILLER_119_1776 ();
 FILLCELL_X32 FILLER_119_1808 ();
 FILLCELL_X32 FILLER_119_1840 ();
 FILLCELL_X32 FILLER_119_1872 ();
 FILLCELL_X32 FILLER_119_1904 ();
 FILLCELL_X32 FILLER_119_1936 ();
 FILLCELL_X32 FILLER_119_1968 ();
 FILLCELL_X32 FILLER_119_2000 ();
 FILLCELL_X32 FILLER_119_2032 ();
 FILLCELL_X32 FILLER_119_2064 ();
 FILLCELL_X32 FILLER_119_2096 ();
 FILLCELL_X32 FILLER_119_2128 ();
 FILLCELL_X32 FILLER_119_2160 ();
 FILLCELL_X32 FILLER_119_2192 ();
 FILLCELL_X32 FILLER_119_2224 ();
 FILLCELL_X32 FILLER_119_2256 ();
 FILLCELL_X32 FILLER_119_2288 ();
 FILLCELL_X32 FILLER_119_2320 ();
 FILLCELL_X32 FILLER_119_2352 ();
 FILLCELL_X32 FILLER_119_2384 ();
 FILLCELL_X16 FILLER_119_2416 ();
 FILLCELL_X4 FILLER_119_2432 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X32 FILLER_120_1016 ();
 FILLCELL_X32 FILLER_120_1048 ();
 FILLCELL_X32 FILLER_120_1080 ();
 FILLCELL_X32 FILLER_120_1112 ();
 FILLCELL_X32 FILLER_120_1144 ();
 FILLCELL_X32 FILLER_120_1176 ();
 FILLCELL_X32 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_120_1240 ();
 FILLCELL_X32 FILLER_120_1272 ();
 FILLCELL_X32 FILLER_120_1304 ();
 FILLCELL_X32 FILLER_120_1336 ();
 FILLCELL_X32 FILLER_120_1368 ();
 FILLCELL_X32 FILLER_120_1400 ();
 FILLCELL_X32 FILLER_120_1432 ();
 FILLCELL_X32 FILLER_120_1464 ();
 FILLCELL_X32 FILLER_120_1496 ();
 FILLCELL_X32 FILLER_120_1528 ();
 FILLCELL_X32 FILLER_120_1560 ();
 FILLCELL_X32 FILLER_120_1592 ();
 FILLCELL_X32 FILLER_120_1624 ();
 FILLCELL_X32 FILLER_120_1656 ();
 FILLCELL_X32 FILLER_120_1688 ();
 FILLCELL_X32 FILLER_120_1720 ();
 FILLCELL_X32 FILLER_120_1752 ();
 FILLCELL_X32 FILLER_120_1784 ();
 FILLCELL_X32 FILLER_120_1816 ();
 FILLCELL_X32 FILLER_120_1848 ();
 FILLCELL_X8 FILLER_120_1880 ();
 FILLCELL_X4 FILLER_120_1888 ();
 FILLCELL_X2 FILLER_120_1892 ();
 FILLCELL_X32 FILLER_120_1895 ();
 FILLCELL_X32 FILLER_120_1927 ();
 FILLCELL_X32 FILLER_120_1959 ();
 FILLCELL_X32 FILLER_120_1991 ();
 FILLCELL_X32 FILLER_120_2023 ();
 FILLCELL_X32 FILLER_120_2055 ();
 FILLCELL_X32 FILLER_120_2087 ();
 FILLCELL_X32 FILLER_120_2119 ();
 FILLCELL_X32 FILLER_120_2151 ();
 FILLCELL_X32 FILLER_120_2183 ();
 FILLCELL_X32 FILLER_120_2215 ();
 FILLCELL_X32 FILLER_120_2247 ();
 FILLCELL_X32 FILLER_120_2279 ();
 FILLCELL_X32 FILLER_120_2311 ();
 FILLCELL_X32 FILLER_120_2343 ();
 FILLCELL_X32 FILLER_120_2375 ();
 FILLCELL_X16 FILLER_120_2407 ();
 FILLCELL_X8 FILLER_120_2423 ();
 FILLCELL_X4 FILLER_120_2431 ();
 FILLCELL_X1 FILLER_120_2435 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X32 FILLER_121_993 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X32 FILLER_121_1057 ();
 FILLCELL_X32 FILLER_121_1089 ();
 FILLCELL_X32 FILLER_121_1121 ();
 FILLCELL_X32 FILLER_121_1153 ();
 FILLCELL_X32 FILLER_121_1185 ();
 FILLCELL_X32 FILLER_121_1217 ();
 FILLCELL_X8 FILLER_121_1249 ();
 FILLCELL_X4 FILLER_121_1257 ();
 FILLCELL_X2 FILLER_121_1261 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X32 FILLER_121_1744 ();
 FILLCELL_X32 FILLER_121_1776 ();
 FILLCELL_X32 FILLER_121_1808 ();
 FILLCELL_X32 FILLER_121_1840 ();
 FILLCELL_X32 FILLER_121_1872 ();
 FILLCELL_X32 FILLER_121_1904 ();
 FILLCELL_X32 FILLER_121_1936 ();
 FILLCELL_X32 FILLER_121_1968 ();
 FILLCELL_X32 FILLER_121_2000 ();
 FILLCELL_X32 FILLER_121_2032 ();
 FILLCELL_X32 FILLER_121_2064 ();
 FILLCELL_X32 FILLER_121_2096 ();
 FILLCELL_X32 FILLER_121_2128 ();
 FILLCELL_X32 FILLER_121_2160 ();
 FILLCELL_X32 FILLER_121_2192 ();
 FILLCELL_X32 FILLER_121_2224 ();
 FILLCELL_X32 FILLER_121_2256 ();
 FILLCELL_X32 FILLER_121_2288 ();
 FILLCELL_X32 FILLER_121_2320 ();
 FILLCELL_X32 FILLER_121_2352 ();
 FILLCELL_X32 FILLER_121_2384 ();
 FILLCELL_X16 FILLER_121_2416 ();
 FILLCELL_X4 FILLER_121_2432 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X32 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_122_1240 ();
 FILLCELL_X32 FILLER_122_1272 ();
 FILLCELL_X32 FILLER_122_1304 ();
 FILLCELL_X32 FILLER_122_1336 ();
 FILLCELL_X32 FILLER_122_1368 ();
 FILLCELL_X32 FILLER_122_1400 ();
 FILLCELL_X32 FILLER_122_1432 ();
 FILLCELL_X32 FILLER_122_1464 ();
 FILLCELL_X32 FILLER_122_1496 ();
 FILLCELL_X32 FILLER_122_1528 ();
 FILLCELL_X32 FILLER_122_1560 ();
 FILLCELL_X32 FILLER_122_1592 ();
 FILLCELL_X32 FILLER_122_1624 ();
 FILLCELL_X32 FILLER_122_1656 ();
 FILLCELL_X32 FILLER_122_1688 ();
 FILLCELL_X32 FILLER_122_1720 ();
 FILLCELL_X32 FILLER_122_1752 ();
 FILLCELL_X32 FILLER_122_1784 ();
 FILLCELL_X32 FILLER_122_1816 ();
 FILLCELL_X32 FILLER_122_1848 ();
 FILLCELL_X8 FILLER_122_1880 ();
 FILLCELL_X4 FILLER_122_1888 ();
 FILLCELL_X2 FILLER_122_1892 ();
 FILLCELL_X32 FILLER_122_1895 ();
 FILLCELL_X32 FILLER_122_1927 ();
 FILLCELL_X32 FILLER_122_1959 ();
 FILLCELL_X32 FILLER_122_1991 ();
 FILLCELL_X32 FILLER_122_2023 ();
 FILLCELL_X32 FILLER_122_2055 ();
 FILLCELL_X32 FILLER_122_2087 ();
 FILLCELL_X32 FILLER_122_2119 ();
 FILLCELL_X32 FILLER_122_2151 ();
 FILLCELL_X32 FILLER_122_2183 ();
 FILLCELL_X32 FILLER_122_2215 ();
 FILLCELL_X32 FILLER_122_2247 ();
 FILLCELL_X32 FILLER_122_2279 ();
 FILLCELL_X32 FILLER_122_2311 ();
 FILLCELL_X32 FILLER_122_2343 ();
 FILLCELL_X32 FILLER_122_2375 ();
 FILLCELL_X16 FILLER_122_2407 ();
 FILLCELL_X8 FILLER_122_2423 ();
 FILLCELL_X4 FILLER_122_2431 ();
 FILLCELL_X1 FILLER_122_2435 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X32 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1121 ();
 FILLCELL_X32 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X32 FILLER_123_1217 ();
 FILLCELL_X8 FILLER_123_1249 ();
 FILLCELL_X4 FILLER_123_1257 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X32 FILLER_123_1744 ();
 FILLCELL_X32 FILLER_123_1776 ();
 FILLCELL_X32 FILLER_123_1808 ();
 FILLCELL_X32 FILLER_123_1840 ();
 FILLCELL_X32 FILLER_123_1872 ();
 FILLCELL_X32 FILLER_123_1904 ();
 FILLCELL_X32 FILLER_123_1936 ();
 FILLCELL_X32 FILLER_123_1968 ();
 FILLCELL_X32 FILLER_123_2000 ();
 FILLCELL_X32 FILLER_123_2032 ();
 FILLCELL_X32 FILLER_123_2064 ();
 FILLCELL_X32 FILLER_123_2096 ();
 FILLCELL_X32 FILLER_123_2128 ();
 FILLCELL_X32 FILLER_123_2160 ();
 FILLCELL_X32 FILLER_123_2192 ();
 FILLCELL_X32 FILLER_123_2224 ();
 FILLCELL_X32 FILLER_123_2256 ();
 FILLCELL_X32 FILLER_123_2288 ();
 FILLCELL_X32 FILLER_123_2320 ();
 FILLCELL_X32 FILLER_123_2352 ();
 FILLCELL_X32 FILLER_123_2384 ();
 FILLCELL_X16 FILLER_123_2416 ();
 FILLCELL_X4 FILLER_123_2432 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X32 FILLER_124_1592 ();
 FILLCELL_X32 FILLER_124_1624 ();
 FILLCELL_X32 FILLER_124_1656 ();
 FILLCELL_X32 FILLER_124_1688 ();
 FILLCELL_X32 FILLER_124_1720 ();
 FILLCELL_X32 FILLER_124_1752 ();
 FILLCELL_X32 FILLER_124_1784 ();
 FILLCELL_X32 FILLER_124_1816 ();
 FILLCELL_X32 FILLER_124_1848 ();
 FILLCELL_X8 FILLER_124_1880 ();
 FILLCELL_X4 FILLER_124_1888 ();
 FILLCELL_X2 FILLER_124_1892 ();
 FILLCELL_X32 FILLER_124_1895 ();
 FILLCELL_X32 FILLER_124_1927 ();
 FILLCELL_X32 FILLER_124_1959 ();
 FILLCELL_X32 FILLER_124_1991 ();
 FILLCELL_X32 FILLER_124_2023 ();
 FILLCELL_X32 FILLER_124_2055 ();
 FILLCELL_X32 FILLER_124_2087 ();
 FILLCELL_X32 FILLER_124_2119 ();
 FILLCELL_X32 FILLER_124_2151 ();
 FILLCELL_X32 FILLER_124_2183 ();
 FILLCELL_X32 FILLER_124_2215 ();
 FILLCELL_X32 FILLER_124_2247 ();
 FILLCELL_X32 FILLER_124_2279 ();
 FILLCELL_X32 FILLER_124_2311 ();
 FILLCELL_X32 FILLER_124_2343 ();
 FILLCELL_X32 FILLER_124_2375 ();
 FILLCELL_X16 FILLER_124_2407 ();
 FILLCELL_X8 FILLER_124_2423 ();
 FILLCELL_X4 FILLER_124_2431 ();
 FILLCELL_X1 FILLER_124_2435 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X32 FILLER_125_1089 ();
 FILLCELL_X32 FILLER_125_1121 ();
 FILLCELL_X32 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1185 ();
 FILLCELL_X32 FILLER_125_1217 ();
 FILLCELL_X8 FILLER_125_1249 ();
 FILLCELL_X4 FILLER_125_1257 ();
 FILLCELL_X2 FILLER_125_1261 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X32 FILLER_125_1712 ();
 FILLCELL_X32 FILLER_125_1744 ();
 FILLCELL_X32 FILLER_125_1776 ();
 FILLCELL_X32 FILLER_125_1808 ();
 FILLCELL_X32 FILLER_125_1840 ();
 FILLCELL_X32 FILLER_125_1872 ();
 FILLCELL_X32 FILLER_125_1904 ();
 FILLCELL_X32 FILLER_125_1936 ();
 FILLCELL_X32 FILLER_125_1968 ();
 FILLCELL_X32 FILLER_125_2000 ();
 FILLCELL_X32 FILLER_125_2032 ();
 FILLCELL_X32 FILLER_125_2064 ();
 FILLCELL_X32 FILLER_125_2096 ();
 FILLCELL_X32 FILLER_125_2128 ();
 FILLCELL_X32 FILLER_125_2160 ();
 FILLCELL_X32 FILLER_125_2192 ();
 FILLCELL_X32 FILLER_125_2224 ();
 FILLCELL_X32 FILLER_125_2256 ();
 FILLCELL_X32 FILLER_125_2288 ();
 FILLCELL_X32 FILLER_125_2320 ();
 FILLCELL_X32 FILLER_125_2352 ();
 FILLCELL_X32 FILLER_125_2384 ();
 FILLCELL_X16 FILLER_125_2416 ();
 FILLCELL_X4 FILLER_125_2432 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X32 FILLER_126_1112 ();
 FILLCELL_X32 FILLER_126_1144 ();
 FILLCELL_X32 FILLER_126_1176 ();
 FILLCELL_X32 FILLER_126_1208 ();
 FILLCELL_X32 FILLER_126_1240 ();
 FILLCELL_X32 FILLER_126_1272 ();
 FILLCELL_X32 FILLER_126_1304 ();
 FILLCELL_X32 FILLER_126_1336 ();
 FILLCELL_X32 FILLER_126_1368 ();
 FILLCELL_X32 FILLER_126_1400 ();
 FILLCELL_X32 FILLER_126_1432 ();
 FILLCELL_X32 FILLER_126_1464 ();
 FILLCELL_X32 FILLER_126_1496 ();
 FILLCELL_X32 FILLER_126_1528 ();
 FILLCELL_X32 FILLER_126_1560 ();
 FILLCELL_X32 FILLER_126_1592 ();
 FILLCELL_X32 FILLER_126_1624 ();
 FILLCELL_X32 FILLER_126_1656 ();
 FILLCELL_X32 FILLER_126_1688 ();
 FILLCELL_X32 FILLER_126_1720 ();
 FILLCELL_X32 FILLER_126_1752 ();
 FILLCELL_X32 FILLER_126_1784 ();
 FILLCELL_X32 FILLER_126_1816 ();
 FILLCELL_X32 FILLER_126_1848 ();
 FILLCELL_X8 FILLER_126_1880 ();
 FILLCELL_X4 FILLER_126_1888 ();
 FILLCELL_X2 FILLER_126_1892 ();
 FILLCELL_X32 FILLER_126_1895 ();
 FILLCELL_X32 FILLER_126_1927 ();
 FILLCELL_X32 FILLER_126_1959 ();
 FILLCELL_X32 FILLER_126_1991 ();
 FILLCELL_X32 FILLER_126_2023 ();
 FILLCELL_X32 FILLER_126_2055 ();
 FILLCELL_X32 FILLER_126_2087 ();
 FILLCELL_X32 FILLER_126_2119 ();
 FILLCELL_X32 FILLER_126_2151 ();
 FILLCELL_X32 FILLER_126_2183 ();
 FILLCELL_X32 FILLER_126_2215 ();
 FILLCELL_X32 FILLER_126_2247 ();
 FILLCELL_X32 FILLER_126_2279 ();
 FILLCELL_X32 FILLER_126_2311 ();
 FILLCELL_X32 FILLER_126_2343 ();
 FILLCELL_X32 FILLER_126_2375 ();
 FILLCELL_X16 FILLER_126_2407 ();
 FILLCELL_X8 FILLER_126_2423 ();
 FILLCELL_X4 FILLER_126_2431 ();
 FILLCELL_X1 FILLER_126_2435 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X32 FILLER_127_1712 ();
 FILLCELL_X32 FILLER_127_1744 ();
 FILLCELL_X32 FILLER_127_1776 ();
 FILLCELL_X32 FILLER_127_1808 ();
 FILLCELL_X32 FILLER_127_1840 ();
 FILLCELL_X32 FILLER_127_1872 ();
 FILLCELL_X32 FILLER_127_1904 ();
 FILLCELL_X32 FILLER_127_1936 ();
 FILLCELL_X32 FILLER_127_1968 ();
 FILLCELL_X32 FILLER_127_2000 ();
 FILLCELL_X32 FILLER_127_2032 ();
 FILLCELL_X32 FILLER_127_2064 ();
 FILLCELL_X32 FILLER_127_2096 ();
 FILLCELL_X32 FILLER_127_2128 ();
 FILLCELL_X32 FILLER_127_2160 ();
 FILLCELL_X32 FILLER_127_2192 ();
 FILLCELL_X32 FILLER_127_2224 ();
 FILLCELL_X32 FILLER_127_2256 ();
 FILLCELL_X32 FILLER_127_2288 ();
 FILLCELL_X32 FILLER_127_2320 ();
 FILLCELL_X32 FILLER_127_2352 ();
 FILLCELL_X32 FILLER_127_2384 ();
 FILLCELL_X16 FILLER_127_2416 ();
 FILLCELL_X4 FILLER_127_2432 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X32 FILLER_128_1112 ();
 FILLCELL_X32 FILLER_128_1144 ();
 FILLCELL_X32 FILLER_128_1176 ();
 FILLCELL_X32 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_128_1240 ();
 FILLCELL_X32 FILLER_128_1272 ();
 FILLCELL_X32 FILLER_128_1304 ();
 FILLCELL_X32 FILLER_128_1336 ();
 FILLCELL_X32 FILLER_128_1368 ();
 FILLCELL_X32 FILLER_128_1400 ();
 FILLCELL_X32 FILLER_128_1432 ();
 FILLCELL_X32 FILLER_128_1464 ();
 FILLCELL_X32 FILLER_128_1496 ();
 FILLCELL_X32 FILLER_128_1528 ();
 FILLCELL_X32 FILLER_128_1560 ();
 FILLCELL_X32 FILLER_128_1592 ();
 FILLCELL_X32 FILLER_128_1624 ();
 FILLCELL_X32 FILLER_128_1656 ();
 FILLCELL_X32 FILLER_128_1688 ();
 FILLCELL_X32 FILLER_128_1720 ();
 FILLCELL_X32 FILLER_128_1752 ();
 FILLCELL_X32 FILLER_128_1784 ();
 FILLCELL_X32 FILLER_128_1816 ();
 FILLCELL_X32 FILLER_128_1848 ();
 FILLCELL_X8 FILLER_128_1880 ();
 FILLCELL_X4 FILLER_128_1888 ();
 FILLCELL_X2 FILLER_128_1892 ();
 FILLCELL_X32 FILLER_128_1895 ();
 FILLCELL_X32 FILLER_128_1927 ();
 FILLCELL_X32 FILLER_128_1959 ();
 FILLCELL_X32 FILLER_128_1991 ();
 FILLCELL_X32 FILLER_128_2023 ();
 FILLCELL_X32 FILLER_128_2055 ();
 FILLCELL_X32 FILLER_128_2087 ();
 FILLCELL_X32 FILLER_128_2119 ();
 FILLCELL_X32 FILLER_128_2151 ();
 FILLCELL_X32 FILLER_128_2183 ();
 FILLCELL_X32 FILLER_128_2215 ();
 FILLCELL_X32 FILLER_128_2247 ();
 FILLCELL_X32 FILLER_128_2279 ();
 FILLCELL_X32 FILLER_128_2311 ();
 FILLCELL_X32 FILLER_128_2343 ();
 FILLCELL_X32 FILLER_128_2375 ();
 FILLCELL_X16 FILLER_128_2407 ();
 FILLCELL_X8 FILLER_128_2423 ();
 FILLCELL_X4 FILLER_128_2431 ();
 FILLCELL_X1 FILLER_128_2435 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X32 FILLER_129_1089 ();
 FILLCELL_X32 FILLER_129_1121 ();
 FILLCELL_X32 FILLER_129_1153 ();
 FILLCELL_X32 FILLER_129_1185 ();
 FILLCELL_X32 FILLER_129_1217 ();
 FILLCELL_X8 FILLER_129_1249 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X32 FILLER_129_1680 ();
 FILLCELL_X32 FILLER_129_1712 ();
 FILLCELL_X32 FILLER_129_1744 ();
 FILLCELL_X32 FILLER_129_1776 ();
 FILLCELL_X32 FILLER_129_1808 ();
 FILLCELL_X32 FILLER_129_1840 ();
 FILLCELL_X32 FILLER_129_1872 ();
 FILLCELL_X32 FILLER_129_1904 ();
 FILLCELL_X32 FILLER_129_1936 ();
 FILLCELL_X32 FILLER_129_1968 ();
 FILLCELL_X32 FILLER_129_2000 ();
 FILLCELL_X32 FILLER_129_2032 ();
 FILLCELL_X32 FILLER_129_2064 ();
 FILLCELL_X32 FILLER_129_2096 ();
 FILLCELL_X32 FILLER_129_2128 ();
 FILLCELL_X32 FILLER_129_2160 ();
 FILLCELL_X32 FILLER_129_2192 ();
 FILLCELL_X32 FILLER_129_2224 ();
 FILLCELL_X32 FILLER_129_2256 ();
 FILLCELL_X32 FILLER_129_2288 ();
 FILLCELL_X32 FILLER_129_2320 ();
 FILLCELL_X32 FILLER_129_2352 ();
 FILLCELL_X32 FILLER_129_2384 ();
 FILLCELL_X16 FILLER_129_2416 ();
 FILLCELL_X4 FILLER_129_2432 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X32 FILLER_130_1080 ();
 FILLCELL_X32 FILLER_130_1112 ();
 FILLCELL_X32 FILLER_130_1144 ();
 FILLCELL_X32 FILLER_130_1176 ();
 FILLCELL_X32 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_130_1240 ();
 FILLCELL_X32 FILLER_130_1272 ();
 FILLCELL_X32 FILLER_130_1304 ();
 FILLCELL_X32 FILLER_130_1336 ();
 FILLCELL_X32 FILLER_130_1368 ();
 FILLCELL_X32 FILLER_130_1400 ();
 FILLCELL_X32 FILLER_130_1432 ();
 FILLCELL_X32 FILLER_130_1464 ();
 FILLCELL_X32 FILLER_130_1496 ();
 FILLCELL_X32 FILLER_130_1528 ();
 FILLCELL_X32 FILLER_130_1560 ();
 FILLCELL_X32 FILLER_130_1592 ();
 FILLCELL_X32 FILLER_130_1624 ();
 FILLCELL_X32 FILLER_130_1656 ();
 FILLCELL_X32 FILLER_130_1688 ();
 FILLCELL_X32 FILLER_130_1720 ();
 FILLCELL_X32 FILLER_130_1752 ();
 FILLCELL_X32 FILLER_130_1784 ();
 FILLCELL_X32 FILLER_130_1816 ();
 FILLCELL_X32 FILLER_130_1848 ();
 FILLCELL_X8 FILLER_130_1880 ();
 FILLCELL_X4 FILLER_130_1888 ();
 FILLCELL_X2 FILLER_130_1892 ();
 FILLCELL_X32 FILLER_130_1895 ();
 FILLCELL_X32 FILLER_130_1927 ();
 FILLCELL_X32 FILLER_130_1959 ();
 FILLCELL_X32 FILLER_130_1991 ();
 FILLCELL_X32 FILLER_130_2023 ();
 FILLCELL_X32 FILLER_130_2055 ();
 FILLCELL_X32 FILLER_130_2087 ();
 FILLCELL_X32 FILLER_130_2119 ();
 FILLCELL_X32 FILLER_130_2151 ();
 FILLCELL_X32 FILLER_130_2183 ();
 FILLCELL_X32 FILLER_130_2215 ();
 FILLCELL_X32 FILLER_130_2247 ();
 FILLCELL_X32 FILLER_130_2279 ();
 FILLCELL_X32 FILLER_130_2311 ();
 FILLCELL_X32 FILLER_130_2343 ();
 FILLCELL_X32 FILLER_130_2375 ();
 FILLCELL_X16 FILLER_130_2407 ();
 FILLCELL_X8 FILLER_130_2423 ();
 FILLCELL_X4 FILLER_130_2431 ();
 FILLCELL_X1 FILLER_130_2435 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X32 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_1025 ();
 FILLCELL_X32 FILLER_131_1057 ();
 FILLCELL_X32 FILLER_131_1089 ();
 FILLCELL_X32 FILLER_131_1121 ();
 FILLCELL_X32 FILLER_131_1153 ();
 FILLCELL_X32 FILLER_131_1185 ();
 FILLCELL_X32 FILLER_131_1217 ();
 FILLCELL_X8 FILLER_131_1249 ();
 FILLCELL_X4 FILLER_131_1257 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X32 FILLER_131_1744 ();
 FILLCELL_X32 FILLER_131_1776 ();
 FILLCELL_X32 FILLER_131_1808 ();
 FILLCELL_X32 FILLER_131_1840 ();
 FILLCELL_X32 FILLER_131_1872 ();
 FILLCELL_X32 FILLER_131_1904 ();
 FILLCELL_X32 FILLER_131_1936 ();
 FILLCELL_X32 FILLER_131_1968 ();
 FILLCELL_X32 FILLER_131_2000 ();
 FILLCELL_X32 FILLER_131_2032 ();
 FILLCELL_X32 FILLER_131_2064 ();
 FILLCELL_X32 FILLER_131_2096 ();
 FILLCELL_X32 FILLER_131_2128 ();
 FILLCELL_X32 FILLER_131_2160 ();
 FILLCELL_X32 FILLER_131_2192 ();
 FILLCELL_X32 FILLER_131_2224 ();
 FILLCELL_X32 FILLER_131_2256 ();
 FILLCELL_X32 FILLER_131_2288 ();
 FILLCELL_X32 FILLER_131_2320 ();
 FILLCELL_X32 FILLER_131_2352 ();
 FILLCELL_X32 FILLER_131_2384 ();
 FILLCELL_X16 FILLER_131_2416 ();
 FILLCELL_X4 FILLER_131_2432 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X32 FILLER_132_1080 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X32 FILLER_132_1144 ();
 FILLCELL_X32 FILLER_132_1176 ();
 FILLCELL_X32 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_132_1240 ();
 FILLCELL_X32 FILLER_132_1272 ();
 FILLCELL_X32 FILLER_132_1304 ();
 FILLCELL_X32 FILLER_132_1336 ();
 FILLCELL_X32 FILLER_132_1368 ();
 FILLCELL_X32 FILLER_132_1400 ();
 FILLCELL_X32 FILLER_132_1432 ();
 FILLCELL_X32 FILLER_132_1464 ();
 FILLCELL_X32 FILLER_132_1496 ();
 FILLCELL_X32 FILLER_132_1528 ();
 FILLCELL_X32 FILLER_132_1560 ();
 FILLCELL_X32 FILLER_132_1592 ();
 FILLCELL_X32 FILLER_132_1624 ();
 FILLCELL_X32 FILLER_132_1656 ();
 FILLCELL_X32 FILLER_132_1688 ();
 FILLCELL_X32 FILLER_132_1720 ();
 FILLCELL_X32 FILLER_132_1752 ();
 FILLCELL_X32 FILLER_132_1784 ();
 FILLCELL_X32 FILLER_132_1816 ();
 FILLCELL_X32 FILLER_132_1848 ();
 FILLCELL_X8 FILLER_132_1880 ();
 FILLCELL_X4 FILLER_132_1888 ();
 FILLCELL_X2 FILLER_132_1892 ();
 FILLCELL_X32 FILLER_132_1895 ();
 FILLCELL_X32 FILLER_132_1927 ();
 FILLCELL_X32 FILLER_132_1959 ();
 FILLCELL_X32 FILLER_132_1991 ();
 FILLCELL_X32 FILLER_132_2023 ();
 FILLCELL_X32 FILLER_132_2055 ();
 FILLCELL_X32 FILLER_132_2087 ();
 FILLCELL_X32 FILLER_132_2119 ();
 FILLCELL_X32 FILLER_132_2151 ();
 FILLCELL_X32 FILLER_132_2183 ();
 FILLCELL_X32 FILLER_132_2215 ();
 FILLCELL_X32 FILLER_132_2247 ();
 FILLCELL_X32 FILLER_132_2279 ();
 FILLCELL_X32 FILLER_132_2311 ();
 FILLCELL_X32 FILLER_132_2343 ();
 FILLCELL_X32 FILLER_132_2375 ();
 FILLCELL_X16 FILLER_132_2407 ();
 FILLCELL_X8 FILLER_132_2423 ();
 FILLCELL_X4 FILLER_132_2431 ();
 FILLCELL_X1 FILLER_132_2435 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X32 FILLER_133_1121 ();
 FILLCELL_X32 FILLER_133_1153 ();
 FILLCELL_X32 FILLER_133_1185 ();
 FILLCELL_X32 FILLER_133_1217 ();
 FILLCELL_X8 FILLER_133_1249 ();
 FILLCELL_X4 FILLER_133_1257 ();
 FILLCELL_X2 FILLER_133_1261 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X32 FILLER_133_1584 ();
 FILLCELL_X32 FILLER_133_1616 ();
 FILLCELL_X32 FILLER_133_1648 ();
 FILLCELL_X32 FILLER_133_1680 ();
 FILLCELL_X32 FILLER_133_1712 ();
 FILLCELL_X32 FILLER_133_1744 ();
 FILLCELL_X32 FILLER_133_1776 ();
 FILLCELL_X32 FILLER_133_1808 ();
 FILLCELL_X32 FILLER_133_1840 ();
 FILLCELL_X32 FILLER_133_1872 ();
 FILLCELL_X32 FILLER_133_1904 ();
 FILLCELL_X32 FILLER_133_1936 ();
 FILLCELL_X32 FILLER_133_1968 ();
 FILLCELL_X32 FILLER_133_2000 ();
 FILLCELL_X32 FILLER_133_2032 ();
 FILLCELL_X32 FILLER_133_2064 ();
 FILLCELL_X32 FILLER_133_2096 ();
 FILLCELL_X32 FILLER_133_2128 ();
 FILLCELL_X32 FILLER_133_2160 ();
 FILLCELL_X32 FILLER_133_2192 ();
 FILLCELL_X32 FILLER_133_2224 ();
 FILLCELL_X32 FILLER_133_2256 ();
 FILLCELL_X32 FILLER_133_2288 ();
 FILLCELL_X32 FILLER_133_2320 ();
 FILLCELL_X32 FILLER_133_2352 ();
 FILLCELL_X32 FILLER_133_2384 ();
 FILLCELL_X16 FILLER_133_2416 ();
 FILLCELL_X4 FILLER_133_2432 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_134_1048 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X32 FILLER_134_1592 ();
 FILLCELL_X32 FILLER_134_1624 ();
 FILLCELL_X32 FILLER_134_1656 ();
 FILLCELL_X32 FILLER_134_1688 ();
 FILLCELL_X32 FILLER_134_1720 ();
 FILLCELL_X32 FILLER_134_1752 ();
 FILLCELL_X32 FILLER_134_1784 ();
 FILLCELL_X32 FILLER_134_1816 ();
 FILLCELL_X32 FILLER_134_1848 ();
 FILLCELL_X8 FILLER_134_1880 ();
 FILLCELL_X4 FILLER_134_1888 ();
 FILLCELL_X2 FILLER_134_1892 ();
 FILLCELL_X32 FILLER_134_1895 ();
 FILLCELL_X32 FILLER_134_1927 ();
 FILLCELL_X32 FILLER_134_1959 ();
 FILLCELL_X32 FILLER_134_1991 ();
 FILLCELL_X32 FILLER_134_2023 ();
 FILLCELL_X32 FILLER_134_2055 ();
 FILLCELL_X32 FILLER_134_2087 ();
 FILLCELL_X32 FILLER_134_2119 ();
 FILLCELL_X32 FILLER_134_2151 ();
 FILLCELL_X32 FILLER_134_2183 ();
 FILLCELL_X32 FILLER_134_2215 ();
 FILLCELL_X32 FILLER_134_2247 ();
 FILLCELL_X32 FILLER_134_2279 ();
 FILLCELL_X32 FILLER_134_2311 ();
 FILLCELL_X32 FILLER_134_2343 ();
 FILLCELL_X32 FILLER_134_2375 ();
 FILLCELL_X16 FILLER_134_2407 ();
 FILLCELL_X8 FILLER_134_2423 ();
 FILLCELL_X4 FILLER_134_2431 ();
 FILLCELL_X1 FILLER_134_2435 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X32 FILLER_135_993 ();
 FILLCELL_X32 FILLER_135_1025 ();
 FILLCELL_X32 FILLER_135_1057 ();
 FILLCELL_X32 FILLER_135_1089 ();
 FILLCELL_X32 FILLER_135_1121 ();
 FILLCELL_X32 FILLER_135_1153 ();
 FILLCELL_X32 FILLER_135_1185 ();
 FILLCELL_X32 FILLER_135_1217 ();
 FILLCELL_X8 FILLER_135_1249 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X32 FILLER_135_1584 ();
 FILLCELL_X32 FILLER_135_1616 ();
 FILLCELL_X32 FILLER_135_1648 ();
 FILLCELL_X32 FILLER_135_1680 ();
 FILLCELL_X32 FILLER_135_1712 ();
 FILLCELL_X32 FILLER_135_1744 ();
 FILLCELL_X32 FILLER_135_1776 ();
 FILLCELL_X32 FILLER_135_1808 ();
 FILLCELL_X32 FILLER_135_1840 ();
 FILLCELL_X32 FILLER_135_1872 ();
 FILLCELL_X32 FILLER_135_1904 ();
 FILLCELL_X32 FILLER_135_1936 ();
 FILLCELL_X32 FILLER_135_1968 ();
 FILLCELL_X32 FILLER_135_2000 ();
 FILLCELL_X32 FILLER_135_2032 ();
 FILLCELL_X32 FILLER_135_2064 ();
 FILLCELL_X32 FILLER_135_2096 ();
 FILLCELL_X32 FILLER_135_2128 ();
 FILLCELL_X32 FILLER_135_2160 ();
 FILLCELL_X32 FILLER_135_2192 ();
 FILLCELL_X32 FILLER_135_2224 ();
 FILLCELL_X32 FILLER_135_2256 ();
 FILLCELL_X32 FILLER_135_2288 ();
 FILLCELL_X32 FILLER_135_2320 ();
 FILLCELL_X32 FILLER_135_2352 ();
 FILLCELL_X32 FILLER_135_2384 ();
 FILLCELL_X16 FILLER_135_2416 ();
 FILLCELL_X4 FILLER_135_2432 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X32 FILLER_136_1016 ();
 FILLCELL_X32 FILLER_136_1048 ();
 FILLCELL_X32 FILLER_136_1080 ();
 FILLCELL_X32 FILLER_136_1112 ();
 FILLCELL_X32 FILLER_136_1144 ();
 FILLCELL_X32 FILLER_136_1176 ();
 FILLCELL_X32 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_136_1240 ();
 FILLCELL_X32 FILLER_136_1272 ();
 FILLCELL_X32 FILLER_136_1304 ();
 FILLCELL_X32 FILLER_136_1336 ();
 FILLCELL_X32 FILLER_136_1368 ();
 FILLCELL_X32 FILLER_136_1400 ();
 FILLCELL_X32 FILLER_136_1432 ();
 FILLCELL_X32 FILLER_136_1464 ();
 FILLCELL_X32 FILLER_136_1496 ();
 FILLCELL_X32 FILLER_136_1528 ();
 FILLCELL_X32 FILLER_136_1560 ();
 FILLCELL_X32 FILLER_136_1592 ();
 FILLCELL_X32 FILLER_136_1624 ();
 FILLCELL_X32 FILLER_136_1656 ();
 FILLCELL_X32 FILLER_136_1688 ();
 FILLCELL_X32 FILLER_136_1720 ();
 FILLCELL_X32 FILLER_136_1752 ();
 FILLCELL_X32 FILLER_136_1784 ();
 FILLCELL_X32 FILLER_136_1816 ();
 FILLCELL_X32 FILLER_136_1848 ();
 FILLCELL_X8 FILLER_136_1880 ();
 FILLCELL_X4 FILLER_136_1888 ();
 FILLCELL_X2 FILLER_136_1892 ();
 FILLCELL_X32 FILLER_136_1895 ();
 FILLCELL_X32 FILLER_136_1927 ();
 FILLCELL_X32 FILLER_136_1959 ();
 FILLCELL_X32 FILLER_136_1991 ();
 FILLCELL_X32 FILLER_136_2023 ();
 FILLCELL_X32 FILLER_136_2055 ();
 FILLCELL_X32 FILLER_136_2087 ();
 FILLCELL_X32 FILLER_136_2119 ();
 FILLCELL_X32 FILLER_136_2151 ();
 FILLCELL_X32 FILLER_136_2183 ();
 FILLCELL_X32 FILLER_136_2215 ();
 FILLCELL_X32 FILLER_136_2247 ();
 FILLCELL_X32 FILLER_136_2279 ();
 FILLCELL_X32 FILLER_136_2311 ();
 FILLCELL_X32 FILLER_136_2343 ();
 FILLCELL_X32 FILLER_136_2375 ();
 FILLCELL_X16 FILLER_136_2407 ();
 FILLCELL_X8 FILLER_136_2423 ();
 FILLCELL_X4 FILLER_136_2431 ();
 FILLCELL_X1 FILLER_136_2435 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X32 FILLER_137_961 ();
 FILLCELL_X32 FILLER_137_993 ();
 FILLCELL_X32 FILLER_137_1025 ();
 FILLCELL_X32 FILLER_137_1057 ();
 FILLCELL_X32 FILLER_137_1089 ();
 FILLCELL_X32 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1153 ();
 FILLCELL_X32 FILLER_137_1185 ();
 FILLCELL_X32 FILLER_137_1217 ();
 FILLCELL_X8 FILLER_137_1249 ();
 FILLCELL_X4 FILLER_137_1257 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X32 FILLER_137_1584 ();
 FILLCELL_X32 FILLER_137_1616 ();
 FILLCELL_X32 FILLER_137_1648 ();
 FILLCELL_X32 FILLER_137_1680 ();
 FILLCELL_X32 FILLER_137_1712 ();
 FILLCELL_X32 FILLER_137_1744 ();
 FILLCELL_X32 FILLER_137_1776 ();
 FILLCELL_X32 FILLER_137_1808 ();
 FILLCELL_X32 FILLER_137_1840 ();
 FILLCELL_X32 FILLER_137_1872 ();
 FILLCELL_X32 FILLER_137_1904 ();
 FILLCELL_X32 FILLER_137_1936 ();
 FILLCELL_X32 FILLER_137_1968 ();
 FILLCELL_X32 FILLER_137_2000 ();
 FILLCELL_X32 FILLER_137_2032 ();
 FILLCELL_X32 FILLER_137_2064 ();
 FILLCELL_X32 FILLER_137_2096 ();
 FILLCELL_X32 FILLER_137_2128 ();
 FILLCELL_X32 FILLER_137_2160 ();
 FILLCELL_X32 FILLER_137_2192 ();
 FILLCELL_X32 FILLER_137_2224 ();
 FILLCELL_X32 FILLER_137_2256 ();
 FILLCELL_X32 FILLER_137_2288 ();
 FILLCELL_X32 FILLER_137_2320 ();
 FILLCELL_X32 FILLER_137_2352 ();
 FILLCELL_X32 FILLER_137_2384 ();
 FILLCELL_X16 FILLER_137_2416 ();
 FILLCELL_X4 FILLER_137_2432 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X32 FILLER_138_984 ();
 FILLCELL_X32 FILLER_138_1016 ();
 FILLCELL_X32 FILLER_138_1048 ();
 FILLCELL_X32 FILLER_138_1080 ();
 FILLCELL_X32 FILLER_138_1112 ();
 FILLCELL_X32 FILLER_138_1144 ();
 FILLCELL_X32 FILLER_138_1176 ();
 FILLCELL_X32 FILLER_138_1208 ();
 FILLCELL_X32 FILLER_138_1240 ();
 FILLCELL_X32 FILLER_138_1272 ();
 FILLCELL_X32 FILLER_138_1304 ();
 FILLCELL_X32 FILLER_138_1336 ();
 FILLCELL_X32 FILLER_138_1368 ();
 FILLCELL_X32 FILLER_138_1400 ();
 FILLCELL_X32 FILLER_138_1432 ();
 FILLCELL_X32 FILLER_138_1464 ();
 FILLCELL_X32 FILLER_138_1496 ();
 FILLCELL_X32 FILLER_138_1528 ();
 FILLCELL_X32 FILLER_138_1560 ();
 FILLCELL_X32 FILLER_138_1592 ();
 FILLCELL_X32 FILLER_138_1624 ();
 FILLCELL_X32 FILLER_138_1656 ();
 FILLCELL_X32 FILLER_138_1688 ();
 FILLCELL_X32 FILLER_138_1720 ();
 FILLCELL_X32 FILLER_138_1752 ();
 FILLCELL_X32 FILLER_138_1784 ();
 FILLCELL_X32 FILLER_138_1816 ();
 FILLCELL_X32 FILLER_138_1848 ();
 FILLCELL_X8 FILLER_138_1880 ();
 FILLCELL_X4 FILLER_138_1888 ();
 FILLCELL_X2 FILLER_138_1892 ();
 FILLCELL_X32 FILLER_138_1895 ();
 FILLCELL_X32 FILLER_138_1927 ();
 FILLCELL_X32 FILLER_138_1959 ();
 FILLCELL_X32 FILLER_138_1991 ();
 FILLCELL_X32 FILLER_138_2023 ();
 FILLCELL_X32 FILLER_138_2055 ();
 FILLCELL_X32 FILLER_138_2087 ();
 FILLCELL_X32 FILLER_138_2119 ();
 FILLCELL_X32 FILLER_138_2151 ();
 FILLCELL_X32 FILLER_138_2183 ();
 FILLCELL_X32 FILLER_138_2215 ();
 FILLCELL_X32 FILLER_138_2247 ();
 FILLCELL_X32 FILLER_138_2279 ();
 FILLCELL_X32 FILLER_138_2311 ();
 FILLCELL_X32 FILLER_138_2343 ();
 FILLCELL_X32 FILLER_138_2375 ();
 FILLCELL_X16 FILLER_138_2407 ();
 FILLCELL_X8 FILLER_138_2423 ();
 FILLCELL_X4 FILLER_138_2431 ();
 FILLCELL_X1 FILLER_138_2435 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X32 FILLER_139_1057 ();
 FILLCELL_X32 FILLER_139_1089 ();
 FILLCELL_X32 FILLER_139_1121 ();
 FILLCELL_X32 FILLER_139_1153 ();
 FILLCELL_X32 FILLER_139_1185 ();
 FILLCELL_X32 FILLER_139_1217 ();
 FILLCELL_X8 FILLER_139_1249 ();
 FILLCELL_X4 FILLER_139_1257 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X32 FILLER_139_1584 ();
 FILLCELL_X32 FILLER_139_1616 ();
 FILLCELL_X32 FILLER_139_1648 ();
 FILLCELL_X32 FILLER_139_1680 ();
 FILLCELL_X32 FILLER_139_1712 ();
 FILLCELL_X32 FILLER_139_1744 ();
 FILLCELL_X32 FILLER_139_1776 ();
 FILLCELL_X32 FILLER_139_1808 ();
 FILLCELL_X32 FILLER_139_1840 ();
 FILLCELL_X32 FILLER_139_1872 ();
 FILLCELL_X32 FILLER_139_1904 ();
 FILLCELL_X32 FILLER_139_1936 ();
 FILLCELL_X32 FILLER_139_1968 ();
 FILLCELL_X32 FILLER_139_2000 ();
 FILLCELL_X32 FILLER_139_2032 ();
 FILLCELL_X32 FILLER_139_2064 ();
 FILLCELL_X32 FILLER_139_2096 ();
 FILLCELL_X32 FILLER_139_2128 ();
 FILLCELL_X32 FILLER_139_2160 ();
 FILLCELL_X32 FILLER_139_2192 ();
 FILLCELL_X32 FILLER_139_2224 ();
 FILLCELL_X32 FILLER_139_2256 ();
 FILLCELL_X32 FILLER_139_2288 ();
 FILLCELL_X32 FILLER_139_2320 ();
 FILLCELL_X32 FILLER_139_2352 ();
 FILLCELL_X32 FILLER_139_2384 ();
 FILLCELL_X16 FILLER_139_2416 ();
 FILLCELL_X4 FILLER_139_2432 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X32 FILLER_140_1592 ();
 FILLCELL_X32 FILLER_140_1624 ();
 FILLCELL_X32 FILLER_140_1656 ();
 FILLCELL_X32 FILLER_140_1688 ();
 FILLCELL_X32 FILLER_140_1720 ();
 FILLCELL_X32 FILLER_140_1752 ();
 FILLCELL_X32 FILLER_140_1784 ();
 FILLCELL_X32 FILLER_140_1816 ();
 FILLCELL_X32 FILLER_140_1848 ();
 FILLCELL_X8 FILLER_140_1880 ();
 FILLCELL_X4 FILLER_140_1888 ();
 FILLCELL_X2 FILLER_140_1892 ();
 FILLCELL_X32 FILLER_140_1895 ();
 FILLCELL_X32 FILLER_140_1927 ();
 FILLCELL_X32 FILLER_140_1959 ();
 FILLCELL_X32 FILLER_140_1991 ();
 FILLCELL_X32 FILLER_140_2023 ();
 FILLCELL_X32 FILLER_140_2055 ();
 FILLCELL_X32 FILLER_140_2087 ();
 FILLCELL_X32 FILLER_140_2119 ();
 FILLCELL_X32 FILLER_140_2151 ();
 FILLCELL_X32 FILLER_140_2183 ();
 FILLCELL_X32 FILLER_140_2215 ();
 FILLCELL_X32 FILLER_140_2247 ();
 FILLCELL_X32 FILLER_140_2279 ();
 FILLCELL_X32 FILLER_140_2311 ();
 FILLCELL_X32 FILLER_140_2343 ();
 FILLCELL_X32 FILLER_140_2375 ();
 FILLCELL_X16 FILLER_140_2407 ();
 FILLCELL_X8 FILLER_140_2423 ();
 FILLCELL_X4 FILLER_140_2431 ();
 FILLCELL_X1 FILLER_140_2435 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X32 FILLER_141_1121 ();
 FILLCELL_X32 FILLER_141_1153 ();
 FILLCELL_X32 FILLER_141_1185 ();
 FILLCELL_X32 FILLER_141_1217 ();
 FILLCELL_X8 FILLER_141_1249 ();
 FILLCELL_X4 FILLER_141_1257 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X32 FILLER_141_1584 ();
 FILLCELL_X32 FILLER_141_1616 ();
 FILLCELL_X32 FILLER_141_1648 ();
 FILLCELL_X32 FILLER_141_1680 ();
 FILLCELL_X32 FILLER_141_1712 ();
 FILLCELL_X32 FILLER_141_1744 ();
 FILLCELL_X32 FILLER_141_1776 ();
 FILLCELL_X32 FILLER_141_1808 ();
 FILLCELL_X32 FILLER_141_1840 ();
 FILLCELL_X32 FILLER_141_1872 ();
 FILLCELL_X32 FILLER_141_1904 ();
 FILLCELL_X32 FILLER_141_1936 ();
 FILLCELL_X32 FILLER_141_1968 ();
 FILLCELL_X32 FILLER_141_2000 ();
 FILLCELL_X32 FILLER_141_2032 ();
 FILLCELL_X32 FILLER_141_2064 ();
 FILLCELL_X32 FILLER_141_2096 ();
 FILLCELL_X32 FILLER_141_2128 ();
 FILLCELL_X32 FILLER_141_2160 ();
 FILLCELL_X32 FILLER_141_2192 ();
 FILLCELL_X32 FILLER_141_2224 ();
 FILLCELL_X32 FILLER_141_2256 ();
 FILLCELL_X32 FILLER_141_2288 ();
 FILLCELL_X32 FILLER_141_2320 ();
 FILLCELL_X32 FILLER_141_2352 ();
 FILLCELL_X32 FILLER_141_2384 ();
 FILLCELL_X16 FILLER_141_2416 ();
 FILLCELL_X4 FILLER_141_2432 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X32 FILLER_142_1624 ();
 FILLCELL_X32 FILLER_142_1656 ();
 FILLCELL_X32 FILLER_142_1688 ();
 FILLCELL_X32 FILLER_142_1720 ();
 FILLCELL_X32 FILLER_142_1752 ();
 FILLCELL_X32 FILLER_142_1784 ();
 FILLCELL_X32 FILLER_142_1816 ();
 FILLCELL_X32 FILLER_142_1848 ();
 FILLCELL_X8 FILLER_142_1880 ();
 FILLCELL_X4 FILLER_142_1888 ();
 FILLCELL_X2 FILLER_142_1892 ();
 FILLCELL_X32 FILLER_142_1895 ();
 FILLCELL_X32 FILLER_142_1927 ();
 FILLCELL_X32 FILLER_142_1959 ();
 FILLCELL_X32 FILLER_142_1991 ();
 FILLCELL_X32 FILLER_142_2023 ();
 FILLCELL_X32 FILLER_142_2055 ();
 FILLCELL_X32 FILLER_142_2087 ();
 FILLCELL_X32 FILLER_142_2119 ();
 FILLCELL_X32 FILLER_142_2151 ();
 FILLCELL_X32 FILLER_142_2183 ();
 FILLCELL_X32 FILLER_142_2215 ();
 FILLCELL_X32 FILLER_142_2247 ();
 FILLCELL_X32 FILLER_142_2279 ();
 FILLCELL_X32 FILLER_142_2311 ();
 FILLCELL_X32 FILLER_142_2343 ();
 FILLCELL_X32 FILLER_142_2375 ();
 FILLCELL_X16 FILLER_142_2407 ();
 FILLCELL_X8 FILLER_142_2423 ();
 FILLCELL_X4 FILLER_142_2431 ();
 FILLCELL_X1 FILLER_142_2435 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X32 FILLER_143_1584 ();
 FILLCELL_X32 FILLER_143_1616 ();
 FILLCELL_X32 FILLER_143_1648 ();
 FILLCELL_X32 FILLER_143_1680 ();
 FILLCELL_X32 FILLER_143_1712 ();
 FILLCELL_X32 FILLER_143_1744 ();
 FILLCELL_X32 FILLER_143_1776 ();
 FILLCELL_X32 FILLER_143_1808 ();
 FILLCELL_X32 FILLER_143_1840 ();
 FILLCELL_X32 FILLER_143_1872 ();
 FILLCELL_X32 FILLER_143_1904 ();
 FILLCELL_X32 FILLER_143_1936 ();
 FILLCELL_X32 FILLER_143_1968 ();
 FILLCELL_X32 FILLER_143_2000 ();
 FILLCELL_X32 FILLER_143_2032 ();
 FILLCELL_X32 FILLER_143_2064 ();
 FILLCELL_X32 FILLER_143_2096 ();
 FILLCELL_X32 FILLER_143_2128 ();
 FILLCELL_X32 FILLER_143_2160 ();
 FILLCELL_X32 FILLER_143_2192 ();
 FILLCELL_X32 FILLER_143_2224 ();
 FILLCELL_X32 FILLER_143_2256 ();
 FILLCELL_X32 FILLER_143_2288 ();
 FILLCELL_X32 FILLER_143_2320 ();
 FILLCELL_X32 FILLER_143_2352 ();
 FILLCELL_X32 FILLER_143_2384 ();
 FILLCELL_X16 FILLER_143_2416 ();
 FILLCELL_X4 FILLER_143_2432 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X32 FILLER_144_1592 ();
 FILLCELL_X32 FILLER_144_1624 ();
 FILLCELL_X32 FILLER_144_1656 ();
 FILLCELL_X32 FILLER_144_1688 ();
 FILLCELL_X32 FILLER_144_1720 ();
 FILLCELL_X32 FILLER_144_1752 ();
 FILLCELL_X32 FILLER_144_1784 ();
 FILLCELL_X32 FILLER_144_1816 ();
 FILLCELL_X32 FILLER_144_1848 ();
 FILLCELL_X8 FILLER_144_1880 ();
 FILLCELL_X4 FILLER_144_1888 ();
 FILLCELL_X2 FILLER_144_1892 ();
 FILLCELL_X32 FILLER_144_1895 ();
 FILLCELL_X32 FILLER_144_1927 ();
 FILLCELL_X32 FILLER_144_1959 ();
 FILLCELL_X32 FILLER_144_1991 ();
 FILLCELL_X32 FILLER_144_2023 ();
 FILLCELL_X32 FILLER_144_2055 ();
 FILLCELL_X32 FILLER_144_2087 ();
 FILLCELL_X32 FILLER_144_2119 ();
 FILLCELL_X32 FILLER_144_2151 ();
 FILLCELL_X32 FILLER_144_2183 ();
 FILLCELL_X32 FILLER_144_2215 ();
 FILLCELL_X32 FILLER_144_2247 ();
 FILLCELL_X32 FILLER_144_2279 ();
 FILLCELL_X32 FILLER_144_2311 ();
 FILLCELL_X32 FILLER_144_2343 ();
 FILLCELL_X32 FILLER_144_2375 ();
 FILLCELL_X16 FILLER_144_2407 ();
 FILLCELL_X8 FILLER_144_2423 ();
 FILLCELL_X4 FILLER_144_2431 ();
 FILLCELL_X1 FILLER_144_2435 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X32 FILLER_145_1776 ();
 FILLCELL_X32 FILLER_145_1808 ();
 FILLCELL_X32 FILLER_145_1840 ();
 FILLCELL_X32 FILLER_145_1872 ();
 FILLCELL_X32 FILLER_145_1904 ();
 FILLCELL_X32 FILLER_145_1936 ();
 FILLCELL_X32 FILLER_145_1968 ();
 FILLCELL_X32 FILLER_145_2000 ();
 FILLCELL_X32 FILLER_145_2032 ();
 FILLCELL_X32 FILLER_145_2064 ();
 FILLCELL_X32 FILLER_145_2096 ();
 FILLCELL_X32 FILLER_145_2128 ();
 FILLCELL_X32 FILLER_145_2160 ();
 FILLCELL_X32 FILLER_145_2192 ();
 FILLCELL_X32 FILLER_145_2224 ();
 FILLCELL_X32 FILLER_145_2256 ();
 FILLCELL_X32 FILLER_145_2288 ();
 FILLCELL_X32 FILLER_145_2320 ();
 FILLCELL_X32 FILLER_145_2352 ();
 FILLCELL_X32 FILLER_145_2384 ();
 FILLCELL_X16 FILLER_145_2416 ();
 FILLCELL_X4 FILLER_145_2432 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X32 FILLER_146_1592 ();
 FILLCELL_X32 FILLER_146_1624 ();
 FILLCELL_X32 FILLER_146_1656 ();
 FILLCELL_X32 FILLER_146_1688 ();
 FILLCELL_X32 FILLER_146_1720 ();
 FILLCELL_X32 FILLER_146_1752 ();
 FILLCELL_X32 FILLER_146_1784 ();
 FILLCELL_X32 FILLER_146_1816 ();
 FILLCELL_X32 FILLER_146_1848 ();
 FILLCELL_X8 FILLER_146_1880 ();
 FILLCELL_X4 FILLER_146_1888 ();
 FILLCELL_X2 FILLER_146_1892 ();
 FILLCELL_X32 FILLER_146_1895 ();
 FILLCELL_X32 FILLER_146_1927 ();
 FILLCELL_X32 FILLER_146_1959 ();
 FILLCELL_X32 FILLER_146_1991 ();
 FILLCELL_X32 FILLER_146_2023 ();
 FILLCELL_X32 FILLER_146_2055 ();
 FILLCELL_X32 FILLER_146_2087 ();
 FILLCELL_X32 FILLER_146_2119 ();
 FILLCELL_X32 FILLER_146_2151 ();
 FILLCELL_X32 FILLER_146_2183 ();
 FILLCELL_X32 FILLER_146_2215 ();
 FILLCELL_X32 FILLER_146_2247 ();
 FILLCELL_X32 FILLER_146_2279 ();
 FILLCELL_X32 FILLER_146_2311 ();
 FILLCELL_X32 FILLER_146_2343 ();
 FILLCELL_X32 FILLER_146_2375 ();
 FILLCELL_X16 FILLER_146_2407 ();
 FILLCELL_X8 FILLER_146_2423 ();
 FILLCELL_X4 FILLER_146_2431 ();
 FILLCELL_X1 FILLER_146_2435 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X32 FILLER_147_1776 ();
 FILLCELL_X32 FILLER_147_1808 ();
 FILLCELL_X32 FILLER_147_1840 ();
 FILLCELL_X32 FILLER_147_1872 ();
 FILLCELL_X32 FILLER_147_1904 ();
 FILLCELL_X32 FILLER_147_1936 ();
 FILLCELL_X32 FILLER_147_1968 ();
 FILLCELL_X32 FILLER_147_2000 ();
 FILLCELL_X32 FILLER_147_2032 ();
 FILLCELL_X32 FILLER_147_2064 ();
 FILLCELL_X32 FILLER_147_2096 ();
 FILLCELL_X32 FILLER_147_2128 ();
 FILLCELL_X32 FILLER_147_2160 ();
 FILLCELL_X32 FILLER_147_2192 ();
 FILLCELL_X32 FILLER_147_2224 ();
 FILLCELL_X32 FILLER_147_2256 ();
 FILLCELL_X32 FILLER_147_2288 ();
 FILLCELL_X32 FILLER_147_2320 ();
 FILLCELL_X32 FILLER_147_2352 ();
 FILLCELL_X32 FILLER_147_2384 ();
 FILLCELL_X16 FILLER_147_2416 ();
 FILLCELL_X4 FILLER_147_2432 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X32 FILLER_148_1592 ();
 FILLCELL_X32 FILLER_148_1624 ();
 FILLCELL_X32 FILLER_148_1656 ();
 FILLCELL_X32 FILLER_148_1688 ();
 FILLCELL_X32 FILLER_148_1720 ();
 FILLCELL_X32 FILLER_148_1752 ();
 FILLCELL_X32 FILLER_148_1784 ();
 FILLCELL_X32 FILLER_148_1816 ();
 FILLCELL_X32 FILLER_148_1848 ();
 FILLCELL_X8 FILLER_148_1880 ();
 FILLCELL_X4 FILLER_148_1888 ();
 FILLCELL_X2 FILLER_148_1892 ();
 FILLCELL_X32 FILLER_148_1895 ();
 FILLCELL_X32 FILLER_148_1927 ();
 FILLCELL_X32 FILLER_148_1959 ();
 FILLCELL_X32 FILLER_148_1991 ();
 FILLCELL_X32 FILLER_148_2023 ();
 FILLCELL_X32 FILLER_148_2055 ();
 FILLCELL_X32 FILLER_148_2087 ();
 FILLCELL_X32 FILLER_148_2119 ();
 FILLCELL_X32 FILLER_148_2151 ();
 FILLCELL_X32 FILLER_148_2183 ();
 FILLCELL_X32 FILLER_148_2215 ();
 FILLCELL_X32 FILLER_148_2247 ();
 FILLCELL_X32 FILLER_148_2279 ();
 FILLCELL_X32 FILLER_148_2311 ();
 FILLCELL_X32 FILLER_148_2343 ();
 FILLCELL_X32 FILLER_148_2375 ();
 FILLCELL_X16 FILLER_148_2407 ();
 FILLCELL_X8 FILLER_148_2423 ();
 FILLCELL_X4 FILLER_148_2431 ();
 FILLCELL_X1 FILLER_148_2435 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X32 FILLER_149_1776 ();
 FILLCELL_X32 FILLER_149_1808 ();
 FILLCELL_X32 FILLER_149_1840 ();
 FILLCELL_X32 FILLER_149_1872 ();
 FILLCELL_X32 FILLER_149_1904 ();
 FILLCELL_X32 FILLER_149_1936 ();
 FILLCELL_X32 FILLER_149_1968 ();
 FILLCELL_X32 FILLER_149_2000 ();
 FILLCELL_X32 FILLER_149_2032 ();
 FILLCELL_X32 FILLER_149_2064 ();
 FILLCELL_X32 FILLER_149_2096 ();
 FILLCELL_X32 FILLER_149_2128 ();
 FILLCELL_X32 FILLER_149_2160 ();
 FILLCELL_X32 FILLER_149_2192 ();
 FILLCELL_X32 FILLER_149_2224 ();
 FILLCELL_X32 FILLER_149_2256 ();
 FILLCELL_X32 FILLER_149_2288 ();
 FILLCELL_X32 FILLER_149_2320 ();
 FILLCELL_X32 FILLER_149_2352 ();
 FILLCELL_X32 FILLER_149_2384 ();
 FILLCELL_X16 FILLER_149_2416 ();
 FILLCELL_X4 FILLER_149_2432 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X32 FILLER_150_1592 ();
 FILLCELL_X32 FILLER_150_1624 ();
 FILLCELL_X32 FILLER_150_1656 ();
 FILLCELL_X32 FILLER_150_1688 ();
 FILLCELL_X32 FILLER_150_1720 ();
 FILLCELL_X32 FILLER_150_1752 ();
 FILLCELL_X32 FILLER_150_1784 ();
 FILLCELL_X32 FILLER_150_1816 ();
 FILLCELL_X32 FILLER_150_1848 ();
 FILLCELL_X8 FILLER_150_1880 ();
 FILLCELL_X4 FILLER_150_1888 ();
 FILLCELL_X2 FILLER_150_1892 ();
 FILLCELL_X32 FILLER_150_1895 ();
 FILLCELL_X32 FILLER_150_1927 ();
 FILLCELL_X32 FILLER_150_1959 ();
 FILLCELL_X32 FILLER_150_1991 ();
 FILLCELL_X32 FILLER_150_2023 ();
 FILLCELL_X32 FILLER_150_2055 ();
 FILLCELL_X32 FILLER_150_2087 ();
 FILLCELL_X32 FILLER_150_2119 ();
 FILLCELL_X32 FILLER_150_2151 ();
 FILLCELL_X32 FILLER_150_2183 ();
 FILLCELL_X32 FILLER_150_2215 ();
 FILLCELL_X32 FILLER_150_2247 ();
 FILLCELL_X32 FILLER_150_2279 ();
 FILLCELL_X32 FILLER_150_2311 ();
 FILLCELL_X32 FILLER_150_2343 ();
 FILLCELL_X32 FILLER_150_2375 ();
 FILLCELL_X16 FILLER_150_2407 ();
 FILLCELL_X8 FILLER_150_2423 ();
 FILLCELL_X4 FILLER_150_2431 ();
 FILLCELL_X1 FILLER_150_2435 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X32 FILLER_151_1776 ();
 FILLCELL_X32 FILLER_151_1808 ();
 FILLCELL_X32 FILLER_151_1840 ();
 FILLCELL_X32 FILLER_151_1872 ();
 FILLCELL_X32 FILLER_151_1904 ();
 FILLCELL_X32 FILLER_151_1936 ();
 FILLCELL_X32 FILLER_151_1968 ();
 FILLCELL_X32 FILLER_151_2000 ();
 FILLCELL_X32 FILLER_151_2032 ();
 FILLCELL_X32 FILLER_151_2064 ();
 FILLCELL_X32 FILLER_151_2096 ();
 FILLCELL_X32 FILLER_151_2128 ();
 FILLCELL_X32 FILLER_151_2160 ();
 FILLCELL_X32 FILLER_151_2192 ();
 FILLCELL_X32 FILLER_151_2224 ();
 FILLCELL_X32 FILLER_151_2256 ();
 FILLCELL_X32 FILLER_151_2288 ();
 FILLCELL_X32 FILLER_151_2320 ();
 FILLCELL_X32 FILLER_151_2352 ();
 FILLCELL_X32 FILLER_151_2384 ();
 FILLCELL_X16 FILLER_151_2416 ();
 FILLCELL_X4 FILLER_151_2432 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X32 FILLER_152_1624 ();
 FILLCELL_X32 FILLER_152_1656 ();
 FILLCELL_X32 FILLER_152_1688 ();
 FILLCELL_X32 FILLER_152_1720 ();
 FILLCELL_X32 FILLER_152_1752 ();
 FILLCELL_X32 FILLER_152_1784 ();
 FILLCELL_X32 FILLER_152_1816 ();
 FILLCELL_X32 FILLER_152_1848 ();
 FILLCELL_X8 FILLER_152_1880 ();
 FILLCELL_X4 FILLER_152_1888 ();
 FILLCELL_X2 FILLER_152_1892 ();
 FILLCELL_X32 FILLER_152_1895 ();
 FILLCELL_X32 FILLER_152_1927 ();
 FILLCELL_X32 FILLER_152_1959 ();
 FILLCELL_X32 FILLER_152_1991 ();
 FILLCELL_X32 FILLER_152_2023 ();
 FILLCELL_X32 FILLER_152_2055 ();
 FILLCELL_X32 FILLER_152_2087 ();
 FILLCELL_X32 FILLER_152_2119 ();
 FILLCELL_X32 FILLER_152_2151 ();
 FILLCELL_X32 FILLER_152_2183 ();
 FILLCELL_X32 FILLER_152_2215 ();
 FILLCELL_X32 FILLER_152_2247 ();
 FILLCELL_X32 FILLER_152_2279 ();
 FILLCELL_X32 FILLER_152_2311 ();
 FILLCELL_X32 FILLER_152_2343 ();
 FILLCELL_X32 FILLER_152_2375 ();
 FILLCELL_X16 FILLER_152_2407 ();
 FILLCELL_X8 FILLER_152_2423 ();
 FILLCELL_X4 FILLER_152_2431 ();
 FILLCELL_X1 FILLER_152_2435 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X32 FILLER_153_1776 ();
 FILLCELL_X32 FILLER_153_1808 ();
 FILLCELL_X32 FILLER_153_1840 ();
 FILLCELL_X32 FILLER_153_1872 ();
 FILLCELL_X32 FILLER_153_1904 ();
 FILLCELL_X32 FILLER_153_1936 ();
 FILLCELL_X32 FILLER_153_1968 ();
 FILLCELL_X32 FILLER_153_2000 ();
 FILLCELL_X32 FILLER_153_2032 ();
 FILLCELL_X32 FILLER_153_2064 ();
 FILLCELL_X32 FILLER_153_2096 ();
 FILLCELL_X32 FILLER_153_2128 ();
 FILLCELL_X32 FILLER_153_2160 ();
 FILLCELL_X32 FILLER_153_2192 ();
 FILLCELL_X32 FILLER_153_2224 ();
 FILLCELL_X32 FILLER_153_2256 ();
 FILLCELL_X32 FILLER_153_2288 ();
 FILLCELL_X32 FILLER_153_2320 ();
 FILLCELL_X32 FILLER_153_2352 ();
 FILLCELL_X32 FILLER_153_2384 ();
 FILLCELL_X16 FILLER_153_2416 ();
 FILLCELL_X4 FILLER_153_2432 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X32 FILLER_154_1592 ();
 FILLCELL_X32 FILLER_154_1624 ();
 FILLCELL_X32 FILLER_154_1656 ();
 FILLCELL_X32 FILLER_154_1688 ();
 FILLCELL_X32 FILLER_154_1720 ();
 FILLCELL_X32 FILLER_154_1752 ();
 FILLCELL_X32 FILLER_154_1784 ();
 FILLCELL_X32 FILLER_154_1816 ();
 FILLCELL_X32 FILLER_154_1848 ();
 FILLCELL_X8 FILLER_154_1880 ();
 FILLCELL_X4 FILLER_154_1888 ();
 FILLCELL_X2 FILLER_154_1892 ();
 FILLCELL_X32 FILLER_154_1895 ();
 FILLCELL_X32 FILLER_154_1927 ();
 FILLCELL_X32 FILLER_154_1959 ();
 FILLCELL_X32 FILLER_154_1991 ();
 FILLCELL_X32 FILLER_154_2023 ();
 FILLCELL_X32 FILLER_154_2055 ();
 FILLCELL_X32 FILLER_154_2087 ();
 FILLCELL_X32 FILLER_154_2119 ();
 FILLCELL_X32 FILLER_154_2151 ();
 FILLCELL_X32 FILLER_154_2183 ();
 FILLCELL_X32 FILLER_154_2215 ();
 FILLCELL_X32 FILLER_154_2247 ();
 FILLCELL_X32 FILLER_154_2279 ();
 FILLCELL_X32 FILLER_154_2311 ();
 FILLCELL_X32 FILLER_154_2343 ();
 FILLCELL_X32 FILLER_154_2375 ();
 FILLCELL_X16 FILLER_154_2407 ();
 FILLCELL_X8 FILLER_154_2423 ();
 FILLCELL_X4 FILLER_154_2431 ();
 FILLCELL_X1 FILLER_154_2435 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X32 FILLER_155_1776 ();
 FILLCELL_X32 FILLER_155_1808 ();
 FILLCELL_X32 FILLER_155_1840 ();
 FILLCELL_X32 FILLER_155_1872 ();
 FILLCELL_X32 FILLER_155_1904 ();
 FILLCELL_X32 FILLER_155_1936 ();
 FILLCELL_X32 FILLER_155_1968 ();
 FILLCELL_X32 FILLER_155_2000 ();
 FILLCELL_X32 FILLER_155_2032 ();
 FILLCELL_X32 FILLER_155_2064 ();
 FILLCELL_X32 FILLER_155_2096 ();
 FILLCELL_X32 FILLER_155_2128 ();
 FILLCELL_X32 FILLER_155_2160 ();
 FILLCELL_X32 FILLER_155_2192 ();
 FILLCELL_X32 FILLER_155_2224 ();
 FILLCELL_X32 FILLER_155_2256 ();
 FILLCELL_X32 FILLER_155_2288 ();
 FILLCELL_X32 FILLER_155_2320 ();
 FILLCELL_X32 FILLER_155_2352 ();
 FILLCELL_X32 FILLER_155_2384 ();
 FILLCELL_X16 FILLER_155_2416 ();
 FILLCELL_X4 FILLER_155_2432 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X32 FILLER_156_1592 ();
 FILLCELL_X32 FILLER_156_1624 ();
 FILLCELL_X32 FILLER_156_1656 ();
 FILLCELL_X32 FILLER_156_1688 ();
 FILLCELL_X32 FILLER_156_1720 ();
 FILLCELL_X32 FILLER_156_1752 ();
 FILLCELL_X32 FILLER_156_1784 ();
 FILLCELL_X32 FILLER_156_1816 ();
 FILLCELL_X32 FILLER_156_1848 ();
 FILLCELL_X8 FILLER_156_1880 ();
 FILLCELL_X4 FILLER_156_1888 ();
 FILLCELL_X2 FILLER_156_1892 ();
 FILLCELL_X32 FILLER_156_1895 ();
 FILLCELL_X32 FILLER_156_1927 ();
 FILLCELL_X32 FILLER_156_1959 ();
 FILLCELL_X32 FILLER_156_1991 ();
 FILLCELL_X32 FILLER_156_2023 ();
 FILLCELL_X32 FILLER_156_2055 ();
 FILLCELL_X32 FILLER_156_2087 ();
 FILLCELL_X32 FILLER_156_2119 ();
 FILLCELL_X32 FILLER_156_2151 ();
 FILLCELL_X32 FILLER_156_2183 ();
 FILLCELL_X32 FILLER_156_2215 ();
 FILLCELL_X32 FILLER_156_2247 ();
 FILLCELL_X32 FILLER_156_2279 ();
 FILLCELL_X32 FILLER_156_2311 ();
 FILLCELL_X32 FILLER_156_2343 ();
 FILLCELL_X32 FILLER_156_2375 ();
 FILLCELL_X16 FILLER_156_2407 ();
 FILLCELL_X8 FILLER_156_2423 ();
 FILLCELL_X4 FILLER_156_2431 ();
 FILLCELL_X1 FILLER_156_2435 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X32 FILLER_157_1776 ();
 FILLCELL_X32 FILLER_157_1808 ();
 FILLCELL_X32 FILLER_157_1840 ();
 FILLCELL_X32 FILLER_157_1872 ();
 FILLCELL_X32 FILLER_157_1904 ();
 FILLCELL_X32 FILLER_157_1936 ();
 FILLCELL_X32 FILLER_157_1968 ();
 FILLCELL_X32 FILLER_157_2000 ();
 FILLCELL_X32 FILLER_157_2032 ();
 FILLCELL_X32 FILLER_157_2064 ();
 FILLCELL_X32 FILLER_157_2096 ();
 FILLCELL_X32 FILLER_157_2128 ();
 FILLCELL_X32 FILLER_157_2160 ();
 FILLCELL_X32 FILLER_157_2192 ();
 FILLCELL_X32 FILLER_157_2224 ();
 FILLCELL_X32 FILLER_157_2256 ();
 FILLCELL_X32 FILLER_157_2288 ();
 FILLCELL_X32 FILLER_157_2320 ();
 FILLCELL_X32 FILLER_157_2352 ();
 FILLCELL_X32 FILLER_157_2384 ();
 FILLCELL_X16 FILLER_157_2416 ();
 FILLCELL_X4 FILLER_157_2432 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X32 FILLER_158_1592 ();
 FILLCELL_X32 FILLER_158_1624 ();
 FILLCELL_X32 FILLER_158_1656 ();
 FILLCELL_X32 FILLER_158_1688 ();
 FILLCELL_X32 FILLER_158_1720 ();
 FILLCELL_X32 FILLER_158_1752 ();
 FILLCELL_X32 FILLER_158_1784 ();
 FILLCELL_X32 FILLER_158_1816 ();
 FILLCELL_X32 FILLER_158_1848 ();
 FILLCELL_X8 FILLER_158_1880 ();
 FILLCELL_X4 FILLER_158_1888 ();
 FILLCELL_X2 FILLER_158_1892 ();
 FILLCELL_X32 FILLER_158_1895 ();
 FILLCELL_X32 FILLER_158_1927 ();
 FILLCELL_X32 FILLER_158_1959 ();
 FILLCELL_X32 FILLER_158_1991 ();
 FILLCELL_X32 FILLER_158_2023 ();
 FILLCELL_X32 FILLER_158_2055 ();
 FILLCELL_X32 FILLER_158_2087 ();
 FILLCELL_X32 FILLER_158_2119 ();
 FILLCELL_X32 FILLER_158_2151 ();
 FILLCELL_X32 FILLER_158_2183 ();
 FILLCELL_X32 FILLER_158_2215 ();
 FILLCELL_X32 FILLER_158_2247 ();
 FILLCELL_X32 FILLER_158_2279 ();
 FILLCELL_X32 FILLER_158_2311 ();
 FILLCELL_X32 FILLER_158_2343 ();
 FILLCELL_X32 FILLER_158_2375 ();
 FILLCELL_X16 FILLER_158_2407 ();
 FILLCELL_X8 FILLER_158_2423 ();
 FILLCELL_X4 FILLER_158_2431 ();
 FILLCELL_X1 FILLER_158_2435 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X32 FILLER_159_1776 ();
 FILLCELL_X32 FILLER_159_1808 ();
 FILLCELL_X32 FILLER_159_1840 ();
 FILLCELL_X32 FILLER_159_1872 ();
 FILLCELL_X32 FILLER_159_1904 ();
 FILLCELL_X32 FILLER_159_1936 ();
 FILLCELL_X32 FILLER_159_1968 ();
 FILLCELL_X32 FILLER_159_2000 ();
 FILLCELL_X32 FILLER_159_2032 ();
 FILLCELL_X32 FILLER_159_2064 ();
 FILLCELL_X32 FILLER_159_2096 ();
 FILLCELL_X32 FILLER_159_2128 ();
 FILLCELL_X32 FILLER_159_2160 ();
 FILLCELL_X32 FILLER_159_2192 ();
 FILLCELL_X32 FILLER_159_2224 ();
 FILLCELL_X32 FILLER_159_2256 ();
 FILLCELL_X32 FILLER_159_2288 ();
 FILLCELL_X32 FILLER_159_2320 ();
 FILLCELL_X32 FILLER_159_2352 ();
 FILLCELL_X32 FILLER_159_2384 ();
 FILLCELL_X16 FILLER_159_2416 ();
 FILLCELL_X4 FILLER_159_2432 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X32 FILLER_160_1592 ();
 FILLCELL_X32 FILLER_160_1624 ();
 FILLCELL_X32 FILLER_160_1656 ();
 FILLCELL_X32 FILLER_160_1688 ();
 FILLCELL_X32 FILLER_160_1720 ();
 FILLCELL_X32 FILLER_160_1752 ();
 FILLCELL_X32 FILLER_160_1784 ();
 FILLCELL_X32 FILLER_160_1816 ();
 FILLCELL_X32 FILLER_160_1848 ();
 FILLCELL_X8 FILLER_160_1880 ();
 FILLCELL_X4 FILLER_160_1888 ();
 FILLCELL_X2 FILLER_160_1892 ();
 FILLCELL_X32 FILLER_160_1895 ();
 FILLCELL_X32 FILLER_160_1927 ();
 FILLCELL_X32 FILLER_160_1959 ();
 FILLCELL_X32 FILLER_160_1991 ();
 FILLCELL_X32 FILLER_160_2023 ();
 FILLCELL_X32 FILLER_160_2055 ();
 FILLCELL_X32 FILLER_160_2087 ();
 FILLCELL_X32 FILLER_160_2119 ();
 FILLCELL_X32 FILLER_160_2151 ();
 FILLCELL_X32 FILLER_160_2183 ();
 FILLCELL_X32 FILLER_160_2215 ();
 FILLCELL_X32 FILLER_160_2247 ();
 FILLCELL_X32 FILLER_160_2279 ();
 FILLCELL_X32 FILLER_160_2311 ();
 FILLCELL_X32 FILLER_160_2343 ();
 FILLCELL_X32 FILLER_160_2375 ();
 FILLCELL_X16 FILLER_160_2407 ();
 FILLCELL_X8 FILLER_160_2423 ();
 FILLCELL_X4 FILLER_160_2431 ();
 FILLCELL_X1 FILLER_160_2435 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X32 FILLER_161_1584 ();
 FILLCELL_X32 FILLER_161_1616 ();
 FILLCELL_X32 FILLER_161_1648 ();
 FILLCELL_X32 FILLER_161_1680 ();
 FILLCELL_X32 FILLER_161_1712 ();
 FILLCELL_X32 FILLER_161_1744 ();
 FILLCELL_X32 FILLER_161_1776 ();
 FILLCELL_X32 FILLER_161_1808 ();
 FILLCELL_X32 FILLER_161_1840 ();
 FILLCELL_X32 FILLER_161_1872 ();
 FILLCELL_X32 FILLER_161_1904 ();
 FILLCELL_X32 FILLER_161_1936 ();
 FILLCELL_X32 FILLER_161_1968 ();
 FILLCELL_X32 FILLER_161_2000 ();
 FILLCELL_X32 FILLER_161_2032 ();
 FILLCELL_X32 FILLER_161_2064 ();
 FILLCELL_X32 FILLER_161_2096 ();
 FILLCELL_X32 FILLER_161_2128 ();
 FILLCELL_X32 FILLER_161_2160 ();
 FILLCELL_X32 FILLER_161_2192 ();
 FILLCELL_X32 FILLER_161_2224 ();
 FILLCELL_X32 FILLER_161_2256 ();
 FILLCELL_X32 FILLER_161_2288 ();
 FILLCELL_X32 FILLER_161_2320 ();
 FILLCELL_X32 FILLER_161_2352 ();
 FILLCELL_X32 FILLER_161_2384 ();
 FILLCELL_X16 FILLER_161_2416 ();
 FILLCELL_X4 FILLER_161_2432 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1304 ();
 FILLCELL_X32 FILLER_162_1336 ();
 FILLCELL_X32 FILLER_162_1368 ();
 FILLCELL_X32 FILLER_162_1400 ();
 FILLCELL_X32 FILLER_162_1432 ();
 FILLCELL_X32 FILLER_162_1464 ();
 FILLCELL_X32 FILLER_162_1496 ();
 FILLCELL_X32 FILLER_162_1528 ();
 FILLCELL_X32 FILLER_162_1560 ();
 FILLCELL_X32 FILLER_162_1592 ();
 FILLCELL_X32 FILLER_162_1624 ();
 FILLCELL_X32 FILLER_162_1656 ();
 FILLCELL_X32 FILLER_162_1688 ();
 FILLCELL_X32 FILLER_162_1720 ();
 FILLCELL_X32 FILLER_162_1752 ();
 FILLCELL_X32 FILLER_162_1784 ();
 FILLCELL_X32 FILLER_162_1816 ();
 FILLCELL_X32 FILLER_162_1848 ();
 FILLCELL_X8 FILLER_162_1880 ();
 FILLCELL_X4 FILLER_162_1888 ();
 FILLCELL_X2 FILLER_162_1892 ();
 FILLCELL_X32 FILLER_162_1895 ();
 FILLCELL_X32 FILLER_162_1927 ();
 FILLCELL_X32 FILLER_162_1959 ();
 FILLCELL_X32 FILLER_162_1991 ();
 FILLCELL_X32 FILLER_162_2023 ();
 FILLCELL_X32 FILLER_162_2055 ();
 FILLCELL_X32 FILLER_162_2087 ();
 FILLCELL_X32 FILLER_162_2119 ();
 FILLCELL_X32 FILLER_162_2151 ();
 FILLCELL_X32 FILLER_162_2183 ();
 FILLCELL_X32 FILLER_162_2215 ();
 FILLCELL_X32 FILLER_162_2247 ();
 FILLCELL_X32 FILLER_162_2279 ();
 FILLCELL_X32 FILLER_162_2311 ();
 FILLCELL_X32 FILLER_162_2343 ();
 FILLCELL_X32 FILLER_162_2375 ();
 FILLCELL_X16 FILLER_162_2407 ();
 FILLCELL_X8 FILLER_162_2423 ();
 FILLCELL_X4 FILLER_162_2431 ();
 FILLCELL_X1 FILLER_162_2435 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X32 FILLER_163_1648 ();
 FILLCELL_X32 FILLER_163_1680 ();
 FILLCELL_X32 FILLER_163_1712 ();
 FILLCELL_X32 FILLER_163_1744 ();
 FILLCELL_X32 FILLER_163_1776 ();
 FILLCELL_X32 FILLER_163_1808 ();
 FILLCELL_X32 FILLER_163_1840 ();
 FILLCELL_X32 FILLER_163_1872 ();
 FILLCELL_X32 FILLER_163_1904 ();
 FILLCELL_X32 FILLER_163_1936 ();
 FILLCELL_X32 FILLER_163_1968 ();
 FILLCELL_X32 FILLER_163_2000 ();
 FILLCELL_X32 FILLER_163_2032 ();
 FILLCELL_X32 FILLER_163_2064 ();
 FILLCELL_X32 FILLER_163_2096 ();
 FILLCELL_X32 FILLER_163_2128 ();
 FILLCELL_X32 FILLER_163_2160 ();
 FILLCELL_X32 FILLER_163_2192 ();
 FILLCELL_X32 FILLER_163_2224 ();
 FILLCELL_X32 FILLER_163_2256 ();
 FILLCELL_X32 FILLER_163_2288 ();
 FILLCELL_X32 FILLER_163_2320 ();
 FILLCELL_X32 FILLER_163_2352 ();
 FILLCELL_X32 FILLER_163_2384 ();
 FILLCELL_X16 FILLER_163_2416 ();
 FILLCELL_X4 FILLER_163_2432 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X32 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1336 ();
 FILLCELL_X32 FILLER_164_1368 ();
 FILLCELL_X32 FILLER_164_1400 ();
 FILLCELL_X32 FILLER_164_1432 ();
 FILLCELL_X32 FILLER_164_1464 ();
 FILLCELL_X32 FILLER_164_1496 ();
 FILLCELL_X32 FILLER_164_1528 ();
 FILLCELL_X32 FILLER_164_1560 ();
 FILLCELL_X32 FILLER_164_1592 ();
 FILLCELL_X32 FILLER_164_1624 ();
 FILLCELL_X32 FILLER_164_1656 ();
 FILLCELL_X32 FILLER_164_1688 ();
 FILLCELL_X32 FILLER_164_1720 ();
 FILLCELL_X32 FILLER_164_1752 ();
 FILLCELL_X32 FILLER_164_1784 ();
 FILLCELL_X32 FILLER_164_1816 ();
 FILLCELL_X32 FILLER_164_1848 ();
 FILLCELL_X8 FILLER_164_1880 ();
 FILLCELL_X4 FILLER_164_1888 ();
 FILLCELL_X2 FILLER_164_1892 ();
 FILLCELL_X32 FILLER_164_1895 ();
 FILLCELL_X32 FILLER_164_1927 ();
 FILLCELL_X32 FILLER_164_1959 ();
 FILLCELL_X32 FILLER_164_1991 ();
 FILLCELL_X32 FILLER_164_2023 ();
 FILLCELL_X32 FILLER_164_2055 ();
 FILLCELL_X32 FILLER_164_2087 ();
 FILLCELL_X32 FILLER_164_2119 ();
 FILLCELL_X32 FILLER_164_2151 ();
 FILLCELL_X32 FILLER_164_2183 ();
 FILLCELL_X32 FILLER_164_2215 ();
 FILLCELL_X32 FILLER_164_2247 ();
 FILLCELL_X32 FILLER_164_2279 ();
 FILLCELL_X32 FILLER_164_2311 ();
 FILLCELL_X32 FILLER_164_2343 ();
 FILLCELL_X32 FILLER_164_2375 ();
 FILLCELL_X16 FILLER_164_2407 ();
 FILLCELL_X8 FILLER_164_2423 ();
 FILLCELL_X4 FILLER_164_2431 ();
 FILLCELL_X1 FILLER_164_2435 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X32 FILLER_165_1648 ();
 FILLCELL_X32 FILLER_165_1680 ();
 FILLCELL_X32 FILLER_165_1712 ();
 FILLCELL_X32 FILLER_165_1744 ();
 FILLCELL_X32 FILLER_165_1776 ();
 FILLCELL_X32 FILLER_165_1808 ();
 FILLCELL_X32 FILLER_165_1840 ();
 FILLCELL_X32 FILLER_165_1872 ();
 FILLCELL_X32 FILLER_165_1904 ();
 FILLCELL_X32 FILLER_165_1936 ();
 FILLCELL_X32 FILLER_165_1968 ();
 FILLCELL_X32 FILLER_165_2000 ();
 FILLCELL_X32 FILLER_165_2032 ();
 FILLCELL_X32 FILLER_165_2064 ();
 FILLCELL_X32 FILLER_165_2096 ();
 FILLCELL_X32 FILLER_165_2128 ();
 FILLCELL_X32 FILLER_165_2160 ();
 FILLCELL_X32 FILLER_165_2192 ();
 FILLCELL_X32 FILLER_165_2224 ();
 FILLCELL_X32 FILLER_165_2256 ();
 FILLCELL_X32 FILLER_165_2288 ();
 FILLCELL_X32 FILLER_165_2320 ();
 FILLCELL_X32 FILLER_165_2352 ();
 FILLCELL_X32 FILLER_165_2384 ();
 FILLCELL_X16 FILLER_165_2416 ();
 FILLCELL_X4 FILLER_165_2432 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X32 FILLER_166_1112 ();
 FILLCELL_X32 FILLER_166_1144 ();
 FILLCELL_X32 FILLER_166_1176 ();
 FILLCELL_X32 FILLER_166_1208 ();
 FILLCELL_X32 FILLER_166_1240 ();
 FILLCELL_X32 FILLER_166_1272 ();
 FILLCELL_X32 FILLER_166_1304 ();
 FILLCELL_X32 FILLER_166_1336 ();
 FILLCELL_X32 FILLER_166_1368 ();
 FILLCELL_X32 FILLER_166_1400 ();
 FILLCELL_X32 FILLER_166_1432 ();
 FILLCELL_X32 FILLER_166_1464 ();
 FILLCELL_X32 FILLER_166_1496 ();
 FILLCELL_X32 FILLER_166_1528 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X32 FILLER_166_1592 ();
 FILLCELL_X32 FILLER_166_1624 ();
 FILLCELL_X32 FILLER_166_1656 ();
 FILLCELL_X32 FILLER_166_1688 ();
 FILLCELL_X32 FILLER_166_1720 ();
 FILLCELL_X32 FILLER_166_1752 ();
 FILLCELL_X32 FILLER_166_1784 ();
 FILLCELL_X32 FILLER_166_1816 ();
 FILLCELL_X32 FILLER_166_1848 ();
 FILLCELL_X8 FILLER_166_1880 ();
 FILLCELL_X4 FILLER_166_1888 ();
 FILLCELL_X2 FILLER_166_1892 ();
 FILLCELL_X32 FILLER_166_1895 ();
 FILLCELL_X32 FILLER_166_1927 ();
 FILLCELL_X32 FILLER_166_1959 ();
 FILLCELL_X32 FILLER_166_1991 ();
 FILLCELL_X32 FILLER_166_2023 ();
 FILLCELL_X32 FILLER_166_2055 ();
 FILLCELL_X32 FILLER_166_2087 ();
 FILLCELL_X32 FILLER_166_2119 ();
 FILLCELL_X32 FILLER_166_2151 ();
 FILLCELL_X32 FILLER_166_2183 ();
 FILLCELL_X32 FILLER_166_2215 ();
 FILLCELL_X32 FILLER_166_2247 ();
 FILLCELL_X32 FILLER_166_2279 ();
 FILLCELL_X32 FILLER_166_2311 ();
 FILLCELL_X32 FILLER_166_2343 ();
 FILLCELL_X32 FILLER_166_2375 ();
 FILLCELL_X16 FILLER_166_2407 ();
 FILLCELL_X8 FILLER_166_2423 ();
 FILLCELL_X4 FILLER_166_2431 ();
 FILLCELL_X1 FILLER_166_2435 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X32 FILLER_167_1648 ();
 FILLCELL_X32 FILLER_167_1680 ();
 FILLCELL_X32 FILLER_167_1712 ();
 FILLCELL_X32 FILLER_167_1744 ();
 FILLCELL_X32 FILLER_167_1776 ();
 FILLCELL_X32 FILLER_167_1808 ();
 FILLCELL_X32 FILLER_167_1840 ();
 FILLCELL_X32 FILLER_167_1872 ();
 FILLCELL_X32 FILLER_167_1904 ();
 FILLCELL_X32 FILLER_167_1936 ();
 FILLCELL_X32 FILLER_167_1968 ();
 FILLCELL_X32 FILLER_167_2000 ();
 FILLCELL_X32 FILLER_167_2032 ();
 FILLCELL_X32 FILLER_167_2064 ();
 FILLCELL_X32 FILLER_167_2096 ();
 FILLCELL_X32 FILLER_167_2128 ();
 FILLCELL_X32 FILLER_167_2160 ();
 FILLCELL_X32 FILLER_167_2192 ();
 FILLCELL_X32 FILLER_167_2224 ();
 FILLCELL_X32 FILLER_167_2256 ();
 FILLCELL_X32 FILLER_167_2288 ();
 FILLCELL_X32 FILLER_167_2320 ();
 FILLCELL_X32 FILLER_167_2352 ();
 FILLCELL_X32 FILLER_167_2384 ();
 FILLCELL_X16 FILLER_167_2416 ();
 FILLCELL_X4 FILLER_167_2432 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X32 FILLER_168_1304 ();
 FILLCELL_X32 FILLER_168_1336 ();
 FILLCELL_X32 FILLER_168_1368 ();
 FILLCELL_X32 FILLER_168_1400 ();
 FILLCELL_X32 FILLER_168_1432 ();
 FILLCELL_X32 FILLER_168_1464 ();
 FILLCELL_X32 FILLER_168_1496 ();
 FILLCELL_X32 FILLER_168_1528 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X32 FILLER_168_1592 ();
 FILLCELL_X32 FILLER_168_1624 ();
 FILLCELL_X32 FILLER_168_1656 ();
 FILLCELL_X32 FILLER_168_1688 ();
 FILLCELL_X32 FILLER_168_1720 ();
 FILLCELL_X32 FILLER_168_1752 ();
 FILLCELL_X32 FILLER_168_1784 ();
 FILLCELL_X32 FILLER_168_1816 ();
 FILLCELL_X32 FILLER_168_1848 ();
 FILLCELL_X8 FILLER_168_1880 ();
 FILLCELL_X4 FILLER_168_1888 ();
 FILLCELL_X2 FILLER_168_1892 ();
 FILLCELL_X32 FILLER_168_1895 ();
 FILLCELL_X32 FILLER_168_1927 ();
 FILLCELL_X32 FILLER_168_1959 ();
 FILLCELL_X32 FILLER_168_1991 ();
 FILLCELL_X32 FILLER_168_2023 ();
 FILLCELL_X32 FILLER_168_2055 ();
 FILLCELL_X32 FILLER_168_2087 ();
 FILLCELL_X32 FILLER_168_2119 ();
 FILLCELL_X32 FILLER_168_2151 ();
 FILLCELL_X32 FILLER_168_2183 ();
 FILLCELL_X32 FILLER_168_2215 ();
 FILLCELL_X32 FILLER_168_2247 ();
 FILLCELL_X32 FILLER_168_2279 ();
 FILLCELL_X32 FILLER_168_2311 ();
 FILLCELL_X32 FILLER_168_2343 ();
 FILLCELL_X32 FILLER_168_2375 ();
 FILLCELL_X16 FILLER_168_2407 ();
 FILLCELL_X8 FILLER_168_2423 ();
 FILLCELL_X4 FILLER_168_2431 ();
 FILLCELL_X1 FILLER_168_2435 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X32 FILLER_169_1089 ();
 FILLCELL_X32 FILLER_169_1121 ();
 FILLCELL_X32 FILLER_169_1153 ();
 FILLCELL_X32 FILLER_169_1185 ();
 FILLCELL_X32 FILLER_169_1217 ();
 FILLCELL_X8 FILLER_169_1249 ();
 FILLCELL_X4 FILLER_169_1257 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X32 FILLER_169_1648 ();
 FILLCELL_X32 FILLER_169_1680 ();
 FILLCELL_X32 FILLER_169_1712 ();
 FILLCELL_X32 FILLER_169_1744 ();
 FILLCELL_X32 FILLER_169_1776 ();
 FILLCELL_X32 FILLER_169_1808 ();
 FILLCELL_X32 FILLER_169_1840 ();
 FILLCELL_X32 FILLER_169_1872 ();
 FILLCELL_X32 FILLER_169_1904 ();
 FILLCELL_X32 FILLER_169_1936 ();
 FILLCELL_X32 FILLER_169_1968 ();
 FILLCELL_X32 FILLER_169_2000 ();
 FILLCELL_X32 FILLER_169_2032 ();
 FILLCELL_X32 FILLER_169_2064 ();
 FILLCELL_X32 FILLER_169_2096 ();
 FILLCELL_X32 FILLER_169_2128 ();
 FILLCELL_X32 FILLER_169_2160 ();
 FILLCELL_X32 FILLER_169_2192 ();
 FILLCELL_X32 FILLER_169_2224 ();
 FILLCELL_X32 FILLER_169_2256 ();
 FILLCELL_X32 FILLER_169_2288 ();
 FILLCELL_X32 FILLER_169_2320 ();
 FILLCELL_X32 FILLER_169_2352 ();
 FILLCELL_X32 FILLER_169_2384 ();
 FILLCELL_X16 FILLER_169_2416 ();
 FILLCELL_X4 FILLER_169_2432 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X32 FILLER_170_1080 ();
 FILLCELL_X32 FILLER_170_1112 ();
 FILLCELL_X32 FILLER_170_1144 ();
 FILLCELL_X32 FILLER_170_1176 ();
 FILLCELL_X32 FILLER_170_1208 ();
 FILLCELL_X32 FILLER_170_1240 ();
 FILLCELL_X32 FILLER_170_1272 ();
 FILLCELL_X32 FILLER_170_1304 ();
 FILLCELL_X32 FILLER_170_1336 ();
 FILLCELL_X32 FILLER_170_1368 ();
 FILLCELL_X32 FILLER_170_1400 ();
 FILLCELL_X32 FILLER_170_1432 ();
 FILLCELL_X32 FILLER_170_1464 ();
 FILLCELL_X32 FILLER_170_1496 ();
 FILLCELL_X32 FILLER_170_1528 ();
 FILLCELL_X32 FILLER_170_1560 ();
 FILLCELL_X32 FILLER_170_1592 ();
 FILLCELL_X32 FILLER_170_1624 ();
 FILLCELL_X32 FILLER_170_1656 ();
 FILLCELL_X32 FILLER_170_1688 ();
 FILLCELL_X32 FILLER_170_1720 ();
 FILLCELL_X32 FILLER_170_1752 ();
 FILLCELL_X32 FILLER_170_1784 ();
 FILLCELL_X32 FILLER_170_1816 ();
 FILLCELL_X32 FILLER_170_1848 ();
 FILLCELL_X8 FILLER_170_1880 ();
 FILLCELL_X4 FILLER_170_1888 ();
 FILLCELL_X2 FILLER_170_1892 ();
 FILLCELL_X32 FILLER_170_1895 ();
 FILLCELL_X32 FILLER_170_1927 ();
 FILLCELL_X32 FILLER_170_1959 ();
 FILLCELL_X32 FILLER_170_1991 ();
 FILLCELL_X32 FILLER_170_2023 ();
 FILLCELL_X32 FILLER_170_2055 ();
 FILLCELL_X32 FILLER_170_2087 ();
 FILLCELL_X32 FILLER_170_2119 ();
 FILLCELL_X32 FILLER_170_2151 ();
 FILLCELL_X32 FILLER_170_2183 ();
 FILLCELL_X32 FILLER_170_2215 ();
 FILLCELL_X32 FILLER_170_2247 ();
 FILLCELL_X32 FILLER_170_2279 ();
 FILLCELL_X32 FILLER_170_2311 ();
 FILLCELL_X32 FILLER_170_2343 ();
 FILLCELL_X32 FILLER_170_2375 ();
 FILLCELL_X16 FILLER_170_2407 ();
 FILLCELL_X8 FILLER_170_2423 ();
 FILLCELL_X4 FILLER_170_2431 ();
 FILLCELL_X1 FILLER_170_2435 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X32 FILLER_171_1185 ();
 FILLCELL_X32 FILLER_171_1217 ();
 FILLCELL_X8 FILLER_171_1249 ();
 FILLCELL_X4 FILLER_171_1257 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X32 FILLER_171_1648 ();
 FILLCELL_X32 FILLER_171_1680 ();
 FILLCELL_X32 FILLER_171_1712 ();
 FILLCELL_X32 FILLER_171_1744 ();
 FILLCELL_X32 FILLER_171_1776 ();
 FILLCELL_X32 FILLER_171_1808 ();
 FILLCELL_X32 FILLER_171_1840 ();
 FILLCELL_X32 FILLER_171_1872 ();
 FILLCELL_X32 FILLER_171_1904 ();
 FILLCELL_X32 FILLER_171_1936 ();
 FILLCELL_X32 FILLER_171_1968 ();
 FILLCELL_X32 FILLER_171_2000 ();
 FILLCELL_X32 FILLER_171_2032 ();
 FILLCELL_X32 FILLER_171_2064 ();
 FILLCELL_X32 FILLER_171_2096 ();
 FILLCELL_X32 FILLER_171_2128 ();
 FILLCELL_X32 FILLER_171_2160 ();
 FILLCELL_X32 FILLER_171_2192 ();
 FILLCELL_X32 FILLER_171_2224 ();
 FILLCELL_X32 FILLER_171_2256 ();
 FILLCELL_X32 FILLER_171_2288 ();
 FILLCELL_X32 FILLER_171_2320 ();
 FILLCELL_X32 FILLER_171_2352 ();
 FILLCELL_X32 FILLER_171_2384 ();
 FILLCELL_X16 FILLER_171_2416 ();
 FILLCELL_X4 FILLER_171_2432 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X32 FILLER_172_1080 ();
 FILLCELL_X32 FILLER_172_1112 ();
 FILLCELL_X32 FILLER_172_1144 ();
 FILLCELL_X32 FILLER_172_1176 ();
 FILLCELL_X32 FILLER_172_1208 ();
 FILLCELL_X32 FILLER_172_1240 ();
 FILLCELL_X32 FILLER_172_1272 ();
 FILLCELL_X32 FILLER_172_1304 ();
 FILLCELL_X32 FILLER_172_1336 ();
 FILLCELL_X32 FILLER_172_1368 ();
 FILLCELL_X32 FILLER_172_1400 ();
 FILLCELL_X32 FILLER_172_1432 ();
 FILLCELL_X32 FILLER_172_1464 ();
 FILLCELL_X32 FILLER_172_1496 ();
 FILLCELL_X32 FILLER_172_1528 ();
 FILLCELL_X32 FILLER_172_1560 ();
 FILLCELL_X32 FILLER_172_1592 ();
 FILLCELL_X32 FILLER_172_1624 ();
 FILLCELL_X32 FILLER_172_1656 ();
 FILLCELL_X32 FILLER_172_1688 ();
 FILLCELL_X32 FILLER_172_1720 ();
 FILLCELL_X32 FILLER_172_1752 ();
 FILLCELL_X32 FILLER_172_1784 ();
 FILLCELL_X32 FILLER_172_1816 ();
 FILLCELL_X32 FILLER_172_1848 ();
 FILLCELL_X8 FILLER_172_1880 ();
 FILLCELL_X4 FILLER_172_1888 ();
 FILLCELL_X2 FILLER_172_1892 ();
 FILLCELL_X32 FILLER_172_1895 ();
 FILLCELL_X32 FILLER_172_1927 ();
 FILLCELL_X32 FILLER_172_1959 ();
 FILLCELL_X32 FILLER_172_1991 ();
 FILLCELL_X32 FILLER_172_2023 ();
 FILLCELL_X32 FILLER_172_2055 ();
 FILLCELL_X32 FILLER_172_2087 ();
 FILLCELL_X32 FILLER_172_2119 ();
 FILLCELL_X32 FILLER_172_2151 ();
 FILLCELL_X32 FILLER_172_2183 ();
 FILLCELL_X32 FILLER_172_2215 ();
 FILLCELL_X32 FILLER_172_2247 ();
 FILLCELL_X32 FILLER_172_2279 ();
 FILLCELL_X32 FILLER_172_2311 ();
 FILLCELL_X32 FILLER_172_2343 ();
 FILLCELL_X32 FILLER_172_2375 ();
 FILLCELL_X16 FILLER_172_2407 ();
 FILLCELL_X8 FILLER_172_2423 ();
 FILLCELL_X4 FILLER_172_2431 ();
 FILLCELL_X1 FILLER_172_2435 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X32 FILLER_173_1648 ();
 FILLCELL_X32 FILLER_173_1680 ();
 FILLCELL_X32 FILLER_173_1712 ();
 FILLCELL_X32 FILLER_173_1744 ();
 FILLCELL_X32 FILLER_173_1776 ();
 FILLCELL_X32 FILLER_173_1808 ();
 FILLCELL_X32 FILLER_173_1840 ();
 FILLCELL_X32 FILLER_173_1872 ();
 FILLCELL_X32 FILLER_173_1904 ();
 FILLCELL_X32 FILLER_173_1936 ();
 FILLCELL_X32 FILLER_173_1968 ();
 FILLCELL_X32 FILLER_173_2000 ();
 FILLCELL_X32 FILLER_173_2032 ();
 FILLCELL_X32 FILLER_173_2064 ();
 FILLCELL_X32 FILLER_173_2096 ();
 FILLCELL_X32 FILLER_173_2128 ();
 FILLCELL_X32 FILLER_173_2160 ();
 FILLCELL_X32 FILLER_173_2192 ();
 FILLCELL_X32 FILLER_173_2224 ();
 FILLCELL_X32 FILLER_173_2256 ();
 FILLCELL_X32 FILLER_173_2288 ();
 FILLCELL_X32 FILLER_173_2320 ();
 FILLCELL_X32 FILLER_173_2352 ();
 FILLCELL_X32 FILLER_173_2384 ();
 FILLCELL_X16 FILLER_173_2416 ();
 FILLCELL_X4 FILLER_173_2432 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X32 FILLER_174_1592 ();
 FILLCELL_X32 FILLER_174_1624 ();
 FILLCELL_X32 FILLER_174_1656 ();
 FILLCELL_X32 FILLER_174_1688 ();
 FILLCELL_X32 FILLER_174_1720 ();
 FILLCELL_X32 FILLER_174_1752 ();
 FILLCELL_X32 FILLER_174_1784 ();
 FILLCELL_X32 FILLER_174_1816 ();
 FILLCELL_X32 FILLER_174_1848 ();
 FILLCELL_X8 FILLER_174_1880 ();
 FILLCELL_X4 FILLER_174_1888 ();
 FILLCELL_X2 FILLER_174_1892 ();
 FILLCELL_X32 FILLER_174_1895 ();
 FILLCELL_X32 FILLER_174_1927 ();
 FILLCELL_X32 FILLER_174_1959 ();
 FILLCELL_X32 FILLER_174_1991 ();
 FILLCELL_X32 FILLER_174_2023 ();
 FILLCELL_X32 FILLER_174_2055 ();
 FILLCELL_X32 FILLER_174_2087 ();
 FILLCELL_X32 FILLER_174_2119 ();
 FILLCELL_X32 FILLER_174_2151 ();
 FILLCELL_X32 FILLER_174_2183 ();
 FILLCELL_X32 FILLER_174_2215 ();
 FILLCELL_X32 FILLER_174_2247 ();
 FILLCELL_X32 FILLER_174_2279 ();
 FILLCELL_X32 FILLER_174_2311 ();
 FILLCELL_X32 FILLER_174_2343 ();
 FILLCELL_X32 FILLER_174_2375 ();
 FILLCELL_X16 FILLER_174_2407 ();
 FILLCELL_X8 FILLER_174_2423 ();
 FILLCELL_X4 FILLER_174_2431 ();
 FILLCELL_X1 FILLER_174_2435 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1648 ();
 FILLCELL_X32 FILLER_175_1680 ();
 FILLCELL_X32 FILLER_175_1712 ();
 FILLCELL_X32 FILLER_175_1744 ();
 FILLCELL_X32 FILLER_175_1776 ();
 FILLCELL_X32 FILLER_175_1808 ();
 FILLCELL_X32 FILLER_175_1840 ();
 FILLCELL_X32 FILLER_175_1872 ();
 FILLCELL_X32 FILLER_175_1904 ();
 FILLCELL_X32 FILLER_175_1936 ();
 FILLCELL_X32 FILLER_175_1968 ();
 FILLCELL_X32 FILLER_175_2000 ();
 FILLCELL_X32 FILLER_175_2032 ();
 FILLCELL_X32 FILLER_175_2064 ();
 FILLCELL_X32 FILLER_175_2096 ();
 FILLCELL_X32 FILLER_175_2128 ();
 FILLCELL_X32 FILLER_175_2160 ();
 FILLCELL_X32 FILLER_175_2192 ();
 FILLCELL_X32 FILLER_175_2224 ();
 FILLCELL_X32 FILLER_175_2256 ();
 FILLCELL_X32 FILLER_175_2288 ();
 FILLCELL_X32 FILLER_175_2320 ();
 FILLCELL_X32 FILLER_175_2352 ();
 FILLCELL_X32 FILLER_175_2384 ();
 FILLCELL_X16 FILLER_175_2416 ();
 FILLCELL_X4 FILLER_175_2432 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X32 FILLER_176_1304 ();
 FILLCELL_X32 FILLER_176_1336 ();
 FILLCELL_X32 FILLER_176_1368 ();
 FILLCELL_X32 FILLER_176_1400 ();
 FILLCELL_X32 FILLER_176_1432 ();
 FILLCELL_X32 FILLER_176_1464 ();
 FILLCELL_X32 FILLER_176_1496 ();
 FILLCELL_X32 FILLER_176_1528 ();
 FILLCELL_X32 FILLER_176_1560 ();
 FILLCELL_X32 FILLER_176_1592 ();
 FILLCELL_X32 FILLER_176_1624 ();
 FILLCELL_X32 FILLER_176_1656 ();
 FILLCELL_X32 FILLER_176_1688 ();
 FILLCELL_X32 FILLER_176_1720 ();
 FILLCELL_X32 FILLER_176_1752 ();
 FILLCELL_X32 FILLER_176_1784 ();
 FILLCELL_X32 FILLER_176_1816 ();
 FILLCELL_X32 FILLER_176_1848 ();
 FILLCELL_X8 FILLER_176_1880 ();
 FILLCELL_X4 FILLER_176_1888 ();
 FILLCELL_X2 FILLER_176_1892 ();
 FILLCELL_X32 FILLER_176_1895 ();
 FILLCELL_X32 FILLER_176_1927 ();
 FILLCELL_X32 FILLER_176_1959 ();
 FILLCELL_X32 FILLER_176_1991 ();
 FILLCELL_X32 FILLER_176_2023 ();
 FILLCELL_X32 FILLER_176_2055 ();
 FILLCELL_X32 FILLER_176_2087 ();
 FILLCELL_X32 FILLER_176_2119 ();
 FILLCELL_X32 FILLER_176_2151 ();
 FILLCELL_X32 FILLER_176_2183 ();
 FILLCELL_X32 FILLER_176_2215 ();
 FILLCELL_X32 FILLER_176_2247 ();
 FILLCELL_X32 FILLER_176_2279 ();
 FILLCELL_X32 FILLER_176_2311 ();
 FILLCELL_X32 FILLER_176_2343 ();
 FILLCELL_X32 FILLER_176_2375 ();
 FILLCELL_X16 FILLER_176_2407 ();
 FILLCELL_X8 FILLER_176_2423 ();
 FILLCELL_X4 FILLER_176_2431 ();
 FILLCELL_X1 FILLER_176_2435 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X32 FILLER_177_1121 ();
 FILLCELL_X32 FILLER_177_1153 ();
 FILLCELL_X32 FILLER_177_1185 ();
 FILLCELL_X32 FILLER_177_1217 ();
 FILLCELL_X8 FILLER_177_1249 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X32 FILLER_177_1648 ();
 FILLCELL_X32 FILLER_177_1680 ();
 FILLCELL_X32 FILLER_177_1712 ();
 FILLCELL_X32 FILLER_177_1744 ();
 FILLCELL_X32 FILLER_177_1776 ();
 FILLCELL_X32 FILLER_177_1808 ();
 FILLCELL_X32 FILLER_177_1840 ();
 FILLCELL_X32 FILLER_177_1872 ();
 FILLCELL_X32 FILLER_177_1904 ();
 FILLCELL_X32 FILLER_177_1936 ();
 FILLCELL_X32 FILLER_177_1968 ();
 FILLCELL_X32 FILLER_177_2000 ();
 FILLCELL_X32 FILLER_177_2032 ();
 FILLCELL_X32 FILLER_177_2064 ();
 FILLCELL_X32 FILLER_177_2096 ();
 FILLCELL_X32 FILLER_177_2128 ();
 FILLCELL_X32 FILLER_177_2160 ();
 FILLCELL_X32 FILLER_177_2192 ();
 FILLCELL_X32 FILLER_177_2224 ();
 FILLCELL_X32 FILLER_177_2256 ();
 FILLCELL_X32 FILLER_177_2288 ();
 FILLCELL_X32 FILLER_177_2320 ();
 FILLCELL_X32 FILLER_177_2352 ();
 FILLCELL_X32 FILLER_177_2384 ();
 FILLCELL_X16 FILLER_177_2416 ();
 FILLCELL_X4 FILLER_177_2432 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X32 FILLER_178_1592 ();
 FILLCELL_X32 FILLER_178_1624 ();
 FILLCELL_X32 FILLER_178_1656 ();
 FILLCELL_X32 FILLER_178_1688 ();
 FILLCELL_X32 FILLER_178_1720 ();
 FILLCELL_X32 FILLER_178_1752 ();
 FILLCELL_X32 FILLER_178_1784 ();
 FILLCELL_X32 FILLER_178_1816 ();
 FILLCELL_X32 FILLER_178_1848 ();
 FILLCELL_X8 FILLER_178_1880 ();
 FILLCELL_X4 FILLER_178_1888 ();
 FILLCELL_X2 FILLER_178_1892 ();
 FILLCELL_X32 FILLER_178_1895 ();
 FILLCELL_X32 FILLER_178_1927 ();
 FILLCELL_X32 FILLER_178_1959 ();
 FILLCELL_X32 FILLER_178_1991 ();
 FILLCELL_X32 FILLER_178_2023 ();
 FILLCELL_X32 FILLER_178_2055 ();
 FILLCELL_X32 FILLER_178_2087 ();
 FILLCELL_X32 FILLER_178_2119 ();
 FILLCELL_X32 FILLER_178_2151 ();
 FILLCELL_X32 FILLER_178_2183 ();
 FILLCELL_X32 FILLER_178_2215 ();
 FILLCELL_X32 FILLER_178_2247 ();
 FILLCELL_X32 FILLER_178_2279 ();
 FILLCELL_X32 FILLER_178_2311 ();
 FILLCELL_X32 FILLER_178_2343 ();
 FILLCELL_X32 FILLER_178_2375 ();
 FILLCELL_X16 FILLER_178_2407 ();
 FILLCELL_X8 FILLER_178_2423 ();
 FILLCELL_X4 FILLER_178_2431 ();
 FILLCELL_X1 FILLER_178_2435 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X32 FILLER_179_1648 ();
 FILLCELL_X32 FILLER_179_1680 ();
 FILLCELL_X32 FILLER_179_1712 ();
 FILLCELL_X32 FILLER_179_1744 ();
 FILLCELL_X32 FILLER_179_1776 ();
 FILLCELL_X32 FILLER_179_1808 ();
 FILLCELL_X32 FILLER_179_1840 ();
 FILLCELL_X32 FILLER_179_1872 ();
 FILLCELL_X32 FILLER_179_1904 ();
 FILLCELL_X32 FILLER_179_1936 ();
 FILLCELL_X32 FILLER_179_1968 ();
 FILLCELL_X32 FILLER_179_2000 ();
 FILLCELL_X32 FILLER_179_2032 ();
 FILLCELL_X32 FILLER_179_2064 ();
 FILLCELL_X32 FILLER_179_2096 ();
 FILLCELL_X32 FILLER_179_2128 ();
 FILLCELL_X32 FILLER_179_2160 ();
 FILLCELL_X32 FILLER_179_2192 ();
 FILLCELL_X32 FILLER_179_2224 ();
 FILLCELL_X32 FILLER_179_2256 ();
 FILLCELL_X32 FILLER_179_2288 ();
 FILLCELL_X32 FILLER_179_2320 ();
 FILLCELL_X32 FILLER_179_2352 ();
 FILLCELL_X32 FILLER_179_2384 ();
 FILLCELL_X16 FILLER_179_2416 ();
 FILLCELL_X4 FILLER_179_2432 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X32 FILLER_180_1592 ();
 FILLCELL_X32 FILLER_180_1624 ();
 FILLCELL_X32 FILLER_180_1656 ();
 FILLCELL_X32 FILLER_180_1688 ();
 FILLCELL_X32 FILLER_180_1720 ();
 FILLCELL_X32 FILLER_180_1752 ();
 FILLCELL_X32 FILLER_180_1784 ();
 FILLCELL_X32 FILLER_180_1816 ();
 FILLCELL_X32 FILLER_180_1848 ();
 FILLCELL_X8 FILLER_180_1880 ();
 FILLCELL_X4 FILLER_180_1888 ();
 FILLCELL_X2 FILLER_180_1892 ();
 FILLCELL_X32 FILLER_180_1895 ();
 FILLCELL_X32 FILLER_180_1927 ();
 FILLCELL_X32 FILLER_180_1959 ();
 FILLCELL_X32 FILLER_180_1991 ();
 FILLCELL_X32 FILLER_180_2023 ();
 FILLCELL_X32 FILLER_180_2055 ();
 FILLCELL_X32 FILLER_180_2087 ();
 FILLCELL_X32 FILLER_180_2119 ();
 FILLCELL_X32 FILLER_180_2151 ();
 FILLCELL_X32 FILLER_180_2183 ();
 FILLCELL_X32 FILLER_180_2215 ();
 FILLCELL_X32 FILLER_180_2247 ();
 FILLCELL_X32 FILLER_180_2279 ();
 FILLCELL_X32 FILLER_180_2311 ();
 FILLCELL_X32 FILLER_180_2343 ();
 FILLCELL_X32 FILLER_180_2375 ();
 FILLCELL_X16 FILLER_180_2407 ();
 FILLCELL_X8 FILLER_180_2423 ();
 FILLCELL_X4 FILLER_180_2431 ();
 FILLCELL_X1 FILLER_180_2435 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X32 FILLER_181_1648 ();
 FILLCELL_X32 FILLER_181_1680 ();
 FILLCELL_X32 FILLER_181_1712 ();
 FILLCELL_X32 FILLER_181_1744 ();
 FILLCELL_X32 FILLER_181_1776 ();
 FILLCELL_X32 FILLER_181_1808 ();
 FILLCELL_X32 FILLER_181_1840 ();
 FILLCELL_X32 FILLER_181_1872 ();
 FILLCELL_X32 FILLER_181_1904 ();
 FILLCELL_X32 FILLER_181_1936 ();
 FILLCELL_X32 FILLER_181_1968 ();
 FILLCELL_X32 FILLER_181_2000 ();
 FILLCELL_X32 FILLER_181_2032 ();
 FILLCELL_X32 FILLER_181_2064 ();
 FILLCELL_X32 FILLER_181_2096 ();
 FILLCELL_X32 FILLER_181_2128 ();
 FILLCELL_X32 FILLER_181_2160 ();
 FILLCELL_X32 FILLER_181_2192 ();
 FILLCELL_X32 FILLER_181_2224 ();
 FILLCELL_X32 FILLER_181_2256 ();
 FILLCELL_X32 FILLER_181_2288 ();
 FILLCELL_X32 FILLER_181_2320 ();
 FILLCELL_X32 FILLER_181_2352 ();
 FILLCELL_X32 FILLER_181_2384 ();
 FILLCELL_X16 FILLER_181_2416 ();
 FILLCELL_X4 FILLER_181_2432 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X32 FILLER_182_1592 ();
 FILLCELL_X32 FILLER_182_1624 ();
 FILLCELL_X32 FILLER_182_1656 ();
 FILLCELL_X32 FILLER_182_1688 ();
 FILLCELL_X32 FILLER_182_1720 ();
 FILLCELL_X32 FILLER_182_1752 ();
 FILLCELL_X32 FILLER_182_1784 ();
 FILLCELL_X32 FILLER_182_1816 ();
 FILLCELL_X32 FILLER_182_1848 ();
 FILLCELL_X8 FILLER_182_1880 ();
 FILLCELL_X4 FILLER_182_1888 ();
 FILLCELL_X2 FILLER_182_1892 ();
 FILLCELL_X32 FILLER_182_1895 ();
 FILLCELL_X32 FILLER_182_1927 ();
 FILLCELL_X32 FILLER_182_1959 ();
 FILLCELL_X32 FILLER_182_1991 ();
 FILLCELL_X32 FILLER_182_2023 ();
 FILLCELL_X32 FILLER_182_2055 ();
 FILLCELL_X32 FILLER_182_2087 ();
 FILLCELL_X32 FILLER_182_2119 ();
 FILLCELL_X32 FILLER_182_2151 ();
 FILLCELL_X32 FILLER_182_2183 ();
 FILLCELL_X32 FILLER_182_2215 ();
 FILLCELL_X32 FILLER_182_2247 ();
 FILLCELL_X32 FILLER_182_2279 ();
 FILLCELL_X32 FILLER_182_2311 ();
 FILLCELL_X32 FILLER_182_2343 ();
 FILLCELL_X32 FILLER_182_2375 ();
 FILLCELL_X16 FILLER_182_2407 ();
 FILLCELL_X8 FILLER_182_2423 ();
 FILLCELL_X4 FILLER_182_2431 ();
 FILLCELL_X1 FILLER_182_2435 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X32 FILLER_183_1648 ();
 FILLCELL_X32 FILLER_183_1680 ();
 FILLCELL_X32 FILLER_183_1712 ();
 FILLCELL_X32 FILLER_183_1744 ();
 FILLCELL_X32 FILLER_183_1776 ();
 FILLCELL_X32 FILLER_183_1808 ();
 FILLCELL_X32 FILLER_183_1840 ();
 FILLCELL_X32 FILLER_183_1872 ();
 FILLCELL_X32 FILLER_183_1904 ();
 FILLCELL_X32 FILLER_183_1936 ();
 FILLCELL_X32 FILLER_183_1968 ();
 FILLCELL_X32 FILLER_183_2000 ();
 FILLCELL_X32 FILLER_183_2032 ();
 FILLCELL_X32 FILLER_183_2064 ();
 FILLCELL_X32 FILLER_183_2096 ();
 FILLCELL_X32 FILLER_183_2128 ();
 FILLCELL_X32 FILLER_183_2160 ();
 FILLCELL_X32 FILLER_183_2192 ();
 FILLCELL_X32 FILLER_183_2224 ();
 FILLCELL_X32 FILLER_183_2256 ();
 FILLCELL_X32 FILLER_183_2288 ();
 FILLCELL_X32 FILLER_183_2320 ();
 FILLCELL_X32 FILLER_183_2352 ();
 FILLCELL_X32 FILLER_183_2384 ();
 FILLCELL_X16 FILLER_183_2416 ();
 FILLCELL_X4 FILLER_183_2432 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X32 FILLER_184_1592 ();
 FILLCELL_X32 FILLER_184_1624 ();
 FILLCELL_X32 FILLER_184_1656 ();
 FILLCELL_X32 FILLER_184_1688 ();
 FILLCELL_X32 FILLER_184_1720 ();
 FILLCELL_X32 FILLER_184_1752 ();
 FILLCELL_X32 FILLER_184_1784 ();
 FILLCELL_X32 FILLER_184_1816 ();
 FILLCELL_X32 FILLER_184_1848 ();
 FILLCELL_X8 FILLER_184_1880 ();
 FILLCELL_X4 FILLER_184_1888 ();
 FILLCELL_X2 FILLER_184_1892 ();
 FILLCELL_X32 FILLER_184_1895 ();
 FILLCELL_X32 FILLER_184_1927 ();
 FILLCELL_X32 FILLER_184_1959 ();
 FILLCELL_X32 FILLER_184_1991 ();
 FILLCELL_X32 FILLER_184_2023 ();
 FILLCELL_X32 FILLER_184_2055 ();
 FILLCELL_X32 FILLER_184_2087 ();
 FILLCELL_X32 FILLER_184_2119 ();
 FILLCELL_X32 FILLER_184_2151 ();
 FILLCELL_X32 FILLER_184_2183 ();
 FILLCELL_X32 FILLER_184_2215 ();
 FILLCELL_X32 FILLER_184_2247 ();
 FILLCELL_X32 FILLER_184_2279 ();
 FILLCELL_X32 FILLER_184_2311 ();
 FILLCELL_X32 FILLER_184_2343 ();
 FILLCELL_X32 FILLER_184_2375 ();
 FILLCELL_X16 FILLER_184_2407 ();
 FILLCELL_X8 FILLER_184_2423 ();
 FILLCELL_X4 FILLER_184_2431 ();
 FILLCELL_X1 FILLER_184_2435 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X32 FILLER_185_1776 ();
 FILLCELL_X32 FILLER_185_1808 ();
 FILLCELL_X32 FILLER_185_1840 ();
 FILLCELL_X32 FILLER_185_1872 ();
 FILLCELL_X32 FILLER_185_1904 ();
 FILLCELL_X32 FILLER_185_1936 ();
 FILLCELL_X32 FILLER_185_1968 ();
 FILLCELL_X32 FILLER_185_2000 ();
 FILLCELL_X32 FILLER_185_2032 ();
 FILLCELL_X32 FILLER_185_2064 ();
 FILLCELL_X32 FILLER_185_2096 ();
 FILLCELL_X32 FILLER_185_2128 ();
 FILLCELL_X32 FILLER_185_2160 ();
 FILLCELL_X32 FILLER_185_2192 ();
 FILLCELL_X32 FILLER_185_2224 ();
 FILLCELL_X32 FILLER_185_2256 ();
 FILLCELL_X32 FILLER_185_2288 ();
 FILLCELL_X32 FILLER_185_2320 ();
 FILLCELL_X32 FILLER_185_2352 ();
 FILLCELL_X32 FILLER_185_2384 ();
 FILLCELL_X16 FILLER_185_2416 ();
 FILLCELL_X4 FILLER_185_2432 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X32 FILLER_186_1592 ();
 FILLCELL_X32 FILLER_186_1624 ();
 FILLCELL_X32 FILLER_186_1656 ();
 FILLCELL_X32 FILLER_186_1688 ();
 FILLCELL_X32 FILLER_186_1720 ();
 FILLCELL_X32 FILLER_186_1752 ();
 FILLCELL_X32 FILLER_186_1784 ();
 FILLCELL_X32 FILLER_186_1816 ();
 FILLCELL_X32 FILLER_186_1848 ();
 FILLCELL_X8 FILLER_186_1880 ();
 FILLCELL_X4 FILLER_186_1888 ();
 FILLCELL_X2 FILLER_186_1892 ();
 FILLCELL_X32 FILLER_186_1895 ();
 FILLCELL_X32 FILLER_186_1927 ();
 FILLCELL_X32 FILLER_186_1959 ();
 FILLCELL_X32 FILLER_186_1991 ();
 FILLCELL_X32 FILLER_186_2023 ();
 FILLCELL_X32 FILLER_186_2055 ();
 FILLCELL_X32 FILLER_186_2087 ();
 FILLCELL_X32 FILLER_186_2119 ();
 FILLCELL_X32 FILLER_186_2151 ();
 FILLCELL_X32 FILLER_186_2183 ();
 FILLCELL_X32 FILLER_186_2215 ();
 FILLCELL_X32 FILLER_186_2247 ();
 FILLCELL_X32 FILLER_186_2279 ();
 FILLCELL_X32 FILLER_186_2311 ();
 FILLCELL_X32 FILLER_186_2343 ();
 FILLCELL_X32 FILLER_186_2375 ();
 FILLCELL_X16 FILLER_186_2407 ();
 FILLCELL_X8 FILLER_186_2423 ();
 FILLCELL_X4 FILLER_186_2431 ();
 FILLCELL_X1 FILLER_186_2435 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X32 FILLER_187_1648 ();
 FILLCELL_X32 FILLER_187_1680 ();
 FILLCELL_X32 FILLER_187_1712 ();
 FILLCELL_X32 FILLER_187_1744 ();
 FILLCELL_X32 FILLER_187_1776 ();
 FILLCELL_X32 FILLER_187_1808 ();
 FILLCELL_X32 FILLER_187_1840 ();
 FILLCELL_X32 FILLER_187_1872 ();
 FILLCELL_X32 FILLER_187_1904 ();
 FILLCELL_X32 FILLER_187_1936 ();
 FILLCELL_X32 FILLER_187_1968 ();
 FILLCELL_X32 FILLER_187_2000 ();
 FILLCELL_X32 FILLER_187_2032 ();
 FILLCELL_X32 FILLER_187_2064 ();
 FILLCELL_X32 FILLER_187_2096 ();
 FILLCELL_X32 FILLER_187_2128 ();
 FILLCELL_X32 FILLER_187_2160 ();
 FILLCELL_X32 FILLER_187_2192 ();
 FILLCELL_X32 FILLER_187_2224 ();
 FILLCELL_X32 FILLER_187_2256 ();
 FILLCELL_X32 FILLER_187_2288 ();
 FILLCELL_X32 FILLER_187_2320 ();
 FILLCELL_X32 FILLER_187_2352 ();
 FILLCELL_X32 FILLER_187_2384 ();
 FILLCELL_X16 FILLER_187_2416 ();
 FILLCELL_X4 FILLER_187_2432 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X32 FILLER_188_1592 ();
 FILLCELL_X32 FILLER_188_1624 ();
 FILLCELL_X32 FILLER_188_1656 ();
 FILLCELL_X32 FILLER_188_1688 ();
 FILLCELL_X32 FILLER_188_1720 ();
 FILLCELL_X32 FILLER_188_1752 ();
 FILLCELL_X32 FILLER_188_1784 ();
 FILLCELL_X32 FILLER_188_1816 ();
 FILLCELL_X32 FILLER_188_1848 ();
 FILLCELL_X8 FILLER_188_1880 ();
 FILLCELL_X4 FILLER_188_1888 ();
 FILLCELL_X2 FILLER_188_1892 ();
 FILLCELL_X32 FILLER_188_1895 ();
 FILLCELL_X32 FILLER_188_1927 ();
 FILLCELL_X32 FILLER_188_1959 ();
 FILLCELL_X32 FILLER_188_1991 ();
 FILLCELL_X32 FILLER_188_2023 ();
 FILLCELL_X32 FILLER_188_2055 ();
 FILLCELL_X32 FILLER_188_2087 ();
 FILLCELL_X32 FILLER_188_2119 ();
 FILLCELL_X32 FILLER_188_2151 ();
 FILLCELL_X32 FILLER_188_2183 ();
 FILLCELL_X32 FILLER_188_2215 ();
 FILLCELL_X32 FILLER_188_2247 ();
 FILLCELL_X32 FILLER_188_2279 ();
 FILLCELL_X32 FILLER_188_2311 ();
 FILLCELL_X32 FILLER_188_2343 ();
 FILLCELL_X32 FILLER_188_2375 ();
 FILLCELL_X1 FILLER_188_2407 ();
 FILLCELL_X16 FILLER_188_2411 ();
 FILLCELL_X8 FILLER_188_2427 ();
 FILLCELL_X1 FILLER_188_2435 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X32 FILLER_189_1648 ();
 FILLCELL_X32 FILLER_189_1680 ();
 FILLCELL_X32 FILLER_189_1712 ();
 FILLCELL_X32 FILLER_189_1744 ();
 FILLCELL_X32 FILLER_189_1776 ();
 FILLCELL_X32 FILLER_189_1808 ();
 FILLCELL_X32 FILLER_189_1840 ();
 FILLCELL_X32 FILLER_189_1872 ();
 FILLCELL_X32 FILLER_189_1904 ();
 FILLCELL_X32 FILLER_189_1936 ();
 FILLCELL_X32 FILLER_189_1968 ();
 FILLCELL_X32 FILLER_189_2000 ();
 FILLCELL_X32 FILLER_189_2032 ();
 FILLCELL_X32 FILLER_189_2064 ();
 FILLCELL_X32 FILLER_189_2096 ();
 FILLCELL_X32 FILLER_189_2128 ();
 FILLCELL_X32 FILLER_189_2160 ();
 FILLCELL_X32 FILLER_189_2192 ();
 FILLCELL_X32 FILLER_189_2224 ();
 FILLCELL_X32 FILLER_189_2256 ();
 FILLCELL_X32 FILLER_189_2288 ();
 FILLCELL_X32 FILLER_189_2320 ();
 FILLCELL_X32 FILLER_189_2352 ();
 FILLCELL_X32 FILLER_189_2384 ();
 FILLCELL_X16 FILLER_189_2416 ();
 FILLCELL_X4 FILLER_189_2432 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X32 FILLER_190_1592 ();
 FILLCELL_X32 FILLER_190_1624 ();
 FILLCELL_X32 FILLER_190_1656 ();
 FILLCELL_X32 FILLER_190_1688 ();
 FILLCELL_X32 FILLER_190_1720 ();
 FILLCELL_X32 FILLER_190_1752 ();
 FILLCELL_X32 FILLER_190_1784 ();
 FILLCELL_X32 FILLER_190_1816 ();
 FILLCELL_X32 FILLER_190_1848 ();
 FILLCELL_X8 FILLER_190_1880 ();
 FILLCELL_X4 FILLER_190_1888 ();
 FILLCELL_X2 FILLER_190_1892 ();
 FILLCELL_X32 FILLER_190_1895 ();
 FILLCELL_X32 FILLER_190_1927 ();
 FILLCELL_X32 FILLER_190_1959 ();
 FILLCELL_X32 FILLER_190_1991 ();
 FILLCELL_X32 FILLER_190_2023 ();
 FILLCELL_X32 FILLER_190_2055 ();
 FILLCELL_X32 FILLER_190_2087 ();
 FILLCELL_X32 FILLER_190_2119 ();
 FILLCELL_X32 FILLER_190_2151 ();
 FILLCELL_X32 FILLER_190_2183 ();
 FILLCELL_X32 FILLER_190_2215 ();
 FILLCELL_X32 FILLER_190_2247 ();
 FILLCELL_X32 FILLER_190_2279 ();
 FILLCELL_X32 FILLER_190_2311 ();
 FILLCELL_X32 FILLER_190_2343 ();
 FILLCELL_X32 FILLER_190_2375 ();
 FILLCELL_X16 FILLER_190_2407 ();
 FILLCELL_X8 FILLER_190_2423 ();
 FILLCELL_X4 FILLER_190_2431 ();
 FILLCELL_X1 FILLER_190_2435 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X32 FILLER_191_1648 ();
 FILLCELL_X32 FILLER_191_1680 ();
 FILLCELL_X32 FILLER_191_1712 ();
 FILLCELL_X32 FILLER_191_1744 ();
 FILLCELL_X32 FILLER_191_1776 ();
 FILLCELL_X32 FILLER_191_1808 ();
 FILLCELL_X32 FILLER_191_1840 ();
 FILLCELL_X32 FILLER_191_1872 ();
 FILLCELL_X32 FILLER_191_1904 ();
 FILLCELL_X32 FILLER_191_1936 ();
 FILLCELL_X32 FILLER_191_1968 ();
 FILLCELL_X32 FILLER_191_2000 ();
 FILLCELL_X32 FILLER_191_2032 ();
 FILLCELL_X32 FILLER_191_2064 ();
 FILLCELL_X32 FILLER_191_2096 ();
 FILLCELL_X32 FILLER_191_2128 ();
 FILLCELL_X32 FILLER_191_2160 ();
 FILLCELL_X32 FILLER_191_2192 ();
 FILLCELL_X32 FILLER_191_2224 ();
 FILLCELL_X32 FILLER_191_2256 ();
 FILLCELL_X32 FILLER_191_2288 ();
 FILLCELL_X32 FILLER_191_2320 ();
 FILLCELL_X32 FILLER_191_2352 ();
 FILLCELL_X32 FILLER_191_2384 ();
 FILLCELL_X16 FILLER_191_2416 ();
 FILLCELL_X4 FILLER_191_2432 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X32 FILLER_192_1592 ();
 FILLCELL_X32 FILLER_192_1624 ();
 FILLCELL_X32 FILLER_192_1656 ();
 FILLCELL_X32 FILLER_192_1688 ();
 FILLCELL_X32 FILLER_192_1720 ();
 FILLCELL_X32 FILLER_192_1752 ();
 FILLCELL_X32 FILLER_192_1784 ();
 FILLCELL_X32 FILLER_192_1816 ();
 FILLCELL_X32 FILLER_192_1848 ();
 FILLCELL_X8 FILLER_192_1880 ();
 FILLCELL_X4 FILLER_192_1888 ();
 FILLCELL_X2 FILLER_192_1892 ();
 FILLCELL_X32 FILLER_192_1895 ();
 FILLCELL_X32 FILLER_192_1927 ();
 FILLCELL_X32 FILLER_192_1959 ();
 FILLCELL_X32 FILLER_192_1991 ();
 FILLCELL_X32 FILLER_192_2023 ();
 FILLCELL_X32 FILLER_192_2055 ();
 FILLCELL_X32 FILLER_192_2087 ();
 FILLCELL_X32 FILLER_192_2119 ();
 FILLCELL_X32 FILLER_192_2151 ();
 FILLCELL_X32 FILLER_192_2183 ();
 FILLCELL_X32 FILLER_192_2215 ();
 FILLCELL_X32 FILLER_192_2247 ();
 FILLCELL_X32 FILLER_192_2279 ();
 FILLCELL_X32 FILLER_192_2311 ();
 FILLCELL_X32 FILLER_192_2343 ();
 FILLCELL_X32 FILLER_192_2375 ();
 FILLCELL_X16 FILLER_192_2407 ();
 FILLCELL_X8 FILLER_192_2423 ();
 FILLCELL_X4 FILLER_192_2431 ();
 FILLCELL_X1 FILLER_192_2435 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X32 FILLER_193_1648 ();
 FILLCELL_X32 FILLER_193_1680 ();
 FILLCELL_X32 FILLER_193_1712 ();
 FILLCELL_X32 FILLER_193_1744 ();
 FILLCELL_X32 FILLER_193_1776 ();
 FILLCELL_X32 FILLER_193_1808 ();
 FILLCELL_X32 FILLER_193_1840 ();
 FILLCELL_X32 FILLER_193_1872 ();
 FILLCELL_X32 FILLER_193_1904 ();
 FILLCELL_X32 FILLER_193_1936 ();
 FILLCELL_X32 FILLER_193_1968 ();
 FILLCELL_X32 FILLER_193_2000 ();
 FILLCELL_X32 FILLER_193_2032 ();
 FILLCELL_X32 FILLER_193_2064 ();
 FILLCELL_X32 FILLER_193_2096 ();
 FILLCELL_X32 FILLER_193_2128 ();
 FILLCELL_X32 FILLER_193_2160 ();
 FILLCELL_X32 FILLER_193_2192 ();
 FILLCELL_X32 FILLER_193_2224 ();
 FILLCELL_X32 FILLER_193_2256 ();
 FILLCELL_X32 FILLER_193_2288 ();
 FILLCELL_X32 FILLER_193_2320 ();
 FILLCELL_X32 FILLER_193_2352 ();
 FILLCELL_X32 FILLER_193_2384 ();
 FILLCELL_X16 FILLER_193_2416 ();
 FILLCELL_X4 FILLER_193_2432 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X32 FILLER_194_1592 ();
 FILLCELL_X32 FILLER_194_1624 ();
 FILLCELL_X32 FILLER_194_1656 ();
 FILLCELL_X32 FILLER_194_1688 ();
 FILLCELL_X32 FILLER_194_1720 ();
 FILLCELL_X32 FILLER_194_1752 ();
 FILLCELL_X32 FILLER_194_1784 ();
 FILLCELL_X32 FILLER_194_1816 ();
 FILLCELL_X32 FILLER_194_1848 ();
 FILLCELL_X8 FILLER_194_1880 ();
 FILLCELL_X4 FILLER_194_1888 ();
 FILLCELL_X2 FILLER_194_1892 ();
 FILLCELL_X32 FILLER_194_1895 ();
 FILLCELL_X32 FILLER_194_1927 ();
 FILLCELL_X32 FILLER_194_1959 ();
 FILLCELL_X32 FILLER_194_1991 ();
 FILLCELL_X32 FILLER_194_2023 ();
 FILLCELL_X32 FILLER_194_2055 ();
 FILLCELL_X32 FILLER_194_2087 ();
 FILLCELL_X32 FILLER_194_2119 ();
 FILLCELL_X32 FILLER_194_2151 ();
 FILLCELL_X32 FILLER_194_2183 ();
 FILLCELL_X32 FILLER_194_2215 ();
 FILLCELL_X32 FILLER_194_2247 ();
 FILLCELL_X32 FILLER_194_2279 ();
 FILLCELL_X32 FILLER_194_2311 ();
 FILLCELL_X32 FILLER_194_2343 ();
 FILLCELL_X32 FILLER_194_2375 ();
 FILLCELL_X16 FILLER_194_2407 ();
 FILLCELL_X8 FILLER_194_2423 ();
 FILLCELL_X4 FILLER_194_2431 ();
 FILLCELL_X1 FILLER_194_2435 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X32 FILLER_195_1648 ();
 FILLCELL_X32 FILLER_195_1680 ();
 FILLCELL_X32 FILLER_195_1712 ();
 FILLCELL_X32 FILLER_195_1744 ();
 FILLCELL_X32 FILLER_195_1776 ();
 FILLCELL_X32 FILLER_195_1808 ();
 FILLCELL_X32 FILLER_195_1840 ();
 FILLCELL_X32 FILLER_195_1872 ();
 FILLCELL_X32 FILLER_195_1904 ();
 FILLCELL_X32 FILLER_195_1936 ();
 FILLCELL_X32 FILLER_195_1968 ();
 FILLCELL_X32 FILLER_195_2000 ();
 FILLCELL_X32 FILLER_195_2032 ();
 FILLCELL_X32 FILLER_195_2064 ();
 FILLCELL_X32 FILLER_195_2096 ();
 FILLCELL_X32 FILLER_195_2128 ();
 FILLCELL_X32 FILLER_195_2160 ();
 FILLCELL_X32 FILLER_195_2192 ();
 FILLCELL_X32 FILLER_195_2224 ();
 FILLCELL_X32 FILLER_195_2256 ();
 FILLCELL_X32 FILLER_195_2288 ();
 FILLCELL_X32 FILLER_195_2320 ();
 FILLCELL_X32 FILLER_195_2352 ();
 FILLCELL_X32 FILLER_195_2384 ();
 FILLCELL_X16 FILLER_195_2416 ();
 FILLCELL_X4 FILLER_195_2432 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X32 FILLER_196_1592 ();
 FILLCELL_X32 FILLER_196_1624 ();
 FILLCELL_X32 FILLER_196_1656 ();
 FILLCELL_X32 FILLER_196_1688 ();
 FILLCELL_X32 FILLER_196_1720 ();
 FILLCELL_X32 FILLER_196_1752 ();
 FILLCELL_X32 FILLER_196_1784 ();
 FILLCELL_X32 FILLER_196_1816 ();
 FILLCELL_X32 FILLER_196_1848 ();
 FILLCELL_X8 FILLER_196_1880 ();
 FILLCELL_X4 FILLER_196_1888 ();
 FILLCELL_X2 FILLER_196_1892 ();
 FILLCELL_X32 FILLER_196_1895 ();
 FILLCELL_X32 FILLER_196_1927 ();
 FILLCELL_X32 FILLER_196_1959 ();
 FILLCELL_X32 FILLER_196_1991 ();
 FILLCELL_X32 FILLER_196_2023 ();
 FILLCELL_X32 FILLER_196_2055 ();
 FILLCELL_X32 FILLER_196_2087 ();
 FILLCELL_X32 FILLER_196_2119 ();
 FILLCELL_X32 FILLER_196_2151 ();
 FILLCELL_X32 FILLER_196_2183 ();
 FILLCELL_X32 FILLER_196_2215 ();
 FILLCELL_X32 FILLER_196_2247 ();
 FILLCELL_X32 FILLER_196_2279 ();
 FILLCELL_X32 FILLER_196_2311 ();
 FILLCELL_X32 FILLER_196_2343 ();
 FILLCELL_X32 FILLER_196_2375 ();
 FILLCELL_X16 FILLER_196_2407 ();
 FILLCELL_X8 FILLER_196_2423 ();
 FILLCELL_X4 FILLER_196_2431 ();
 FILLCELL_X1 FILLER_196_2435 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X32 FILLER_197_1648 ();
 FILLCELL_X32 FILLER_197_1680 ();
 FILLCELL_X32 FILLER_197_1712 ();
 FILLCELL_X32 FILLER_197_1744 ();
 FILLCELL_X32 FILLER_197_1776 ();
 FILLCELL_X32 FILLER_197_1808 ();
 FILLCELL_X32 FILLER_197_1840 ();
 FILLCELL_X32 FILLER_197_1872 ();
 FILLCELL_X32 FILLER_197_1904 ();
 FILLCELL_X32 FILLER_197_1936 ();
 FILLCELL_X32 FILLER_197_1968 ();
 FILLCELL_X32 FILLER_197_2000 ();
 FILLCELL_X32 FILLER_197_2032 ();
 FILLCELL_X32 FILLER_197_2064 ();
 FILLCELL_X32 FILLER_197_2096 ();
 FILLCELL_X32 FILLER_197_2128 ();
 FILLCELL_X32 FILLER_197_2160 ();
 FILLCELL_X32 FILLER_197_2192 ();
 FILLCELL_X32 FILLER_197_2224 ();
 FILLCELL_X32 FILLER_197_2256 ();
 FILLCELL_X32 FILLER_197_2288 ();
 FILLCELL_X32 FILLER_197_2320 ();
 FILLCELL_X32 FILLER_197_2352 ();
 FILLCELL_X32 FILLER_197_2384 ();
 FILLCELL_X16 FILLER_197_2416 ();
 FILLCELL_X4 FILLER_197_2432 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X32 FILLER_198_1592 ();
 FILLCELL_X32 FILLER_198_1624 ();
 FILLCELL_X32 FILLER_198_1656 ();
 FILLCELL_X32 FILLER_198_1688 ();
 FILLCELL_X32 FILLER_198_1720 ();
 FILLCELL_X32 FILLER_198_1752 ();
 FILLCELL_X32 FILLER_198_1784 ();
 FILLCELL_X32 FILLER_198_1816 ();
 FILLCELL_X32 FILLER_198_1848 ();
 FILLCELL_X8 FILLER_198_1880 ();
 FILLCELL_X4 FILLER_198_1888 ();
 FILLCELL_X2 FILLER_198_1892 ();
 FILLCELL_X32 FILLER_198_1895 ();
 FILLCELL_X32 FILLER_198_1927 ();
 FILLCELL_X32 FILLER_198_1959 ();
 FILLCELL_X32 FILLER_198_1991 ();
 FILLCELL_X32 FILLER_198_2023 ();
 FILLCELL_X32 FILLER_198_2055 ();
 FILLCELL_X32 FILLER_198_2087 ();
 FILLCELL_X32 FILLER_198_2119 ();
 FILLCELL_X32 FILLER_198_2151 ();
 FILLCELL_X32 FILLER_198_2183 ();
 FILLCELL_X32 FILLER_198_2215 ();
 FILLCELL_X32 FILLER_198_2247 ();
 FILLCELL_X32 FILLER_198_2279 ();
 FILLCELL_X32 FILLER_198_2311 ();
 FILLCELL_X32 FILLER_198_2343 ();
 FILLCELL_X32 FILLER_198_2375 ();
 FILLCELL_X16 FILLER_198_2407 ();
 FILLCELL_X8 FILLER_198_2423 ();
 FILLCELL_X4 FILLER_198_2431 ();
 FILLCELL_X1 FILLER_198_2435 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X32 FILLER_199_1648 ();
 FILLCELL_X32 FILLER_199_1680 ();
 FILLCELL_X32 FILLER_199_1712 ();
 FILLCELL_X32 FILLER_199_1744 ();
 FILLCELL_X32 FILLER_199_1776 ();
 FILLCELL_X32 FILLER_199_1808 ();
 FILLCELL_X32 FILLER_199_1840 ();
 FILLCELL_X32 FILLER_199_1872 ();
 FILLCELL_X32 FILLER_199_1904 ();
 FILLCELL_X32 FILLER_199_1936 ();
 FILLCELL_X32 FILLER_199_1968 ();
 FILLCELL_X32 FILLER_199_2000 ();
 FILLCELL_X32 FILLER_199_2032 ();
 FILLCELL_X32 FILLER_199_2064 ();
 FILLCELL_X32 FILLER_199_2096 ();
 FILLCELL_X32 FILLER_199_2128 ();
 FILLCELL_X32 FILLER_199_2160 ();
 FILLCELL_X32 FILLER_199_2192 ();
 FILLCELL_X32 FILLER_199_2224 ();
 FILLCELL_X32 FILLER_199_2256 ();
 FILLCELL_X32 FILLER_199_2288 ();
 FILLCELL_X32 FILLER_199_2320 ();
 FILLCELL_X32 FILLER_199_2352 ();
 FILLCELL_X32 FILLER_199_2384 ();
 FILLCELL_X16 FILLER_199_2416 ();
 FILLCELL_X4 FILLER_199_2432 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X32 FILLER_200_1592 ();
 FILLCELL_X32 FILLER_200_1624 ();
 FILLCELL_X32 FILLER_200_1656 ();
 FILLCELL_X32 FILLER_200_1688 ();
 FILLCELL_X32 FILLER_200_1720 ();
 FILLCELL_X32 FILLER_200_1752 ();
 FILLCELL_X32 FILLER_200_1784 ();
 FILLCELL_X32 FILLER_200_1816 ();
 FILLCELL_X32 FILLER_200_1848 ();
 FILLCELL_X8 FILLER_200_1880 ();
 FILLCELL_X4 FILLER_200_1888 ();
 FILLCELL_X2 FILLER_200_1892 ();
 FILLCELL_X32 FILLER_200_1895 ();
 FILLCELL_X32 FILLER_200_1927 ();
 FILLCELL_X32 FILLER_200_1959 ();
 FILLCELL_X32 FILLER_200_1991 ();
 FILLCELL_X32 FILLER_200_2023 ();
 FILLCELL_X32 FILLER_200_2055 ();
 FILLCELL_X32 FILLER_200_2087 ();
 FILLCELL_X32 FILLER_200_2119 ();
 FILLCELL_X32 FILLER_200_2151 ();
 FILLCELL_X32 FILLER_200_2183 ();
 FILLCELL_X32 FILLER_200_2215 ();
 FILLCELL_X32 FILLER_200_2247 ();
 FILLCELL_X32 FILLER_200_2279 ();
 FILLCELL_X32 FILLER_200_2311 ();
 FILLCELL_X32 FILLER_200_2343 ();
 FILLCELL_X32 FILLER_200_2375 ();
 FILLCELL_X16 FILLER_200_2407 ();
 FILLCELL_X8 FILLER_200_2423 ();
 FILLCELL_X4 FILLER_200_2431 ();
 FILLCELL_X1 FILLER_200_2435 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X32 FILLER_201_1776 ();
 FILLCELL_X32 FILLER_201_1808 ();
 FILLCELL_X32 FILLER_201_1840 ();
 FILLCELL_X32 FILLER_201_1872 ();
 FILLCELL_X32 FILLER_201_1904 ();
 FILLCELL_X32 FILLER_201_1936 ();
 FILLCELL_X32 FILLER_201_1968 ();
 FILLCELL_X32 FILLER_201_2000 ();
 FILLCELL_X32 FILLER_201_2032 ();
 FILLCELL_X32 FILLER_201_2064 ();
 FILLCELL_X32 FILLER_201_2096 ();
 FILLCELL_X32 FILLER_201_2128 ();
 FILLCELL_X32 FILLER_201_2160 ();
 FILLCELL_X32 FILLER_201_2192 ();
 FILLCELL_X32 FILLER_201_2224 ();
 FILLCELL_X32 FILLER_201_2256 ();
 FILLCELL_X32 FILLER_201_2288 ();
 FILLCELL_X32 FILLER_201_2320 ();
 FILLCELL_X32 FILLER_201_2352 ();
 FILLCELL_X32 FILLER_201_2384 ();
 FILLCELL_X16 FILLER_201_2416 ();
 FILLCELL_X4 FILLER_201_2432 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_202_1784 ();
 FILLCELL_X32 FILLER_202_1816 ();
 FILLCELL_X32 FILLER_202_1848 ();
 FILLCELL_X8 FILLER_202_1880 ();
 FILLCELL_X4 FILLER_202_1888 ();
 FILLCELL_X2 FILLER_202_1892 ();
 FILLCELL_X32 FILLER_202_1895 ();
 FILLCELL_X32 FILLER_202_1927 ();
 FILLCELL_X32 FILLER_202_1959 ();
 FILLCELL_X32 FILLER_202_1991 ();
 FILLCELL_X32 FILLER_202_2023 ();
 FILLCELL_X32 FILLER_202_2055 ();
 FILLCELL_X32 FILLER_202_2087 ();
 FILLCELL_X32 FILLER_202_2119 ();
 FILLCELL_X32 FILLER_202_2151 ();
 FILLCELL_X32 FILLER_202_2183 ();
 FILLCELL_X32 FILLER_202_2215 ();
 FILLCELL_X32 FILLER_202_2247 ();
 FILLCELL_X32 FILLER_202_2279 ();
 FILLCELL_X32 FILLER_202_2311 ();
 FILLCELL_X32 FILLER_202_2343 ();
 FILLCELL_X32 FILLER_202_2375 ();
 FILLCELL_X16 FILLER_202_2407 ();
 FILLCELL_X8 FILLER_202_2423 ();
 FILLCELL_X4 FILLER_202_2431 ();
 FILLCELL_X1 FILLER_202_2435 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X32 FILLER_203_1776 ();
 FILLCELL_X32 FILLER_203_1808 ();
 FILLCELL_X32 FILLER_203_1840 ();
 FILLCELL_X32 FILLER_203_1872 ();
 FILLCELL_X32 FILLER_203_1904 ();
 FILLCELL_X32 FILLER_203_1936 ();
 FILLCELL_X32 FILLER_203_1968 ();
 FILLCELL_X32 FILLER_203_2000 ();
 FILLCELL_X32 FILLER_203_2032 ();
 FILLCELL_X32 FILLER_203_2064 ();
 FILLCELL_X32 FILLER_203_2096 ();
 FILLCELL_X32 FILLER_203_2128 ();
 FILLCELL_X32 FILLER_203_2160 ();
 FILLCELL_X32 FILLER_203_2192 ();
 FILLCELL_X32 FILLER_203_2224 ();
 FILLCELL_X32 FILLER_203_2256 ();
 FILLCELL_X32 FILLER_203_2288 ();
 FILLCELL_X32 FILLER_203_2320 ();
 FILLCELL_X32 FILLER_203_2352 ();
 FILLCELL_X32 FILLER_203_2384 ();
 FILLCELL_X16 FILLER_203_2416 ();
 FILLCELL_X4 FILLER_203_2432 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X32 FILLER_204_1784 ();
 FILLCELL_X32 FILLER_204_1816 ();
 FILLCELL_X32 FILLER_204_1848 ();
 FILLCELL_X8 FILLER_204_1880 ();
 FILLCELL_X4 FILLER_204_1888 ();
 FILLCELL_X2 FILLER_204_1892 ();
 FILLCELL_X32 FILLER_204_1895 ();
 FILLCELL_X32 FILLER_204_1927 ();
 FILLCELL_X32 FILLER_204_1959 ();
 FILLCELL_X32 FILLER_204_1991 ();
 FILLCELL_X32 FILLER_204_2023 ();
 FILLCELL_X32 FILLER_204_2055 ();
 FILLCELL_X32 FILLER_204_2087 ();
 FILLCELL_X32 FILLER_204_2119 ();
 FILLCELL_X32 FILLER_204_2151 ();
 FILLCELL_X32 FILLER_204_2183 ();
 FILLCELL_X32 FILLER_204_2215 ();
 FILLCELL_X32 FILLER_204_2247 ();
 FILLCELL_X32 FILLER_204_2279 ();
 FILLCELL_X32 FILLER_204_2311 ();
 FILLCELL_X32 FILLER_204_2343 ();
 FILLCELL_X32 FILLER_204_2375 ();
 FILLCELL_X16 FILLER_204_2407 ();
 FILLCELL_X8 FILLER_204_2423 ();
 FILLCELL_X4 FILLER_204_2431 ();
 FILLCELL_X1 FILLER_204_2435 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X32 FILLER_205_1776 ();
 FILLCELL_X32 FILLER_205_1808 ();
 FILLCELL_X32 FILLER_205_1840 ();
 FILLCELL_X32 FILLER_205_1872 ();
 FILLCELL_X32 FILLER_205_1904 ();
 FILLCELL_X32 FILLER_205_1936 ();
 FILLCELL_X32 FILLER_205_1968 ();
 FILLCELL_X32 FILLER_205_2000 ();
 FILLCELL_X32 FILLER_205_2032 ();
 FILLCELL_X32 FILLER_205_2064 ();
 FILLCELL_X32 FILLER_205_2096 ();
 FILLCELL_X32 FILLER_205_2128 ();
 FILLCELL_X32 FILLER_205_2160 ();
 FILLCELL_X32 FILLER_205_2192 ();
 FILLCELL_X32 FILLER_205_2224 ();
 FILLCELL_X32 FILLER_205_2256 ();
 FILLCELL_X32 FILLER_205_2288 ();
 FILLCELL_X32 FILLER_205_2320 ();
 FILLCELL_X32 FILLER_205_2352 ();
 FILLCELL_X32 FILLER_205_2384 ();
 FILLCELL_X16 FILLER_205_2416 ();
 FILLCELL_X4 FILLER_205_2432 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X32 FILLER_206_1784 ();
 FILLCELL_X32 FILLER_206_1816 ();
 FILLCELL_X32 FILLER_206_1848 ();
 FILLCELL_X8 FILLER_206_1880 ();
 FILLCELL_X4 FILLER_206_1888 ();
 FILLCELL_X2 FILLER_206_1892 ();
 FILLCELL_X32 FILLER_206_1895 ();
 FILLCELL_X32 FILLER_206_1927 ();
 FILLCELL_X32 FILLER_206_1959 ();
 FILLCELL_X32 FILLER_206_1991 ();
 FILLCELL_X32 FILLER_206_2023 ();
 FILLCELL_X32 FILLER_206_2055 ();
 FILLCELL_X32 FILLER_206_2087 ();
 FILLCELL_X32 FILLER_206_2119 ();
 FILLCELL_X32 FILLER_206_2151 ();
 FILLCELL_X32 FILLER_206_2183 ();
 FILLCELL_X32 FILLER_206_2215 ();
 FILLCELL_X32 FILLER_206_2247 ();
 FILLCELL_X32 FILLER_206_2279 ();
 FILLCELL_X32 FILLER_206_2311 ();
 FILLCELL_X32 FILLER_206_2343 ();
 FILLCELL_X32 FILLER_206_2375 ();
 FILLCELL_X16 FILLER_206_2407 ();
 FILLCELL_X8 FILLER_206_2423 ();
 FILLCELL_X4 FILLER_206_2431 ();
 FILLCELL_X1 FILLER_206_2435 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X32 FILLER_207_1776 ();
 FILLCELL_X32 FILLER_207_1808 ();
 FILLCELL_X32 FILLER_207_1840 ();
 FILLCELL_X32 FILLER_207_1872 ();
 FILLCELL_X32 FILLER_207_1904 ();
 FILLCELL_X32 FILLER_207_1936 ();
 FILLCELL_X32 FILLER_207_1968 ();
 FILLCELL_X32 FILLER_207_2000 ();
 FILLCELL_X32 FILLER_207_2032 ();
 FILLCELL_X32 FILLER_207_2064 ();
 FILLCELL_X32 FILLER_207_2096 ();
 FILLCELL_X32 FILLER_207_2128 ();
 FILLCELL_X32 FILLER_207_2160 ();
 FILLCELL_X32 FILLER_207_2192 ();
 FILLCELL_X32 FILLER_207_2224 ();
 FILLCELL_X32 FILLER_207_2256 ();
 FILLCELL_X32 FILLER_207_2288 ();
 FILLCELL_X32 FILLER_207_2320 ();
 FILLCELL_X32 FILLER_207_2352 ();
 FILLCELL_X32 FILLER_207_2384 ();
 FILLCELL_X16 FILLER_207_2416 ();
 FILLCELL_X4 FILLER_207_2432 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X32 FILLER_208_1784 ();
 FILLCELL_X32 FILLER_208_1816 ();
 FILLCELL_X32 FILLER_208_1848 ();
 FILLCELL_X8 FILLER_208_1880 ();
 FILLCELL_X4 FILLER_208_1888 ();
 FILLCELL_X2 FILLER_208_1892 ();
 FILLCELL_X32 FILLER_208_1895 ();
 FILLCELL_X32 FILLER_208_1927 ();
 FILLCELL_X32 FILLER_208_1959 ();
 FILLCELL_X32 FILLER_208_1991 ();
 FILLCELL_X32 FILLER_208_2023 ();
 FILLCELL_X32 FILLER_208_2055 ();
 FILLCELL_X32 FILLER_208_2087 ();
 FILLCELL_X32 FILLER_208_2119 ();
 FILLCELL_X32 FILLER_208_2151 ();
 FILLCELL_X32 FILLER_208_2183 ();
 FILLCELL_X32 FILLER_208_2215 ();
 FILLCELL_X32 FILLER_208_2247 ();
 FILLCELL_X32 FILLER_208_2279 ();
 FILLCELL_X32 FILLER_208_2311 ();
 FILLCELL_X32 FILLER_208_2343 ();
 FILLCELL_X32 FILLER_208_2375 ();
 FILLCELL_X16 FILLER_208_2407 ();
 FILLCELL_X8 FILLER_208_2423 ();
 FILLCELL_X4 FILLER_208_2431 ();
 FILLCELL_X1 FILLER_208_2435 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X32 FILLER_209_1776 ();
 FILLCELL_X32 FILLER_209_1808 ();
 FILLCELL_X32 FILLER_209_1840 ();
 FILLCELL_X32 FILLER_209_1872 ();
 FILLCELL_X32 FILLER_209_1904 ();
 FILLCELL_X32 FILLER_209_1936 ();
 FILLCELL_X32 FILLER_209_1968 ();
 FILLCELL_X32 FILLER_209_2000 ();
 FILLCELL_X32 FILLER_209_2032 ();
 FILLCELL_X32 FILLER_209_2064 ();
 FILLCELL_X32 FILLER_209_2096 ();
 FILLCELL_X32 FILLER_209_2128 ();
 FILLCELL_X32 FILLER_209_2160 ();
 FILLCELL_X32 FILLER_209_2192 ();
 FILLCELL_X32 FILLER_209_2224 ();
 FILLCELL_X32 FILLER_209_2256 ();
 FILLCELL_X32 FILLER_209_2288 ();
 FILLCELL_X32 FILLER_209_2320 ();
 FILLCELL_X32 FILLER_209_2352 ();
 FILLCELL_X32 FILLER_209_2384 ();
 FILLCELL_X16 FILLER_209_2416 ();
 FILLCELL_X4 FILLER_209_2432 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_210_1784 ();
 FILLCELL_X32 FILLER_210_1816 ();
 FILLCELL_X32 FILLER_210_1848 ();
 FILLCELL_X8 FILLER_210_1880 ();
 FILLCELL_X4 FILLER_210_1888 ();
 FILLCELL_X2 FILLER_210_1892 ();
 FILLCELL_X32 FILLER_210_1895 ();
 FILLCELL_X32 FILLER_210_1927 ();
 FILLCELL_X32 FILLER_210_1959 ();
 FILLCELL_X32 FILLER_210_1991 ();
 FILLCELL_X32 FILLER_210_2023 ();
 FILLCELL_X32 FILLER_210_2055 ();
 FILLCELL_X32 FILLER_210_2087 ();
 FILLCELL_X32 FILLER_210_2119 ();
 FILLCELL_X32 FILLER_210_2151 ();
 FILLCELL_X32 FILLER_210_2183 ();
 FILLCELL_X32 FILLER_210_2215 ();
 FILLCELL_X32 FILLER_210_2247 ();
 FILLCELL_X32 FILLER_210_2279 ();
 FILLCELL_X32 FILLER_210_2311 ();
 FILLCELL_X32 FILLER_210_2343 ();
 FILLCELL_X32 FILLER_210_2375 ();
 FILLCELL_X16 FILLER_210_2407 ();
 FILLCELL_X8 FILLER_210_2423 ();
 FILLCELL_X4 FILLER_210_2431 ();
 FILLCELL_X1 FILLER_210_2435 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X32 FILLER_211_1776 ();
 FILLCELL_X32 FILLER_211_1808 ();
 FILLCELL_X32 FILLER_211_1840 ();
 FILLCELL_X32 FILLER_211_1872 ();
 FILLCELL_X32 FILLER_211_1904 ();
 FILLCELL_X32 FILLER_211_1936 ();
 FILLCELL_X32 FILLER_211_1968 ();
 FILLCELL_X32 FILLER_211_2000 ();
 FILLCELL_X32 FILLER_211_2032 ();
 FILLCELL_X32 FILLER_211_2064 ();
 FILLCELL_X32 FILLER_211_2096 ();
 FILLCELL_X32 FILLER_211_2128 ();
 FILLCELL_X32 FILLER_211_2160 ();
 FILLCELL_X32 FILLER_211_2192 ();
 FILLCELL_X32 FILLER_211_2224 ();
 FILLCELL_X32 FILLER_211_2256 ();
 FILLCELL_X32 FILLER_211_2288 ();
 FILLCELL_X32 FILLER_211_2320 ();
 FILLCELL_X32 FILLER_211_2352 ();
 FILLCELL_X32 FILLER_211_2384 ();
 FILLCELL_X16 FILLER_211_2416 ();
 FILLCELL_X4 FILLER_211_2432 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_212_1784 ();
 FILLCELL_X32 FILLER_212_1816 ();
 FILLCELL_X32 FILLER_212_1848 ();
 FILLCELL_X8 FILLER_212_1880 ();
 FILLCELL_X4 FILLER_212_1888 ();
 FILLCELL_X2 FILLER_212_1892 ();
 FILLCELL_X32 FILLER_212_1895 ();
 FILLCELL_X32 FILLER_212_1927 ();
 FILLCELL_X32 FILLER_212_1959 ();
 FILLCELL_X32 FILLER_212_1991 ();
 FILLCELL_X32 FILLER_212_2023 ();
 FILLCELL_X32 FILLER_212_2055 ();
 FILLCELL_X32 FILLER_212_2087 ();
 FILLCELL_X32 FILLER_212_2119 ();
 FILLCELL_X32 FILLER_212_2151 ();
 FILLCELL_X32 FILLER_212_2183 ();
 FILLCELL_X32 FILLER_212_2215 ();
 FILLCELL_X32 FILLER_212_2247 ();
 FILLCELL_X32 FILLER_212_2279 ();
 FILLCELL_X32 FILLER_212_2311 ();
 FILLCELL_X32 FILLER_212_2343 ();
 FILLCELL_X32 FILLER_212_2375 ();
 FILLCELL_X16 FILLER_212_2407 ();
 FILLCELL_X8 FILLER_212_2423 ();
 FILLCELL_X4 FILLER_212_2431 ();
 FILLCELL_X1 FILLER_212_2435 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X32 FILLER_213_1776 ();
 FILLCELL_X32 FILLER_213_1808 ();
 FILLCELL_X32 FILLER_213_1840 ();
 FILLCELL_X32 FILLER_213_1872 ();
 FILLCELL_X32 FILLER_213_1904 ();
 FILLCELL_X32 FILLER_213_1936 ();
 FILLCELL_X32 FILLER_213_1968 ();
 FILLCELL_X32 FILLER_213_2000 ();
 FILLCELL_X32 FILLER_213_2032 ();
 FILLCELL_X32 FILLER_213_2064 ();
 FILLCELL_X32 FILLER_213_2096 ();
 FILLCELL_X32 FILLER_213_2128 ();
 FILLCELL_X32 FILLER_213_2160 ();
 FILLCELL_X32 FILLER_213_2192 ();
 FILLCELL_X32 FILLER_213_2224 ();
 FILLCELL_X32 FILLER_213_2256 ();
 FILLCELL_X32 FILLER_213_2288 ();
 FILLCELL_X32 FILLER_213_2320 ();
 FILLCELL_X32 FILLER_213_2352 ();
 FILLCELL_X32 FILLER_213_2384 ();
 FILLCELL_X16 FILLER_213_2416 ();
 FILLCELL_X4 FILLER_213_2432 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_214_1784 ();
 FILLCELL_X32 FILLER_214_1816 ();
 FILLCELL_X32 FILLER_214_1848 ();
 FILLCELL_X8 FILLER_214_1880 ();
 FILLCELL_X4 FILLER_214_1888 ();
 FILLCELL_X2 FILLER_214_1892 ();
 FILLCELL_X32 FILLER_214_1895 ();
 FILLCELL_X32 FILLER_214_1927 ();
 FILLCELL_X32 FILLER_214_1959 ();
 FILLCELL_X32 FILLER_214_1991 ();
 FILLCELL_X32 FILLER_214_2023 ();
 FILLCELL_X32 FILLER_214_2055 ();
 FILLCELL_X32 FILLER_214_2087 ();
 FILLCELL_X32 FILLER_214_2119 ();
 FILLCELL_X32 FILLER_214_2151 ();
 FILLCELL_X32 FILLER_214_2183 ();
 FILLCELL_X32 FILLER_214_2215 ();
 FILLCELL_X32 FILLER_214_2247 ();
 FILLCELL_X32 FILLER_214_2279 ();
 FILLCELL_X32 FILLER_214_2311 ();
 FILLCELL_X32 FILLER_214_2343 ();
 FILLCELL_X32 FILLER_214_2375 ();
 FILLCELL_X16 FILLER_214_2407 ();
 FILLCELL_X8 FILLER_214_2423 ();
 FILLCELL_X4 FILLER_214_2431 ();
 FILLCELL_X1 FILLER_214_2435 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X32 FILLER_215_1776 ();
 FILLCELL_X32 FILLER_215_1808 ();
 FILLCELL_X32 FILLER_215_1840 ();
 FILLCELL_X32 FILLER_215_1872 ();
 FILLCELL_X32 FILLER_215_1904 ();
 FILLCELL_X32 FILLER_215_1936 ();
 FILLCELL_X32 FILLER_215_1968 ();
 FILLCELL_X32 FILLER_215_2000 ();
 FILLCELL_X32 FILLER_215_2032 ();
 FILLCELL_X32 FILLER_215_2064 ();
 FILLCELL_X32 FILLER_215_2096 ();
 FILLCELL_X32 FILLER_215_2128 ();
 FILLCELL_X32 FILLER_215_2160 ();
 FILLCELL_X32 FILLER_215_2192 ();
 FILLCELL_X32 FILLER_215_2224 ();
 FILLCELL_X32 FILLER_215_2256 ();
 FILLCELL_X32 FILLER_215_2288 ();
 FILLCELL_X32 FILLER_215_2320 ();
 FILLCELL_X32 FILLER_215_2352 ();
 FILLCELL_X32 FILLER_215_2384 ();
 FILLCELL_X16 FILLER_215_2416 ();
 FILLCELL_X4 FILLER_215_2432 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X32 FILLER_216_1784 ();
 FILLCELL_X32 FILLER_216_1816 ();
 FILLCELL_X32 FILLER_216_1848 ();
 FILLCELL_X8 FILLER_216_1880 ();
 FILLCELL_X4 FILLER_216_1888 ();
 FILLCELL_X2 FILLER_216_1892 ();
 FILLCELL_X32 FILLER_216_1895 ();
 FILLCELL_X32 FILLER_216_1927 ();
 FILLCELL_X32 FILLER_216_1959 ();
 FILLCELL_X32 FILLER_216_1991 ();
 FILLCELL_X32 FILLER_216_2023 ();
 FILLCELL_X32 FILLER_216_2055 ();
 FILLCELL_X32 FILLER_216_2087 ();
 FILLCELL_X32 FILLER_216_2119 ();
 FILLCELL_X32 FILLER_216_2151 ();
 FILLCELL_X32 FILLER_216_2183 ();
 FILLCELL_X32 FILLER_216_2215 ();
 FILLCELL_X32 FILLER_216_2247 ();
 FILLCELL_X32 FILLER_216_2279 ();
 FILLCELL_X32 FILLER_216_2311 ();
 FILLCELL_X32 FILLER_216_2343 ();
 FILLCELL_X32 FILLER_216_2375 ();
 FILLCELL_X16 FILLER_216_2407 ();
 FILLCELL_X8 FILLER_216_2423 ();
 FILLCELL_X4 FILLER_216_2431 ();
 FILLCELL_X1 FILLER_216_2435 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X32 FILLER_217_1776 ();
 FILLCELL_X32 FILLER_217_1808 ();
 FILLCELL_X32 FILLER_217_1840 ();
 FILLCELL_X32 FILLER_217_1872 ();
 FILLCELL_X32 FILLER_217_1904 ();
 FILLCELL_X32 FILLER_217_1936 ();
 FILLCELL_X32 FILLER_217_1968 ();
 FILLCELL_X32 FILLER_217_2000 ();
 FILLCELL_X32 FILLER_217_2032 ();
 FILLCELL_X32 FILLER_217_2064 ();
 FILLCELL_X32 FILLER_217_2096 ();
 FILLCELL_X32 FILLER_217_2128 ();
 FILLCELL_X32 FILLER_217_2160 ();
 FILLCELL_X32 FILLER_217_2192 ();
 FILLCELL_X32 FILLER_217_2224 ();
 FILLCELL_X32 FILLER_217_2256 ();
 FILLCELL_X32 FILLER_217_2288 ();
 FILLCELL_X32 FILLER_217_2320 ();
 FILLCELL_X32 FILLER_217_2352 ();
 FILLCELL_X32 FILLER_217_2384 ();
 FILLCELL_X16 FILLER_217_2416 ();
 FILLCELL_X4 FILLER_217_2432 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_218_1784 ();
 FILLCELL_X32 FILLER_218_1816 ();
 FILLCELL_X32 FILLER_218_1848 ();
 FILLCELL_X8 FILLER_218_1880 ();
 FILLCELL_X4 FILLER_218_1888 ();
 FILLCELL_X2 FILLER_218_1892 ();
 FILLCELL_X32 FILLER_218_1895 ();
 FILLCELL_X32 FILLER_218_1927 ();
 FILLCELL_X32 FILLER_218_1959 ();
 FILLCELL_X32 FILLER_218_1991 ();
 FILLCELL_X32 FILLER_218_2023 ();
 FILLCELL_X32 FILLER_218_2055 ();
 FILLCELL_X32 FILLER_218_2087 ();
 FILLCELL_X32 FILLER_218_2119 ();
 FILLCELL_X32 FILLER_218_2151 ();
 FILLCELL_X32 FILLER_218_2183 ();
 FILLCELL_X32 FILLER_218_2215 ();
 FILLCELL_X32 FILLER_218_2247 ();
 FILLCELL_X32 FILLER_218_2279 ();
 FILLCELL_X32 FILLER_218_2311 ();
 FILLCELL_X32 FILLER_218_2343 ();
 FILLCELL_X32 FILLER_218_2375 ();
 FILLCELL_X16 FILLER_218_2407 ();
 FILLCELL_X8 FILLER_218_2423 ();
 FILLCELL_X4 FILLER_218_2431 ();
 FILLCELL_X1 FILLER_218_2435 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X32 FILLER_219_1776 ();
 FILLCELL_X32 FILLER_219_1808 ();
 FILLCELL_X32 FILLER_219_1840 ();
 FILLCELL_X32 FILLER_219_1872 ();
 FILLCELL_X32 FILLER_219_1904 ();
 FILLCELL_X32 FILLER_219_1936 ();
 FILLCELL_X32 FILLER_219_1968 ();
 FILLCELL_X32 FILLER_219_2000 ();
 FILLCELL_X32 FILLER_219_2032 ();
 FILLCELL_X32 FILLER_219_2064 ();
 FILLCELL_X32 FILLER_219_2096 ();
 FILLCELL_X32 FILLER_219_2128 ();
 FILLCELL_X32 FILLER_219_2160 ();
 FILLCELL_X32 FILLER_219_2192 ();
 FILLCELL_X32 FILLER_219_2224 ();
 FILLCELL_X32 FILLER_219_2256 ();
 FILLCELL_X32 FILLER_219_2288 ();
 FILLCELL_X32 FILLER_219_2320 ();
 FILLCELL_X32 FILLER_219_2352 ();
 FILLCELL_X32 FILLER_219_2384 ();
 FILLCELL_X16 FILLER_219_2416 ();
 FILLCELL_X4 FILLER_219_2432 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_220_1784 ();
 FILLCELL_X32 FILLER_220_1816 ();
 FILLCELL_X32 FILLER_220_1848 ();
 FILLCELL_X8 FILLER_220_1880 ();
 FILLCELL_X4 FILLER_220_1888 ();
 FILLCELL_X2 FILLER_220_1892 ();
 FILLCELL_X32 FILLER_220_1895 ();
 FILLCELL_X32 FILLER_220_1927 ();
 FILLCELL_X32 FILLER_220_1959 ();
 FILLCELL_X32 FILLER_220_1991 ();
 FILLCELL_X32 FILLER_220_2023 ();
 FILLCELL_X32 FILLER_220_2055 ();
 FILLCELL_X32 FILLER_220_2087 ();
 FILLCELL_X32 FILLER_220_2119 ();
 FILLCELL_X32 FILLER_220_2151 ();
 FILLCELL_X32 FILLER_220_2183 ();
 FILLCELL_X32 FILLER_220_2215 ();
 FILLCELL_X32 FILLER_220_2247 ();
 FILLCELL_X32 FILLER_220_2279 ();
 FILLCELL_X32 FILLER_220_2311 ();
 FILLCELL_X32 FILLER_220_2343 ();
 FILLCELL_X32 FILLER_220_2375 ();
 FILLCELL_X16 FILLER_220_2407 ();
 FILLCELL_X8 FILLER_220_2423 ();
 FILLCELL_X4 FILLER_220_2431 ();
 FILLCELL_X1 FILLER_220_2435 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X32 FILLER_221_1776 ();
 FILLCELL_X32 FILLER_221_1808 ();
 FILLCELL_X32 FILLER_221_1840 ();
 FILLCELL_X32 FILLER_221_1872 ();
 FILLCELL_X32 FILLER_221_1904 ();
 FILLCELL_X32 FILLER_221_1936 ();
 FILLCELL_X32 FILLER_221_1968 ();
 FILLCELL_X32 FILLER_221_2000 ();
 FILLCELL_X32 FILLER_221_2032 ();
 FILLCELL_X32 FILLER_221_2064 ();
 FILLCELL_X32 FILLER_221_2096 ();
 FILLCELL_X32 FILLER_221_2128 ();
 FILLCELL_X32 FILLER_221_2160 ();
 FILLCELL_X32 FILLER_221_2192 ();
 FILLCELL_X32 FILLER_221_2224 ();
 FILLCELL_X32 FILLER_221_2256 ();
 FILLCELL_X32 FILLER_221_2288 ();
 FILLCELL_X32 FILLER_221_2320 ();
 FILLCELL_X32 FILLER_221_2352 ();
 FILLCELL_X32 FILLER_221_2384 ();
 FILLCELL_X16 FILLER_221_2416 ();
 FILLCELL_X4 FILLER_221_2432 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_222_1784 ();
 FILLCELL_X32 FILLER_222_1816 ();
 FILLCELL_X32 FILLER_222_1848 ();
 FILLCELL_X8 FILLER_222_1880 ();
 FILLCELL_X4 FILLER_222_1888 ();
 FILLCELL_X2 FILLER_222_1892 ();
 FILLCELL_X32 FILLER_222_1895 ();
 FILLCELL_X32 FILLER_222_1927 ();
 FILLCELL_X32 FILLER_222_1959 ();
 FILLCELL_X32 FILLER_222_1991 ();
 FILLCELL_X32 FILLER_222_2023 ();
 FILLCELL_X32 FILLER_222_2055 ();
 FILLCELL_X32 FILLER_222_2087 ();
 FILLCELL_X32 FILLER_222_2119 ();
 FILLCELL_X32 FILLER_222_2151 ();
 FILLCELL_X32 FILLER_222_2183 ();
 FILLCELL_X32 FILLER_222_2215 ();
 FILLCELL_X32 FILLER_222_2247 ();
 FILLCELL_X32 FILLER_222_2279 ();
 FILLCELL_X32 FILLER_222_2311 ();
 FILLCELL_X32 FILLER_222_2343 ();
 FILLCELL_X32 FILLER_222_2375 ();
 FILLCELL_X16 FILLER_222_2407 ();
 FILLCELL_X8 FILLER_222_2423 ();
 FILLCELL_X4 FILLER_222_2431 ();
 FILLCELL_X1 FILLER_222_2435 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X32 FILLER_223_1776 ();
 FILLCELL_X32 FILLER_223_1808 ();
 FILLCELL_X32 FILLER_223_1840 ();
 FILLCELL_X32 FILLER_223_1872 ();
 FILLCELL_X32 FILLER_223_1904 ();
 FILLCELL_X32 FILLER_223_1936 ();
 FILLCELL_X32 FILLER_223_1968 ();
 FILLCELL_X32 FILLER_223_2000 ();
 FILLCELL_X32 FILLER_223_2032 ();
 FILLCELL_X32 FILLER_223_2064 ();
 FILLCELL_X32 FILLER_223_2096 ();
 FILLCELL_X32 FILLER_223_2128 ();
 FILLCELL_X32 FILLER_223_2160 ();
 FILLCELL_X32 FILLER_223_2192 ();
 FILLCELL_X32 FILLER_223_2224 ();
 FILLCELL_X32 FILLER_223_2256 ();
 FILLCELL_X32 FILLER_223_2288 ();
 FILLCELL_X32 FILLER_223_2320 ();
 FILLCELL_X32 FILLER_223_2352 ();
 FILLCELL_X32 FILLER_223_2384 ();
 FILLCELL_X16 FILLER_223_2416 ();
 FILLCELL_X4 FILLER_223_2432 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_224_1784 ();
 FILLCELL_X32 FILLER_224_1816 ();
 FILLCELL_X32 FILLER_224_1848 ();
 FILLCELL_X8 FILLER_224_1880 ();
 FILLCELL_X4 FILLER_224_1888 ();
 FILLCELL_X2 FILLER_224_1892 ();
 FILLCELL_X32 FILLER_224_1895 ();
 FILLCELL_X32 FILLER_224_1927 ();
 FILLCELL_X32 FILLER_224_1959 ();
 FILLCELL_X32 FILLER_224_1991 ();
 FILLCELL_X32 FILLER_224_2023 ();
 FILLCELL_X32 FILLER_224_2055 ();
 FILLCELL_X32 FILLER_224_2087 ();
 FILLCELL_X32 FILLER_224_2119 ();
 FILLCELL_X32 FILLER_224_2151 ();
 FILLCELL_X32 FILLER_224_2183 ();
 FILLCELL_X32 FILLER_224_2215 ();
 FILLCELL_X32 FILLER_224_2247 ();
 FILLCELL_X32 FILLER_224_2279 ();
 FILLCELL_X32 FILLER_224_2311 ();
 FILLCELL_X32 FILLER_224_2343 ();
 FILLCELL_X32 FILLER_224_2375 ();
 FILLCELL_X16 FILLER_224_2407 ();
 FILLCELL_X8 FILLER_224_2423 ();
 FILLCELL_X4 FILLER_224_2431 ();
 FILLCELL_X1 FILLER_224_2435 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X32 FILLER_225_1776 ();
 FILLCELL_X32 FILLER_225_1808 ();
 FILLCELL_X32 FILLER_225_1840 ();
 FILLCELL_X32 FILLER_225_1872 ();
 FILLCELL_X32 FILLER_225_1904 ();
 FILLCELL_X32 FILLER_225_1936 ();
 FILLCELL_X32 FILLER_225_1968 ();
 FILLCELL_X32 FILLER_225_2000 ();
 FILLCELL_X32 FILLER_225_2032 ();
 FILLCELL_X32 FILLER_225_2064 ();
 FILLCELL_X32 FILLER_225_2096 ();
 FILLCELL_X32 FILLER_225_2128 ();
 FILLCELL_X32 FILLER_225_2160 ();
 FILLCELL_X32 FILLER_225_2192 ();
 FILLCELL_X32 FILLER_225_2224 ();
 FILLCELL_X32 FILLER_225_2256 ();
 FILLCELL_X32 FILLER_225_2288 ();
 FILLCELL_X32 FILLER_225_2320 ();
 FILLCELL_X32 FILLER_225_2352 ();
 FILLCELL_X32 FILLER_225_2384 ();
 FILLCELL_X16 FILLER_225_2416 ();
 FILLCELL_X4 FILLER_225_2432 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_226_1784 ();
 FILLCELL_X32 FILLER_226_1816 ();
 FILLCELL_X32 FILLER_226_1848 ();
 FILLCELL_X8 FILLER_226_1880 ();
 FILLCELL_X4 FILLER_226_1888 ();
 FILLCELL_X2 FILLER_226_1892 ();
 FILLCELL_X32 FILLER_226_1895 ();
 FILLCELL_X32 FILLER_226_1927 ();
 FILLCELL_X32 FILLER_226_1959 ();
 FILLCELL_X32 FILLER_226_1991 ();
 FILLCELL_X32 FILLER_226_2023 ();
 FILLCELL_X32 FILLER_226_2055 ();
 FILLCELL_X32 FILLER_226_2087 ();
 FILLCELL_X32 FILLER_226_2119 ();
 FILLCELL_X32 FILLER_226_2151 ();
 FILLCELL_X32 FILLER_226_2183 ();
 FILLCELL_X32 FILLER_226_2215 ();
 FILLCELL_X32 FILLER_226_2247 ();
 FILLCELL_X32 FILLER_226_2279 ();
 FILLCELL_X32 FILLER_226_2311 ();
 FILLCELL_X32 FILLER_226_2343 ();
 FILLCELL_X32 FILLER_226_2375 ();
 FILLCELL_X16 FILLER_226_2407 ();
 FILLCELL_X8 FILLER_226_2423 ();
 FILLCELL_X4 FILLER_226_2431 ();
 FILLCELL_X1 FILLER_226_2435 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X32 FILLER_227_1776 ();
 FILLCELL_X32 FILLER_227_1808 ();
 FILLCELL_X32 FILLER_227_1840 ();
 FILLCELL_X32 FILLER_227_1872 ();
 FILLCELL_X32 FILLER_227_1904 ();
 FILLCELL_X32 FILLER_227_1936 ();
 FILLCELL_X32 FILLER_227_1968 ();
 FILLCELL_X32 FILLER_227_2000 ();
 FILLCELL_X32 FILLER_227_2032 ();
 FILLCELL_X32 FILLER_227_2064 ();
 FILLCELL_X32 FILLER_227_2096 ();
 FILLCELL_X32 FILLER_227_2128 ();
 FILLCELL_X32 FILLER_227_2160 ();
 FILLCELL_X32 FILLER_227_2192 ();
 FILLCELL_X32 FILLER_227_2224 ();
 FILLCELL_X32 FILLER_227_2256 ();
 FILLCELL_X32 FILLER_227_2288 ();
 FILLCELL_X32 FILLER_227_2320 ();
 FILLCELL_X32 FILLER_227_2352 ();
 FILLCELL_X32 FILLER_227_2384 ();
 FILLCELL_X16 FILLER_227_2416 ();
 FILLCELL_X4 FILLER_227_2432 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_228_1784 ();
 FILLCELL_X32 FILLER_228_1816 ();
 FILLCELL_X32 FILLER_228_1848 ();
 FILLCELL_X8 FILLER_228_1880 ();
 FILLCELL_X4 FILLER_228_1888 ();
 FILLCELL_X2 FILLER_228_1892 ();
 FILLCELL_X32 FILLER_228_1895 ();
 FILLCELL_X32 FILLER_228_1927 ();
 FILLCELL_X32 FILLER_228_1959 ();
 FILLCELL_X32 FILLER_228_1991 ();
 FILLCELL_X32 FILLER_228_2023 ();
 FILLCELL_X32 FILLER_228_2055 ();
 FILLCELL_X32 FILLER_228_2087 ();
 FILLCELL_X32 FILLER_228_2119 ();
 FILLCELL_X32 FILLER_228_2151 ();
 FILLCELL_X32 FILLER_228_2183 ();
 FILLCELL_X32 FILLER_228_2215 ();
 FILLCELL_X32 FILLER_228_2247 ();
 FILLCELL_X32 FILLER_228_2279 ();
 FILLCELL_X32 FILLER_228_2311 ();
 FILLCELL_X32 FILLER_228_2343 ();
 FILLCELL_X32 FILLER_228_2375 ();
 FILLCELL_X16 FILLER_228_2407 ();
 FILLCELL_X8 FILLER_228_2423 ();
 FILLCELL_X4 FILLER_228_2431 ();
 FILLCELL_X1 FILLER_228_2435 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X32 FILLER_229_1776 ();
 FILLCELL_X32 FILLER_229_1808 ();
 FILLCELL_X32 FILLER_229_1840 ();
 FILLCELL_X32 FILLER_229_1872 ();
 FILLCELL_X32 FILLER_229_1904 ();
 FILLCELL_X32 FILLER_229_1936 ();
 FILLCELL_X32 FILLER_229_1968 ();
 FILLCELL_X32 FILLER_229_2000 ();
 FILLCELL_X32 FILLER_229_2032 ();
 FILLCELL_X32 FILLER_229_2064 ();
 FILLCELL_X32 FILLER_229_2096 ();
 FILLCELL_X32 FILLER_229_2128 ();
 FILLCELL_X32 FILLER_229_2160 ();
 FILLCELL_X32 FILLER_229_2192 ();
 FILLCELL_X32 FILLER_229_2224 ();
 FILLCELL_X32 FILLER_229_2256 ();
 FILLCELL_X32 FILLER_229_2288 ();
 FILLCELL_X32 FILLER_229_2320 ();
 FILLCELL_X32 FILLER_229_2352 ();
 FILLCELL_X32 FILLER_229_2384 ();
 FILLCELL_X16 FILLER_229_2416 ();
 FILLCELL_X4 FILLER_229_2432 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_230_1784 ();
 FILLCELL_X32 FILLER_230_1816 ();
 FILLCELL_X32 FILLER_230_1848 ();
 FILLCELL_X8 FILLER_230_1880 ();
 FILLCELL_X4 FILLER_230_1888 ();
 FILLCELL_X2 FILLER_230_1892 ();
 FILLCELL_X32 FILLER_230_1895 ();
 FILLCELL_X32 FILLER_230_1927 ();
 FILLCELL_X32 FILLER_230_1959 ();
 FILLCELL_X32 FILLER_230_1991 ();
 FILLCELL_X32 FILLER_230_2023 ();
 FILLCELL_X32 FILLER_230_2055 ();
 FILLCELL_X32 FILLER_230_2087 ();
 FILLCELL_X32 FILLER_230_2119 ();
 FILLCELL_X32 FILLER_230_2151 ();
 FILLCELL_X32 FILLER_230_2183 ();
 FILLCELL_X32 FILLER_230_2215 ();
 FILLCELL_X32 FILLER_230_2247 ();
 FILLCELL_X32 FILLER_230_2279 ();
 FILLCELL_X32 FILLER_230_2311 ();
 FILLCELL_X32 FILLER_230_2343 ();
 FILLCELL_X32 FILLER_230_2375 ();
 FILLCELL_X16 FILLER_230_2407 ();
 FILLCELL_X8 FILLER_230_2423 ();
 FILLCELL_X4 FILLER_230_2431 ();
 FILLCELL_X1 FILLER_230_2435 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X32 FILLER_231_1776 ();
 FILLCELL_X32 FILLER_231_1808 ();
 FILLCELL_X32 FILLER_231_1840 ();
 FILLCELL_X32 FILLER_231_1872 ();
 FILLCELL_X32 FILLER_231_1904 ();
 FILLCELL_X32 FILLER_231_1936 ();
 FILLCELL_X32 FILLER_231_1968 ();
 FILLCELL_X32 FILLER_231_2000 ();
 FILLCELL_X32 FILLER_231_2032 ();
 FILLCELL_X32 FILLER_231_2064 ();
 FILLCELL_X32 FILLER_231_2096 ();
 FILLCELL_X32 FILLER_231_2128 ();
 FILLCELL_X32 FILLER_231_2160 ();
 FILLCELL_X32 FILLER_231_2192 ();
 FILLCELL_X32 FILLER_231_2224 ();
 FILLCELL_X32 FILLER_231_2256 ();
 FILLCELL_X32 FILLER_231_2288 ();
 FILLCELL_X32 FILLER_231_2320 ();
 FILLCELL_X32 FILLER_231_2352 ();
 FILLCELL_X32 FILLER_231_2384 ();
 FILLCELL_X16 FILLER_231_2416 ();
 FILLCELL_X4 FILLER_231_2432 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X32 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_232_1784 ();
 FILLCELL_X32 FILLER_232_1816 ();
 FILLCELL_X32 FILLER_232_1848 ();
 FILLCELL_X8 FILLER_232_1880 ();
 FILLCELL_X4 FILLER_232_1888 ();
 FILLCELL_X2 FILLER_232_1892 ();
 FILLCELL_X32 FILLER_232_1895 ();
 FILLCELL_X32 FILLER_232_1927 ();
 FILLCELL_X32 FILLER_232_1959 ();
 FILLCELL_X32 FILLER_232_1991 ();
 FILLCELL_X32 FILLER_232_2023 ();
 FILLCELL_X32 FILLER_232_2055 ();
 FILLCELL_X32 FILLER_232_2087 ();
 FILLCELL_X32 FILLER_232_2119 ();
 FILLCELL_X32 FILLER_232_2151 ();
 FILLCELL_X32 FILLER_232_2183 ();
 FILLCELL_X32 FILLER_232_2215 ();
 FILLCELL_X32 FILLER_232_2247 ();
 FILLCELL_X32 FILLER_232_2279 ();
 FILLCELL_X32 FILLER_232_2311 ();
 FILLCELL_X32 FILLER_232_2343 ();
 FILLCELL_X32 FILLER_232_2375 ();
 FILLCELL_X16 FILLER_232_2407 ();
 FILLCELL_X8 FILLER_232_2423 ();
 FILLCELL_X4 FILLER_232_2431 ();
 FILLCELL_X1 FILLER_232_2435 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X32 FILLER_233_1776 ();
 FILLCELL_X32 FILLER_233_1808 ();
 FILLCELL_X32 FILLER_233_1840 ();
 FILLCELL_X32 FILLER_233_1872 ();
 FILLCELL_X32 FILLER_233_1904 ();
 FILLCELL_X32 FILLER_233_1936 ();
 FILLCELL_X32 FILLER_233_1968 ();
 FILLCELL_X32 FILLER_233_2000 ();
 FILLCELL_X32 FILLER_233_2032 ();
 FILLCELL_X32 FILLER_233_2064 ();
 FILLCELL_X32 FILLER_233_2096 ();
 FILLCELL_X32 FILLER_233_2128 ();
 FILLCELL_X32 FILLER_233_2160 ();
 FILLCELL_X32 FILLER_233_2192 ();
 FILLCELL_X32 FILLER_233_2224 ();
 FILLCELL_X32 FILLER_233_2256 ();
 FILLCELL_X32 FILLER_233_2288 ();
 FILLCELL_X32 FILLER_233_2320 ();
 FILLCELL_X32 FILLER_233_2352 ();
 FILLCELL_X32 FILLER_233_2384 ();
 FILLCELL_X16 FILLER_233_2416 ();
 FILLCELL_X4 FILLER_233_2432 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X32 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_234_1784 ();
 FILLCELL_X32 FILLER_234_1816 ();
 FILLCELL_X32 FILLER_234_1848 ();
 FILLCELL_X8 FILLER_234_1880 ();
 FILLCELL_X4 FILLER_234_1888 ();
 FILLCELL_X2 FILLER_234_1892 ();
 FILLCELL_X32 FILLER_234_1895 ();
 FILLCELL_X32 FILLER_234_1927 ();
 FILLCELL_X32 FILLER_234_1959 ();
 FILLCELL_X32 FILLER_234_1991 ();
 FILLCELL_X32 FILLER_234_2023 ();
 FILLCELL_X32 FILLER_234_2055 ();
 FILLCELL_X32 FILLER_234_2087 ();
 FILLCELL_X32 FILLER_234_2119 ();
 FILLCELL_X32 FILLER_234_2151 ();
 FILLCELL_X32 FILLER_234_2183 ();
 FILLCELL_X32 FILLER_234_2215 ();
 FILLCELL_X32 FILLER_234_2247 ();
 FILLCELL_X32 FILLER_234_2279 ();
 FILLCELL_X32 FILLER_234_2311 ();
 FILLCELL_X32 FILLER_234_2343 ();
 FILLCELL_X32 FILLER_234_2375 ();
 FILLCELL_X16 FILLER_234_2407 ();
 FILLCELL_X8 FILLER_234_2423 ();
 FILLCELL_X4 FILLER_234_2431 ();
 FILLCELL_X1 FILLER_234_2435 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X32 FILLER_235_1776 ();
 FILLCELL_X32 FILLER_235_1808 ();
 FILLCELL_X32 FILLER_235_1840 ();
 FILLCELL_X32 FILLER_235_1872 ();
 FILLCELL_X32 FILLER_235_1904 ();
 FILLCELL_X32 FILLER_235_1936 ();
 FILLCELL_X32 FILLER_235_1968 ();
 FILLCELL_X32 FILLER_235_2000 ();
 FILLCELL_X32 FILLER_235_2032 ();
 FILLCELL_X32 FILLER_235_2064 ();
 FILLCELL_X32 FILLER_235_2096 ();
 FILLCELL_X32 FILLER_235_2128 ();
 FILLCELL_X32 FILLER_235_2160 ();
 FILLCELL_X32 FILLER_235_2192 ();
 FILLCELL_X32 FILLER_235_2224 ();
 FILLCELL_X32 FILLER_235_2256 ();
 FILLCELL_X32 FILLER_235_2288 ();
 FILLCELL_X32 FILLER_235_2320 ();
 FILLCELL_X32 FILLER_235_2352 ();
 FILLCELL_X32 FILLER_235_2384 ();
 FILLCELL_X16 FILLER_235_2416 ();
 FILLCELL_X4 FILLER_235_2432 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X32 FILLER_236_1752 ();
 FILLCELL_X32 FILLER_236_1784 ();
 FILLCELL_X32 FILLER_236_1816 ();
 FILLCELL_X32 FILLER_236_1848 ();
 FILLCELL_X8 FILLER_236_1880 ();
 FILLCELL_X4 FILLER_236_1888 ();
 FILLCELL_X2 FILLER_236_1892 ();
 FILLCELL_X32 FILLER_236_1895 ();
 FILLCELL_X32 FILLER_236_1927 ();
 FILLCELL_X32 FILLER_236_1959 ();
 FILLCELL_X32 FILLER_236_1991 ();
 FILLCELL_X32 FILLER_236_2023 ();
 FILLCELL_X32 FILLER_236_2055 ();
 FILLCELL_X32 FILLER_236_2087 ();
 FILLCELL_X32 FILLER_236_2119 ();
 FILLCELL_X32 FILLER_236_2151 ();
 FILLCELL_X32 FILLER_236_2183 ();
 FILLCELL_X32 FILLER_236_2215 ();
 FILLCELL_X32 FILLER_236_2247 ();
 FILLCELL_X32 FILLER_236_2279 ();
 FILLCELL_X32 FILLER_236_2311 ();
 FILLCELL_X32 FILLER_236_2343 ();
 FILLCELL_X32 FILLER_236_2375 ();
 FILLCELL_X16 FILLER_236_2407 ();
 FILLCELL_X8 FILLER_236_2423 ();
 FILLCELL_X4 FILLER_236_2431 ();
 FILLCELL_X1 FILLER_236_2435 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X32 FILLER_237_865 ();
 FILLCELL_X32 FILLER_237_897 ();
 FILLCELL_X32 FILLER_237_929 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X32 FILLER_237_1776 ();
 FILLCELL_X32 FILLER_237_1808 ();
 FILLCELL_X32 FILLER_237_1840 ();
 FILLCELL_X32 FILLER_237_1872 ();
 FILLCELL_X32 FILLER_237_1904 ();
 FILLCELL_X32 FILLER_237_1936 ();
 FILLCELL_X32 FILLER_237_1968 ();
 FILLCELL_X32 FILLER_237_2000 ();
 FILLCELL_X32 FILLER_237_2032 ();
 FILLCELL_X32 FILLER_237_2064 ();
 FILLCELL_X32 FILLER_237_2096 ();
 FILLCELL_X32 FILLER_237_2128 ();
 FILLCELL_X32 FILLER_237_2160 ();
 FILLCELL_X32 FILLER_237_2192 ();
 FILLCELL_X32 FILLER_237_2224 ();
 FILLCELL_X32 FILLER_237_2256 ();
 FILLCELL_X32 FILLER_237_2288 ();
 FILLCELL_X32 FILLER_237_2320 ();
 FILLCELL_X32 FILLER_237_2352 ();
 FILLCELL_X32 FILLER_237_2384 ();
 FILLCELL_X16 FILLER_237_2416 ();
 FILLCELL_X4 FILLER_237_2432 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X32 FILLER_238_856 ();
 FILLCELL_X32 FILLER_238_888 ();
 FILLCELL_X32 FILLER_238_920 ();
 FILLCELL_X32 FILLER_238_952 ();
 FILLCELL_X32 FILLER_238_984 ();
 FILLCELL_X32 FILLER_238_1016 ();
 FILLCELL_X32 FILLER_238_1048 ();
 FILLCELL_X32 FILLER_238_1080 ();
 FILLCELL_X32 FILLER_238_1112 ();
 FILLCELL_X32 FILLER_238_1144 ();
 FILLCELL_X32 FILLER_238_1176 ();
 FILLCELL_X32 FILLER_238_1208 ();
 FILLCELL_X32 FILLER_238_1240 ();
 FILLCELL_X32 FILLER_238_1272 ();
 FILLCELL_X32 FILLER_238_1304 ();
 FILLCELL_X32 FILLER_238_1336 ();
 FILLCELL_X32 FILLER_238_1368 ();
 FILLCELL_X32 FILLER_238_1400 ();
 FILLCELL_X32 FILLER_238_1432 ();
 FILLCELL_X32 FILLER_238_1464 ();
 FILLCELL_X32 FILLER_238_1496 ();
 FILLCELL_X32 FILLER_238_1528 ();
 FILLCELL_X32 FILLER_238_1560 ();
 FILLCELL_X32 FILLER_238_1592 ();
 FILLCELL_X32 FILLER_238_1624 ();
 FILLCELL_X32 FILLER_238_1656 ();
 FILLCELL_X32 FILLER_238_1688 ();
 FILLCELL_X32 FILLER_238_1720 ();
 FILLCELL_X32 FILLER_238_1752 ();
 FILLCELL_X32 FILLER_238_1784 ();
 FILLCELL_X32 FILLER_238_1816 ();
 FILLCELL_X32 FILLER_238_1848 ();
 FILLCELL_X8 FILLER_238_1880 ();
 FILLCELL_X4 FILLER_238_1888 ();
 FILLCELL_X2 FILLER_238_1892 ();
 FILLCELL_X32 FILLER_238_1895 ();
 FILLCELL_X32 FILLER_238_1927 ();
 FILLCELL_X32 FILLER_238_1959 ();
 FILLCELL_X32 FILLER_238_1991 ();
 FILLCELL_X32 FILLER_238_2023 ();
 FILLCELL_X32 FILLER_238_2055 ();
 FILLCELL_X32 FILLER_238_2087 ();
 FILLCELL_X32 FILLER_238_2119 ();
 FILLCELL_X32 FILLER_238_2151 ();
 FILLCELL_X32 FILLER_238_2183 ();
 FILLCELL_X32 FILLER_238_2215 ();
 FILLCELL_X32 FILLER_238_2247 ();
 FILLCELL_X32 FILLER_238_2279 ();
 FILLCELL_X32 FILLER_238_2311 ();
 FILLCELL_X32 FILLER_238_2343 ();
 FILLCELL_X32 FILLER_238_2375 ();
 FILLCELL_X16 FILLER_238_2407 ();
 FILLCELL_X8 FILLER_238_2423 ();
 FILLCELL_X4 FILLER_238_2431 ();
 FILLCELL_X1 FILLER_238_2435 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X32 FILLER_239_833 ();
 FILLCELL_X32 FILLER_239_865 ();
 FILLCELL_X32 FILLER_239_897 ();
 FILLCELL_X32 FILLER_239_929 ();
 FILLCELL_X32 FILLER_239_961 ();
 FILLCELL_X32 FILLER_239_993 ();
 FILLCELL_X32 FILLER_239_1025 ();
 FILLCELL_X32 FILLER_239_1057 ();
 FILLCELL_X32 FILLER_239_1089 ();
 FILLCELL_X32 FILLER_239_1121 ();
 FILLCELL_X32 FILLER_239_1153 ();
 FILLCELL_X32 FILLER_239_1185 ();
 FILLCELL_X32 FILLER_239_1217 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X32 FILLER_239_1776 ();
 FILLCELL_X32 FILLER_239_1808 ();
 FILLCELL_X32 FILLER_239_1840 ();
 FILLCELL_X32 FILLER_239_1872 ();
 FILLCELL_X32 FILLER_239_1904 ();
 FILLCELL_X32 FILLER_239_1936 ();
 FILLCELL_X32 FILLER_239_1968 ();
 FILLCELL_X32 FILLER_239_2000 ();
 FILLCELL_X32 FILLER_239_2032 ();
 FILLCELL_X32 FILLER_239_2064 ();
 FILLCELL_X32 FILLER_239_2096 ();
 FILLCELL_X32 FILLER_239_2128 ();
 FILLCELL_X32 FILLER_239_2160 ();
 FILLCELL_X32 FILLER_239_2192 ();
 FILLCELL_X32 FILLER_239_2224 ();
 FILLCELL_X32 FILLER_239_2256 ();
 FILLCELL_X32 FILLER_239_2288 ();
 FILLCELL_X32 FILLER_239_2320 ();
 FILLCELL_X32 FILLER_239_2352 ();
 FILLCELL_X32 FILLER_239_2384 ();
 FILLCELL_X16 FILLER_239_2416 ();
 FILLCELL_X4 FILLER_239_2432 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X32 FILLER_240_824 ();
 FILLCELL_X32 FILLER_240_856 ();
 FILLCELL_X32 FILLER_240_888 ();
 FILLCELL_X32 FILLER_240_920 ();
 FILLCELL_X32 FILLER_240_952 ();
 FILLCELL_X32 FILLER_240_984 ();
 FILLCELL_X32 FILLER_240_1016 ();
 FILLCELL_X32 FILLER_240_1048 ();
 FILLCELL_X32 FILLER_240_1080 ();
 FILLCELL_X32 FILLER_240_1112 ();
 FILLCELL_X32 FILLER_240_1144 ();
 FILLCELL_X32 FILLER_240_1176 ();
 FILLCELL_X32 FILLER_240_1208 ();
 FILLCELL_X32 FILLER_240_1240 ();
 FILLCELL_X32 FILLER_240_1272 ();
 FILLCELL_X32 FILLER_240_1304 ();
 FILLCELL_X32 FILLER_240_1336 ();
 FILLCELL_X32 FILLER_240_1368 ();
 FILLCELL_X32 FILLER_240_1400 ();
 FILLCELL_X32 FILLER_240_1432 ();
 FILLCELL_X32 FILLER_240_1464 ();
 FILLCELL_X32 FILLER_240_1496 ();
 FILLCELL_X32 FILLER_240_1528 ();
 FILLCELL_X32 FILLER_240_1560 ();
 FILLCELL_X32 FILLER_240_1592 ();
 FILLCELL_X32 FILLER_240_1624 ();
 FILLCELL_X32 FILLER_240_1656 ();
 FILLCELL_X32 FILLER_240_1688 ();
 FILLCELL_X32 FILLER_240_1720 ();
 FILLCELL_X32 FILLER_240_1752 ();
 FILLCELL_X32 FILLER_240_1784 ();
 FILLCELL_X32 FILLER_240_1816 ();
 FILLCELL_X32 FILLER_240_1848 ();
 FILLCELL_X8 FILLER_240_1880 ();
 FILLCELL_X4 FILLER_240_1888 ();
 FILLCELL_X2 FILLER_240_1892 ();
 FILLCELL_X32 FILLER_240_1895 ();
 FILLCELL_X32 FILLER_240_1927 ();
 FILLCELL_X32 FILLER_240_1959 ();
 FILLCELL_X32 FILLER_240_1991 ();
 FILLCELL_X32 FILLER_240_2023 ();
 FILLCELL_X32 FILLER_240_2055 ();
 FILLCELL_X32 FILLER_240_2087 ();
 FILLCELL_X32 FILLER_240_2119 ();
 FILLCELL_X32 FILLER_240_2151 ();
 FILLCELL_X32 FILLER_240_2183 ();
 FILLCELL_X32 FILLER_240_2215 ();
 FILLCELL_X32 FILLER_240_2247 ();
 FILLCELL_X32 FILLER_240_2279 ();
 FILLCELL_X32 FILLER_240_2311 ();
 FILLCELL_X32 FILLER_240_2343 ();
 FILLCELL_X32 FILLER_240_2375 ();
 FILLCELL_X16 FILLER_240_2407 ();
 FILLCELL_X8 FILLER_240_2423 ();
 FILLCELL_X4 FILLER_240_2431 ();
 FILLCELL_X1 FILLER_240_2435 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X32 FILLER_241_833 ();
 FILLCELL_X32 FILLER_241_865 ();
 FILLCELL_X32 FILLER_241_897 ();
 FILLCELL_X32 FILLER_241_929 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X32 FILLER_241_993 ();
 FILLCELL_X32 FILLER_241_1025 ();
 FILLCELL_X32 FILLER_241_1057 ();
 FILLCELL_X32 FILLER_241_1089 ();
 FILLCELL_X32 FILLER_241_1121 ();
 FILLCELL_X32 FILLER_241_1153 ();
 FILLCELL_X32 FILLER_241_1185 ();
 FILLCELL_X32 FILLER_241_1217 ();
 FILLCELL_X8 FILLER_241_1249 ();
 FILLCELL_X4 FILLER_241_1257 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X32 FILLER_241_1776 ();
 FILLCELL_X32 FILLER_241_1808 ();
 FILLCELL_X32 FILLER_241_1840 ();
 FILLCELL_X32 FILLER_241_1872 ();
 FILLCELL_X32 FILLER_241_1904 ();
 FILLCELL_X32 FILLER_241_1936 ();
 FILLCELL_X32 FILLER_241_1968 ();
 FILLCELL_X32 FILLER_241_2000 ();
 FILLCELL_X32 FILLER_241_2032 ();
 FILLCELL_X32 FILLER_241_2064 ();
 FILLCELL_X32 FILLER_241_2096 ();
 FILLCELL_X32 FILLER_241_2128 ();
 FILLCELL_X32 FILLER_241_2160 ();
 FILLCELL_X32 FILLER_241_2192 ();
 FILLCELL_X32 FILLER_241_2224 ();
 FILLCELL_X32 FILLER_241_2256 ();
 FILLCELL_X32 FILLER_241_2288 ();
 FILLCELL_X32 FILLER_241_2320 ();
 FILLCELL_X32 FILLER_241_2352 ();
 FILLCELL_X32 FILLER_241_2384 ();
 FILLCELL_X16 FILLER_241_2416 ();
 FILLCELL_X4 FILLER_241_2432 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X32 FILLER_242_824 ();
 FILLCELL_X32 FILLER_242_856 ();
 FILLCELL_X32 FILLER_242_888 ();
 FILLCELL_X32 FILLER_242_920 ();
 FILLCELL_X32 FILLER_242_952 ();
 FILLCELL_X32 FILLER_242_984 ();
 FILLCELL_X32 FILLER_242_1016 ();
 FILLCELL_X32 FILLER_242_1048 ();
 FILLCELL_X32 FILLER_242_1080 ();
 FILLCELL_X32 FILLER_242_1112 ();
 FILLCELL_X32 FILLER_242_1144 ();
 FILLCELL_X32 FILLER_242_1176 ();
 FILLCELL_X32 FILLER_242_1208 ();
 FILLCELL_X32 FILLER_242_1240 ();
 FILLCELL_X32 FILLER_242_1272 ();
 FILLCELL_X32 FILLER_242_1304 ();
 FILLCELL_X32 FILLER_242_1336 ();
 FILLCELL_X32 FILLER_242_1368 ();
 FILLCELL_X32 FILLER_242_1400 ();
 FILLCELL_X32 FILLER_242_1432 ();
 FILLCELL_X32 FILLER_242_1464 ();
 FILLCELL_X32 FILLER_242_1496 ();
 FILLCELL_X32 FILLER_242_1528 ();
 FILLCELL_X32 FILLER_242_1560 ();
 FILLCELL_X32 FILLER_242_1592 ();
 FILLCELL_X32 FILLER_242_1624 ();
 FILLCELL_X32 FILLER_242_1656 ();
 FILLCELL_X32 FILLER_242_1688 ();
 FILLCELL_X32 FILLER_242_1720 ();
 FILLCELL_X32 FILLER_242_1752 ();
 FILLCELL_X32 FILLER_242_1784 ();
 FILLCELL_X32 FILLER_242_1816 ();
 FILLCELL_X32 FILLER_242_1848 ();
 FILLCELL_X8 FILLER_242_1880 ();
 FILLCELL_X4 FILLER_242_1888 ();
 FILLCELL_X2 FILLER_242_1892 ();
 FILLCELL_X32 FILLER_242_1895 ();
 FILLCELL_X32 FILLER_242_1927 ();
 FILLCELL_X32 FILLER_242_1959 ();
 FILLCELL_X32 FILLER_242_1991 ();
 FILLCELL_X32 FILLER_242_2023 ();
 FILLCELL_X32 FILLER_242_2055 ();
 FILLCELL_X32 FILLER_242_2087 ();
 FILLCELL_X32 FILLER_242_2119 ();
 FILLCELL_X32 FILLER_242_2151 ();
 FILLCELL_X32 FILLER_242_2183 ();
 FILLCELL_X32 FILLER_242_2215 ();
 FILLCELL_X32 FILLER_242_2247 ();
 FILLCELL_X32 FILLER_242_2279 ();
 FILLCELL_X32 FILLER_242_2311 ();
 FILLCELL_X32 FILLER_242_2343 ();
 FILLCELL_X32 FILLER_242_2375 ();
 FILLCELL_X16 FILLER_242_2407 ();
 FILLCELL_X8 FILLER_242_2423 ();
 FILLCELL_X4 FILLER_242_2431 ();
 FILLCELL_X1 FILLER_242_2435 ();
 FILLCELL_X32 FILLER_243_1 ();
 FILLCELL_X32 FILLER_243_33 ();
 FILLCELL_X32 FILLER_243_65 ();
 FILLCELL_X32 FILLER_243_97 ();
 FILLCELL_X32 FILLER_243_129 ();
 FILLCELL_X32 FILLER_243_161 ();
 FILLCELL_X32 FILLER_243_193 ();
 FILLCELL_X32 FILLER_243_225 ();
 FILLCELL_X32 FILLER_243_257 ();
 FILLCELL_X32 FILLER_243_289 ();
 FILLCELL_X32 FILLER_243_321 ();
 FILLCELL_X32 FILLER_243_353 ();
 FILLCELL_X32 FILLER_243_385 ();
 FILLCELL_X32 FILLER_243_417 ();
 FILLCELL_X32 FILLER_243_449 ();
 FILLCELL_X32 FILLER_243_481 ();
 FILLCELL_X32 FILLER_243_513 ();
 FILLCELL_X32 FILLER_243_545 ();
 FILLCELL_X32 FILLER_243_577 ();
 FILLCELL_X32 FILLER_243_609 ();
 FILLCELL_X32 FILLER_243_641 ();
 FILLCELL_X32 FILLER_243_673 ();
 FILLCELL_X32 FILLER_243_705 ();
 FILLCELL_X32 FILLER_243_737 ();
 FILLCELL_X32 FILLER_243_769 ();
 FILLCELL_X32 FILLER_243_801 ();
 FILLCELL_X32 FILLER_243_833 ();
 FILLCELL_X32 FILLER_243_865 ();
 FILLCELL_X32 FILLER_243_897 ();
 FILLCELL_X32 FILLER_243_929 ();
 FILLCELL_X32 FILLER_243_961 ();
 FILLCELL_X32 FILLER_243_993 ();
 FILLCELL_X32 FILLER_243_1025 ();
 FILLCELL_X32 FILLER_243_1057 ();
 FILLCELL_X32 FILLER_243_1089 ();
 FILLCELL_X32 FILLER_243_1121 ();
 FILLCELL_X32 FILLER_243_1153 ();
 FILLCELL_X32 FILLER_243_1185 ();
 FILLCELL_X32 FILLER_243_1217 ();
 FILLCELL_X8 FILLER_243_1249 ();
 FILLCELL_X4 FILLER_243_1257 ();
 FILLCELL_X2 FILLER_243_1261 ();
 FILLCELL_X32 FILLER_243_1264 ();
 FILLCELL_X32 FILLER_243_1296 ();
 FILLCELL_X32 FILLER_243_1328 ();
 FILLCELL_X32 FILLER_243_1360 ();
 FILLCELL_X32 FILLER_243_1392 ();
 FILLCELL_X32 FILLER_243_1424 ();
 FILLCELL_X32 FILLER_243_1456 ();
 FILLCELL_X32 FILLER_243_1488 ();
 FILLCELL_X32 FILLER_243_1520 ();
 FILLCELL_X32 FILLER_243_1552 ();
 FILLCELL_X32 FILLER_243_1584 ();
 FILLCELL_X32 FILLER_243_1616 ();
 FILLCELL_X32 FILLER_243_1648 ();
 FILLCELL_X32 FILLER_243_1680 ();
 FILLCELL_X32 FILLER_243_1712 ();
 FILLCELL_X32 FILLER_243_1744 ();
 FILLCELL_X32 FILLER_243_1776 ();
 FILLCELL_X32 FILLER_243_1808 ();
 FILLCELL_X32 FILLER_243_1840 ();
 FILLCELL_X32 FILLER_243_1872 ();
 FILLCELL_X32 FILLER_243_1904 ();
 FILLCELL_X32 FILLER_243_1936 ();
 FILLCELL_X32 FILLER_243_1968 ();
 FILLCELL_X32 FILLER_243_2000 ();
 FILLCELL_X32 FILLER_243_2032 ();
 FILLCELL_X32 FILLER_243_2064 ();
 FILLCELL_X32 FILLER_243_2096 ();
 FILLCELL_X32 FILLER_243_2128 ();
 FILLCELL_X32 FILLER_243_2160 ();
 FILLCELL_X32 FILLER_243_2192 ();
 FILLCELL_X32 FILLER_243_2224 ();
 FILLCELL_X32 FILLER_243_2256 ();
 FILLCELL_X32 FILLER_243_2288 ();
 FILLCELL_X32 FILLER_243_2320 ();
 FILLCELL_X32 FILLER_243_2352 ();
 FILLCELL_X32 FILLER_243_2384 ();
 FILLCELL_X16 FILLER_243_2416 ();
 FILLCELL_X4 FILLER_243_2432 ();
 FILLCELL_X32 FILLER_244_1 ();
 FILLCELL_X32 FILLER_244_33 ();
 FILLCELL_X32 FILLER_244_65 ();
 FILLCELL_X32 FILLER_244_97 ();
 FILLCELL_X32 FILLER_244_129 ();
 FILLCELL_X32 FILLER_244_161 ();
 FILLCELL_X32 FILLER_244_193 ();
 FILLCELL_X32 FILLER_244_225 ();
 FILLCELL_X32 FILLER_244_257 ();
 FILLCELL_X32 FILLER_244_289 ();
 FILLCELL_X32 FILLER_244_321 ();
 FILLCELL_X32 FILLER_244_353 ();
 FILLCELL_X32 FILLER_244_385 ();
 FILLCELL_X32 FILLER_244_417 ();
 FILLCELL_X32 FILLER_244_449 ();
 FILLCELL_X32 FILLER_244_481 ();
 FILLCELL_X32 FILLER_244_513 ();
 FILLCELL_X32 FILLER_244_545 ();
 FILLCELL_X32 FILLER_244_577 ();
 FILLCELL_X16 FILLER_244_609 ();
 FILLCELL_X4 FILLER_244_625 ();
 FILLCELL_X2 FILLER_244_629 ();
 FILLCELL_X32 FILLER_244_632 ();
 FILLCELL_X32 FILLER_244_664 ();
 FILLCELL_X32 FILLER_244_696 ();
 FILLCELL_X32 FILLER_244_728 ();
 FILLCELL_X32 FILLER_244_760 ();
 FILLCELL_X32 FILLER_244_792 ();
 FILLCELL_X32 FILLER_244_824 ();
 FILLCELL_X32 FILLER_244_856 ();
 FILLCELL_X32 FILLER_244_888 ();
 FILLCELL_X32 FILLER_244_920 ();
 FILLCELL_X32 FILLER_244_952 ();
 FILLCELL_X32 FILLER_244_984 ();
 FILLCELL_X32 FILLER_244_1016 ();
 FILLCELL_X32 FILLER_244_1048 ();
 FILLCELL_X32 FILLER_244_1080 ();
 FILLCELL_X32 FILLER_244_1112 ();
 FILLCELL_X32 FILLER_244_1144 ();
 FILLCELL_X32 FILLER_244_1176 ();
 FILLCELL_X32 FILLER_244_1208 ();
 FILLCELL_X32 FILLER_244_1240 ();
 FILLCELL_X32 FILLER_244_1272 ();
 FILLCELL_X32 FILLER_244_1304 ();
 FILLCELL_X32 FILLER_244_1336 ();
 FILLCELL_X32 FILLER_244_1368 ();
 FILLCELL_X32 FILLER_244_1400 ();
 FILLCELL_X32 FILLER_244_1432 ();
 FILLCELL_X32 FILLER_244_1464 ();
 FILLCELL_X32 FILLER_244_1496 ();
 FILLCELL_X32 FILLER_244_1528 ();
 FILLCELL_X32 FILLER_244_1560 ();
 FILLCELL_X32 FILLER_244_1592 ();
 FILLCELL_X32 FILLER_244_1624 ();
 FILLCELL_X32 FILLER_244_1656 ();
 FILLCELL_X32 FILLER_244_1688 ();
 FILLCELL_X32 FILLER_244_1720 ();
 FILLCELL_X32 FILLER_244_1752 ();
 FILLCELL_X32 FILLER_244_1784 ();
 FILLCELL_X32 FILLER_244_1816 ();
 FILLCELL_X32 FILLER_244_1848 ();
 FILLCELL_X8 FILLER_244_1880 ();
 FILLCELL_X4 FILLER_244_1888 ();
 FILLCELL_X2 FILLER_244_1892 ();
 FILLCELL_X32 FILLER_244_1895 ();
 FILLCELL_X32 FILLER_244_1927 ();
 FILLCELL_X32 FILLER_244_1959 ();
 FILLCELL_X32 FILLER_244_1991 ();
 FILLCELL_X32 FILLER_244_2023 ();
 FILLCELL_X32 FILLER_244_2055 ();
 FILLCELL_X32 FILLER_244_2087 ();
 FILLCELL_X32 FILLER_244_2119 ();
 FILLCELL_X32 FILLER_244_2151 ();
 FILLCELL_X32 FILLER_244_2183 ();
 FILLCELL_X32 FILLER_244_2215 ();
 FILLCELL_X32 FILLER_244_2247 ();
 FILLCELL_X32 FILLER_244_2279 ();
 FILLCELL_X32 FILLER_244_2311 ();
 FILLCELL_X32 FILLER_244_2343 ();
 FILLCELL_X32 FILLER_244_2375 ();
 FILLCELL_X16 FILLER_244_2407 ();
 FILLCELL_X8 FILLER_244_2423 ();
 FILLCELL_X4 FILLER_244_2431 ();
 FILLCELL_X1 FILLER_244_2435 ();
 FILLCELL_X32 FILLER_245_1 ();
 FILLCELL_X32 FILLER_245_33 ();
 FILLCELL_X32 FILLER_245_65 ();
 FILLCELL_X32 FILLER_245_97 ();
 FILLCELL_X32 FILLER_245_129 ();
 FILLCELL_X32 FILLER_245_161 ();
 FILLCELL_X32 FILLER_245_193 ();
 FILLCELL_X32 FILLER_245_225 ();
 FILLCELL_X32 FILLER_245_257 ();
 FILLCELL_X32 FILLER_245_289 ();
 FILLCELL_X32 FILLER_245_321 ();
 FILLCELL_X32 FILLER_245_353 ();
 FILLCELL_X32 FILLER_245_385 ();
 FILLCELL_X32 FILLER_245_417 ();
 FILLCELL_X32 FILLER_245_449 ();
 FILLCELL_X32 FILLER_245_481 ();
 FILLCELL_X32 FILLER_245_513 ();
 FILLCELL_X32 FILLER_245_545 ();
 FILLCELL_X32 FILLER_245_577 ();
 FILLCELL_X32 FILLER_245_609 ();
 FILLCELL_X32 FILLER_245_641 ();
 FILLCELL_X32 FILLER_245_673 ();
 FILLCELL_X32 FILLER_245_705 ();
 FILLCELL_X32 FILLER_245_737 ();
 FILLCELL_X32 FILLER_245_769 ();
 FILLCELL_X32 FILLER_245_801 ();
 FILLCELL_X32 FILLER_245_833 ();
 FILLCELL_X32 FILLER_245_865 ();
 FILLCELL_X32 FILLER_245_897 ();
 FILLCELL_X32 FILLER_245_929 ();
 FILLCELL_X32 FILLER_245_961 ();
 FILLCELL_X32 FILLER_245_993 ();
 FILLCELL_X32 FILLER_245_1025 ();
 FILLCELL_X32 FILLER_245_1057 ();
 FILLCELL_X32 FILLER_245_1089 ();
 FILLCELL_X32 FILLER_245_1121 ();
 FILLCELL_X32 FILLER_245_1153 ();
 FILLCELL_X32 FILLER_245_1185 ();
 FILLCELL_X32 FILLER_245_1217 ();
 FILLCELL_X8 FILLER_245_1249 ();
 FILLCELL_X4 FILLER_245_1257 ();
 FILLCELL_X2 FILLER_245_1261 ();
 FILLCELL_X32 FILLER_245_1264 ();
 FILLCELL_X32 FILLER_245_1296 ();
 FILLCELL_X32 FILLER_245_1328 ();
 FILLCELL_X32 FILLER_245_1360 ();
 FILLCELL_X32 FILLER_245_1392 ();
 FILLCELL_X32 FILLER_245_1424 ();
 FILLCELL_X32 FILLER_245_1456 ();
 FILLCELL_X32 FILLER_245_1488 ();
 FILLCELL_X32 FILLER_245_1520 ();
 FILLCELL_X32 FILLER_245_1552 ();
 FILLCELL_X32 FILLER_245_1584 ();
 FILLCELL_X32 FILLER_245_1616 ();
 FILLCELL_X32 FILLER_245_1648 ();
 FILLCELL_X32 FILLER_245_1680 ();
 FILLCELL_X32 FILLER_245_1712 ();
 FILLCELL_X32 FILLER_245_1744 ();
 FILLCELL_X32 FILLER_245_1776 ();
 FILLCELL_X32 FILLER_245_1808 ();
 FILLCELL_X32 FILLER_245_1840 ();
 FILLCELL_X32 FILLER_245_1872 ();
 FILLCELL_X32 FILLER_245_1904 ();
 FILLCELL_X32 FILLER_245_1936 ();
 FILLCELL_X32 FILLER_245_1968 ();
 FILLCELL_X32 FILLER_245_2000 ();
 FILLCELL_X32 FILLER_245_2032 ();
 FILLCELL_X32 FILLER_245_2064 ();
 FILLCELL_X32 FILLER_245_2096 ();
 FILLCELL_X32 FILLER_245_2128 ();
 FILLCELL_X32 FILLER_245_2160 ();
 FILLCELL_X32 FILLER_245_2192 ();
 FILLCELL_X32 FILLER_245_2224 ();
 FILLCELL_X32 FILLER_245_2256 ();
 FILLCELL_X32 FILLER_245_2288 ();
 FILLCELL_X32 FILLER_245_2320 ();
 FILLCELL_X32 FILLER_245_2352 ();
 FILLCELL_X32 FILLER_245_2384 ();
 FILLCELL_X16 FILLER_245_2416 ();
 FILLCELL_X4 FILLER_245_2432 ();
 FILLCELL_X32 FILLER_246_1 ();
 FILLCELL_X32 FILLER_246_33 ();
 FILLCELL_X32 FILLER_246_65 ();
 FILLCELL_X32 FILLER_246_97 ();
 FILLCELL_X32 FILLER_246_129 ();
 FILLCELL_X32 FILLER_246_161 ();
 FILLCELL_X32 FILLER_246_193 ();
 FILLCELL_X32 FILLER_246_225 ();
 FILLCELL_X32 FILLER_246_257 ();
 FILLCELL_X32 FILLER_246_289 ();
 FILLCELL_X32 FILLER_246_321 ();
 FILLCELL_X32 FILLER_246_353 ();
 FILLCELL_X32 FILLER_246_385 ();
 FILLCELL_X32 FILLER_246_417 ();
 FILLCELL_X32 FILLER_246_449 ();
 FILLCELL_X32 FILLER_246_481 ();
 FILLCELL_X32 FILLER_246_513 ();
 FILLCELL_X32 FILLER_246_545 ();
 FILLCELL_X32 FILLER_246_577 ();
 FILLCELL_X16 FILLER_246_609 ();
 FILLCELL_X4 FILLER_246_625 ();
 FILLCELL_X2 FILLER_246_629 ();
 FILLCELL_X32 FILLER_246_632 ();
 FILLCELL_X32 FILLER_246_664 ();
 FILLCELL_X32 FILLER_246_696 ();
 FILLCELL_X32 FILLER_246_728 ();
 FILLCELL_X32 FILLER_246_760 ();
 FILLCELL_X32 FILLER_246_792 ();
 FILLCELL_X32 FILLER_246_824 ();
 FILLCELL_X32 FILLER_246_856 ();
 FILLCELL_X32 FILLER_246_888 ();
 FILLCELL_X32 FILLER_246_920 ();
 FILLCELL_X32 FILLER_246_952 ();
 FILLCELL_X32 FILLER_246_984 ();
 FILLCELL_X32 FILLER_246_1016 ();
 FILLCELL_X32 FILLER_246_1048 ();
 FILLCELL_X32 FILLER_246_1080 ();
 FILLCELL_X32 FILLER_246_1112 ();
 FILLCELL_X32 FILLER_246_1144 ();
 FILLCELL_X32 FILLER_246_1176 ();
 FILLCELL_X32 FILLER_246_1208 ();
 FILLCELL_X32 FILLER_246_1240 ();
 FILLCELL_X32 FILLER_246_1272 ();
 FILLCELL_X32 FILLER_246_1304 ();
 FILLCELL_X32 FILLER_246_1336 ();
 FILLCELL_X32 FILLER_246_1368 ();
 FILLCELL_X32 FILLER_246_1400 ();
 FILLCELL_X32 FILLER_246_1432 ();
 FILLCELL_X32 FILLER_246_1464 ();
 FILLCELL_X32 FILLER_246_1496 ();
 FILLCELL_X32 FILLER_246_1528 ();
 FILLCELL_X32 FILLER_246_1560 ();
 FILLCELL_X32 FILLER_246_1592 ();
 FILLCELL_X32 FILLER_246_1624 ();
 FILLCELL_X32 FILLER_246_1656 ();
 FILLCELL_X32 FILLER_246_1688 ();
 FILLCELL_X32 FILLER_246_1720 ();
 FILLCELL_X32 FILLER_246_1752 ();
 FILLCELL_X32 FILLER_246_1784 ();
 FILLCELL_X32 FILLER_246_1816 ();
 FILLCELL_X32 FILLER_246_1848 ();
 FILLCELL_X8 FILLER_246_1880 ();
 FILLCELL_X4 FILLER_246_1888 ();
 FILLCELL_X2 FILLER_246_1892 ();
 FILLCELL_X32 FILLER_246_1895 ();
 FILLCELL_X32 FILLER_246_1927 ();
 FILLCELL_X32 FILLER_246_1959 ();
 FILLCELL_X32 FILLER_246_1991 ();
 FILLCELL_X32 FILLER_246_2023 ();
 FILLCELL_X32 FILLER_246_2055 ();
 FILLCELL_X32 FILLER_246_2087 ();
 FILLCELL_X32 FILLER_246_2119 ();
 FILLCELL_X32 FILLER_246_2151 ();
 FILLCELL_X32 FILLER_246_2183 ();
 FILLCELL_X32 FILLER_246_2215 ();
 FILLCELL_X32 FILLER_246_2247 ();
 FILLCELL_X32 FILLER_246_2279 ();
 FILLCELL_X32 FILLER_246_2311 ();
 FILLCELL_X32 FILLER_246_2343 ();
 FILLCELL_X32 FILLER_246_2375 ();
 FILLCELL_X16 FILLER_246_2407 ();
 FILLCELL_X8 FILLER_246_2423 ();
 FILLCELL_X4 FILLER_246_2431 ();
 FILLCELL_X1 FILLER_246_2435 ();
 FILLCELL_X32 FILLER_247_1 ();
 FILLCELL_X32 FILLER_247_33 ();
 FILLCELL_X32 FILLER_247_65 ();
 FILLCELL_X32 FILLER_247_97 ();
 FILLCELL_X32 FILLER_247_129 ();
 FILLCELL_X32 FILLER_247_161 ();
 FILLCELL_X32 FILLER_247_193 ();
 FILLCELL_X32 FILLER_247_225 ();
 FILLCELL_X32 FILLER_247_257 ();
 FILLCELL_X32 FILLER_247_289 ();
 FILLCELL_X32 FILLER_247_321 ();
 FILLCELL_X32 FILLER_247_353 ();
 FILLCELL_X32 FILLER_247_385 ();
 FILLCELL_X32 FILLER_247_417 ();
 FILLCELL_X32 FILLER_247_449 ();
 FILLCELL_X32 FILLER_247_481 ();
 FILLCELL_X32 FILLER_247_513 ();
 FILLCELL_X32 FILLER_247_545 ();
 FILLCELL_X32 FILLER_247_577 ();
 FILLCELL_X32 FILLER_247_609 ();
 FILLCELL_X32 FILLER_247_641 ();
 FILLCELL_X32 FILLER_247_673 ();
 FILLCELL_X32 FILLER_247_705 ();
 FILLCELL_X32 FILLER_247_737 ();
 FILLCELL_X32 FILLER_247_769 ();
 FILLCELL_X32 FILLER_247_801 ();
 FILLCELL_X32 FILLER_247_833 ();
 FILLCELL_X32 FILLER_247_865 ();
 FILLCELL_X32 FILLER_247_897 ();
 FILLCELL_X32 FILLER_247_929 ();
 FILLCELL_X32 FILLER_247_961 ();
 FILLCELL_X32 FILLER_247_993 ();
 FILLCELL_X32 FILLER_247_1025 ();
 FILLCELL_X32 FILLER_247_1057 ();
 FILLCELL_X32 FILLER_247_1089 ();
 FILLCELL_X32 FILLER_247_1121 ();
 FILLCELL_X32 FILLER_247_1153 ();
 FILLCELL_X32 FILLER_247_1185 ();
 FILLCELL_X32 FILLER_247_1217 ();
 FILLCELL_X8 FILLER_247_1249 ();
 FILLCELL_X4 FILLER_247_1257 ();
 FILLCELL_X2 FILLER_247_1261 ();
 FILLCELL_X32 FILLER_247_1264 ();
 FILLCELL_X32 FILLER_247_1296 ();
 FILLCELL_X32 FILLER_247_1328 ();
 FILLCELL_X32 FILLER_247_1360 ();
 FILLCELL_X32 FILLER_247_1392 ();
 FILLCELL_X32 FILLER_247_1424 ();
 FILLCELL_X32 FILLER_247_1456 ();
 FILLCELL_X32 FILLER_247_1488 ();
 FILLCELL_X32 FILLER_247_1520 ();
 FILLCELL_X32 FILLER_247_1552 ();
 FILLCELL_X32 FILLER_247_1584 ();
 FILLCELL_X32 FILLER_247_1616 ();
 FILLCELL_X32 FILLER_247_1648 ();
 FILLCELL_X32 FILLER_247_1680 ();
 FILLCELL_X32 FILLER_247_1712 ();
 FILLCELL_X32 FILLER_247_1744 ();
 FILLCELL_X32 FILLER_247_1776 ();
 FILLCELL_X32 FILLER_247_1808 ();
 FILLCELL_X32 FILLER_247_1840 ();
 FILLCELL_X32 FILLER_247_1872 ();
 FILLCELL_X32 FILLER_247_1904 ();
 FILLCELL_X32 FILLER_247_1936 ();
 FILLCELL_X32 FILLER_247_1968 ();
 FILLCELL_X32 FILLER_247_2000 ();
 FILLCELL_X32 FILLER_247_2032 ();
 FILLCELL_X32 FILLER_247_2064 ();
 FILLCELL_X32 FILLER_247_2096 ();
 FILLCELL_X32 FILLER_247_2128 ();
 FILLCELL_X32 FILLER_247_2160 ();
 FILLCELL_X32 FILLER_247_2192 ();
 FILLCELL_X32 FILLER_247_2224 ();
 FILLCELL_X32 FILLER_247_2256 ();
 FILLCELL_X32 FILLER_247_2288 ();
 FILLCELL_X32 FILLER_247_2320 ();
 FILLCELL_X32 FILLER_247_2352 ();
 FILLCELL_X32 FILLER_247_2384 ();
 FILLCELL_X16 FILLER_247_2416 ();
 FILLCELL_X4 FILLER_247_2432 ();
 FILLCELL_X32 FILLER_248_1 ();
 FILLCELL_X32 FILLER_248_33 ();
 FILLCELL_X32 FILLER_248_65 ();
 FILLCELL_X32 FILLER_248_97 ();
 FILLCELL_X32 FILLER_248_129 ();
 FILLCELL_X32 FILLER_248_161 ();
 FILLCELL_X32 FILLER_248_193 ();
 FILLCELL_X32 FILLER_248_225 ();
 FILLCELL_X32 FILLER_248_257 ();
 FILLCELL_X32 FILLER_248_289 ();
 FILLCELL_X32 FILLER_248_321 ();
 FILLCELL_X32 FILLER_248_353 ();
 FILLCELL_X32 FILLER_248_385 ();
 FILLCELL_X32 FILLER_248_417 ();
 FILLCELL_X32 FILLER_248_449 ();
 FILLCELL_X32 FILLER_248_481 ();
 FILLCELL_X32 FILLER_248_513 ();
 FILLCELL_X32 FILLER_248_545 ();
 FILLCELL_X32 FILLER_248_577 ();
 FILLCELL_X16 FILLER_248_609 ();
 FILLCELL_X4 FILLER_248_625 ();
 FILLCELL_X2 FILLER_248_629 ();
 FILLCELL_X32 FILLER_248_632 ();
 FILLCELL_X32 FILLER_248_664 ();
 FILLCELL_X32 FILLER_248_696 ();
 FILLCELL_X32 FILLER_248_728 ();
 FILLCELL_X32 FILLER_248_760 ();
 FILLCELL_X32 FILLER_248_792 ();
 FILLCELL_X32 FILLER_248_824 ();
 FILLCELL_X32 FILLER_248_856 ();
 FILLCELL_X32 FILLER_248_888 ();
 FILLCELL_X32 FILLER_248_920 ();
 FILLCELL_X32 FILLER_248_952 ();
 FILLCELL_X32 FILLER_248_984 ();
 FILLCELL_X32 FILLER_248_1016 ();
 FILLCELL_X32 FILLER_248_1048 ();
 FILLCELL_X32 FILLER_248_1080 ();
 FILLCELL_X32 FILLER_248_1112 ();
 FILLCELL_X32 FILLER_248_1144 ();
 FILLCELL_X32 FILLER_248_1176 ();
 FILLCELL_X32 FILLER_248_1208 ();
 FILLCELL_X32 FILLER_248_1240 ();
 FILLCELL_X32 FILLER_248_1272 ();
 FILLCELL_X32 FILLER_248_1304 ();
 FILLCELL_X32 FILLER_248_1336 ();
 FILLCELL_X32 FILLER_248_1368 ();
 FILLCELL_X32 FILLER_248_1400 ();
 FILLCELL_X32 FILLER_248_1432 ();
 FILLCELL_X32 FILLER_248_1464 ();
 FILLCELL_X32 FILLER_248_1496 ();
 FILLCELL_X32 FILLER_248_1528 ();
 FILLCELL_X32 FILLER_248_1560 ();
 FILLCELL_X32 FILLER_248_1592 ();
 FILLCELL_X32 FILLER_248_1624 ();
 FILLCELL_X32 FILLER_248_1656 ();
 FILLCELL_X32 FILLER_248_1688 ();
 FILLCELL_X32 FILLER_248_1720 ();
 FILLCELL_X32 FILLER_248_1752 ();
 FILLCELL_X32 FILLER_248_1784 ();
 FILLCELL_X32 FILLER_248_1816 ();
 FILLCELL_X32 FILLER_248_1848 ();
 FILLCELL_X8 FILLER_248_1880 ();
 FILLCELL_X4 FILLER_248_1888 ();
 FILLCELL_X2 FILLER_248_1892 ();
 FILLCELL_X32 FILLER_248_1895 ();
 FILLCELL_X32 FILLER_248_1927 ();
 FILLCELL_X32 FILLER_248_1959 ();
 FILLCELL_X32 FILLER_248_1991 ();
 FILLCELL_X32 FILLER_248_2023 ();
 FILLCELL_X32 FILLER_248_2055 ();
 FILLCELL_X32 FILLER_248_2087 ();
 FILLCELL_X32 FILLER_248_2119 ();
 FILLCELL_X32 FILLER_248_2151 ();
 FILLCELL_X32 FILLER_248_2183 ();
 FILLCELL_X32 FILLER_248_2215 ();
 FILLCELL_X32 FILLER_248_2247 ();
 FILLCELL_X32 FILLER_248_2279 ();
 FILLCELL_X32 FILLER_248_2311 ();
 FILLCELL_X32 FILLER_248_2343 ();
 FILLCELL_X32 FILLER_248_2375 ();
 FILLCELL_X16 FILLER_248_2407 ();
 FILLCELL_X8 FILLER_248_2423 ();
 FILLCELL_X4 FILLER_248_2431 ();
 FILLCELL_X1 FILLER_248_2435 ();
 FILLCELL_X32 FILLER_249_1 ();
 FILLCELL_X32 FILLER_249_33 ();
 FILLCELL_X32 FILLER_249_65 ();
 FILLCELL_X32 FILLER_249_97 ();
 FILLCELL_X32 FILLER_249_129 ();
 FILLCELL_X32 FILLER_249_161 ();
 FILLCELL_X32 FILLER_249_193 ();
 FILLCELL_X32 FILLER_249_225 ();
 FILLCELL_X32 FILLER_249_257 ();
 FILLCELL_X32 FILLER_249_289 ();
 FILLCELL_X32 FILLER_249_321 ();
 FILLCELL_X32 FILLER_249_353 ();
 FILLCELL_X32 FILLER_249_385 ();
 FILLCELL_X32 FILLER_249_417 ();
 FILLCELL_X32 FILLER_249_449 ();
 FILLCELL_X32 FILLER_249_481 ();
 FILLCELL_X32 FILLER_249_513 ();
 FILLCELL_X32 FILLER_249_545 ();
 FILLCELL_X32 FILLER_249_577 ();
 FILLCELL_X32 FILLER_249_609 ();
 FILLCELL_X32 FILLER_249_641 ();
 FILLCELL_X32 FILLER_249_673 ();
 FILLCELL_X32 FILLER_249_705 ();
 FILLCELL_X32 FILLER_249_737 ();
 FILLCELL_X32 FILLER_249_769 ();
 FILLCELL_X32 FILLER_249_801 ();
 FILLCELL_X32 FILLER_249_833 ();
 FILLCELL_X32 FILLER_249_865 ();
 FILLCELL_X32 FILLER_249_897 ();
 FILLCELL_X32 FILLER_249_929 ();
 FILLCELL_X32 FILLER_249_961 ();
 FILLCELL_X32 FILLER_249_993 ();
 FILLCELL_X32 FILLER_249_1025 ();
 FILLCELL_X32 FILLER_249_1057 ();
 FILLCELL_X32 FILLER_249_1089 ();
 FILLCELL_X32 FILLER_249_1121 ();
 FILLCELL_X32 FILLER_249_1153 ();
 FILLCELL_X32 FILLER_249_1185 ();
 FILLCELL_X32 FILLER_249_1217 ();
 FILLCELL_X8 FILLER_249_1249 ();
 FILLCELL_X4 FILLER_249_1257 ();
 FILLCELL_X2 FILLER_249_1261 ();
 FILLCELL_X32 FILLER_249_1264 ();
 FILLCELL_X32 FILLER_249_1296 ();
 FILLCELL_X32 FILLER_249_1328 ();
 FILLCELL_X32 FILLER_249_1360 ();
 FILLCELL_X32 FILLER_249_1392 ();
 FILLCELL_X32 FILLER_249_1424 ();
 FILLCELL_X32 FILLER_249_1456 ();
 FILLCELL_X32 FILLER_249_1488 ();
 FILLCELL_X32 FILLER_249_1520 ();
 FILLCELL_X32 FILLER_249_1552 ();
 FILLCELL_X32 FILLER_249_1584 ();
 FILLCELL_X32 FILLER_249_1616 ();
 FILLCELL_X32 FILLER_249_1648 ();
 FILLCELL_X32 FILLER_249_1680 ();
 FILLCELL_X32 FILLER_249_1712 ();
 FILLCELL_X32 FILLER_249_1744 ();
 FILLCELL_X32 FILLER_249_1776 ();
 FILLCELL_X32 FILLER_249_1808 ();
 FILLCELL_X32 FILLER_249_1840 ();
 FILLCELL_X32 FILLER_249_1872 ();
 FILLCELL_X32 FILLER_249_1904 ();
 FILLCELL_X32 FILLER_249_1936 ();
 FILLCELL_X32 FILLER_249_1968 ();
 FILLCELL_X32 FILLER_249_2000 ();
 FILLCELL_X32 FILLER_249_2032 ();
 FILLCELL_X32 FILLER_249_2064 ();
 FILLCELL_X32 FILLER_249_2096 ();
 FILLCELL_X32 FILLER_249_2128 ();
 FILLCELL_X32 FILLER_249_2160 ();
 FILLCELL_X32 FILLER_249_2192 ();
 FILLCELL_X32 FILLER_249_2224 ();
 FILLCELL_X32 FILLER_249_2256 ();
 FILLCELL_X32 FILLER_249_2288 ();
 FILLCELL_X32 FILLER_249_2320 ();
 FILLCELL_X32 FILLER_249_2352 ();
 FILLCELL_X32 FILLER_249_2384 ();
 FILLCELL_X16 FILLER_249_2416 ();
 FILLCELL_X4 FILLER_249_2432 ();
 FILLCELL_X32 FILLER_250_1 ();
 FILLCELL_X32 FILLER_250_33 ();
 FILLCELL_X32 FILLER_250_65 ();
 FILLCELL_X32 FILLER_250_97 ();
 FILLCELL_X32 FILLER_250_129 ();
 FILLCELL_X32 FILLER_250_161 ();
 FILLCELL_X32 FILLER_250_193 ();
 FILLCELL_X32 FILLER_250_225 ();
 FILLCELL_X32 FILLER_250_257 ();
 FILLCELL_X32 FILLER_250_289 ();
 FILLCELL_X32 FILLER_250_321 ();
 FILLCELL_X32 FILLER_250_353 ();
 FILLCELL_X32 FILLER_250_385 ();
 FILLCELL_X32 FILLER_250_417 ();
 FILLCELL_X32 FILLER_250_449 ();
 FILLCELL_X32 FILLER_250_481 ();
 FILLCELL_X32 FILLER_250_513 ();
 FILLCELL_X32 FILLER_250_545 ();
 FILLCELL_X32 FILLER_250_577 ();
 FILLCELL_X16 FILLER_250_609 ();
 FILLCELL_X4 FILLER_250_625 ();
 FILLCELL_X2 FILLER_250_629 ();
 FILLCELL_X32 FILLER_250_632 ();
 FILLCELL_X32 FILLER_250_664 ();
 FILLCELL_X32 FILLER_250_696 ();
 FILLCELL_X32 FILLER_250_728 ();
 FILLCELL_X32 FILLER_250_760 ();
 FILLCELL_X32 FILLER_250_792 ();
 FILLCELL_X32 FILLER_250_824 ();
 FILLCELL_X32 FILLER_250_856 ();
 FILLCELL_X32 FILLER_250_888 ();
 FILLCELL_X32 FILLER_250_920 ();
 FILLCELL_X32 FILLER_250_952 ();
 FILLCELL_X32 FILLER_250_984 ();
 FILLCELL_X32 FILLER_250_1016 ();
 FILLCELL_X32 FILLER_250_1048 ();
 FILLCELL_X32 FILLER_250_1080 ();
 FILLCELL_X32 FILLER_250_1112 ();
 FILLCELL_X32 FILLER_250_1144 ();
 FILLCELL_X32 FILLER_250_1176 ();
 FILLCELL_X32 FILLER_250_1208 ();
 FILLCELL_X32 FILLER_250_1240 ();
 FILLCELL_X32 FILLER_250_1272 ();
 FILLCELL_X32 FILLER_250_1304 ();
 FILLCELL_X32 FILLER_250_1336 ();
 FILLCELL_X32 FILLER_250_1368 ();
 FILLCELL_X32 FILLER_250_1400 ();
 FILLCELL_X32 FILLER_250_1432 ();
 FILLCELL_X32 FILLER_250_1464 ();
 FILLCELL_X32 FILLER_250_1496 ();
 FILLCELL_X32 FILLER_250_1528 ();
 FILLCELL_X32 FILLER_250_1560 ();
 FILLCELL_X32 FILLER_250_1592 ();
 FILLCELL_X32 FILLER_250_1624 ();
 FILLCELL_X32 FILLER_250_1656 ();
 FILLCELL_X32 FILLER_250_1688 ();
 FILLCELL_X32 FILLER_250_1720 ();
 FILLCELL_X32 FILLER_250_1752 ();
 FILLCELL_X32 FILLER_250_1784 ();
 FILLCELL_X32 FILLER_250_1816 ();
 FILLCELL_X32 FILLER_250_1848 ();
 FILLCELL_X8 FILLER_250_1880 ();
 FILLCELL_X4 FILLER_250_1888 ();
 FILLCELL_X2 FILLER_250_1892 ();
 FILLCELL_X32 FILLER_250_1895 ();
 FILLCELL_X32 FILLER_250_1927 ();
 FILLCELL_X32 FILLER_250_1959 ();
 FILLCELL_X32 FILLER_250_1991 ();
 FILLCELL_X32 FILLER_250_2023 ();
 FILLCELL_X32 FILLER_250_2055 ();
 FILLCELL_X32 FILLER_250_2087 ();
 FILLCELL_X32 FILLER_250_2119 ();
 FILLCELL_X32 FILLER_250_2151 ();
 FILLCELL_X32 FILLER_250_2183 ();
 FILLCELL_X32 FILLER_250_2215 ();
 FILLCELL_X32 FILLER_250_2247 ();
 FILLCELL_X32 FILLER_250_2279 ();
 FILLCELL_X32 FILLER_250_2311 ();
 FILLCELL_X32 FILLER_250_2343 ();
 FILLCELL_X32 FILLER_250_2375 ();
 FILLCELL_X16 FILLER_250_2407 ();
 FILLCELL_X8 FILLER_250_2423 ();
 FILLCELL_X4 FILLER_250_2431 ();
 FILLCELL_X1 FILLER_250_2435 ();
 FILLCELL_X32 FILLER_251_1 ();
 FILLCELL_X32 FILLER_251_33 ();
 FILLCELL_X32 FILLER_251_65 ();
 FILLCELL_X32 FILLER_251_97 ();
 FILLCELL_X32 FILLER_251_129 ();
 FILLCELL_X32 FILLER_251_161 ();
 FILLCELL_X32 FILLER_251_193 ();
 FILLCELL_X32 FILLER_251_225 ();
 FILLCELL_X32 FILLER_251_257 ();
 FILLCELL_X32 FILLER_251_289 ();
 FILLCELL_X32 FILLER_251_321 ();
 FILLCELL_X32 FILLER_251_353 ();
 FILLCELL_X32 FILLER_251_385 ();
 FILLCELL_X32 FILLER_251_417 ();
 FILLCELL_X32 FILLER_251_449 ();
 FILLCELL_X32 FILLER_251_481 ();
 FILLCELL_X32 FILLER_251_513 ();
 FILLCELL_X32 FILLER_251_545 ();
 FILLCELL_X32 FILLER_251_577 ();
 FILLCELL_X32 FILLER_251_609 ();
 FILLCELL_X32 FILLER_251_641 ();
 FILLCELL_X32 FILLER_251_673 ();
 FILLCELL_X32 FILLER_251_705 ();
 FILLCELL_X32 FILLER_251_737 ();
 FILLCELL_X32 FILLER_251_769 ();
 FILLCELL_X32 FILLER_251_801 ();
 FILLCELL_X32 FILLER_251_833 ();
 FILLCELL_X32 FILLER_251_865 ();
 FILLCELL_X32 FILLER_251_897 ();
 FILLCELL_X32 FILLER_251_929 ();
 FILLCELL_X32 FILLER_251_961 ();
 FILLCELL_X32 FILLER_251_993 ();
 FILLCELL_X32 FILLER_251_1025 ();
 FILLCELL_X32 FILLER_251_1057 ();
 FILLCELL_X32 FILLER_251_1089 ();
 FILLCELL_X32 FILLER_251_1121 ();
 FILLCELL_X32 FILLER_251_1153 ();
 FILLCELL_X32 FILLER_251_1185 ();
 FILLCELL_X32 FILLER_251_1217 ();
 FILLCELL_X8 FILLER_251_1249 ();
 FILLCELL_X4 FILLER_251_1257 ();
 FILLCELL_X2 FILLER_251_1261 ();
 FILLCELL_X32 FILLER_251_1264 ();
 FILLCELL_X32 FILLER_251_1296 ();
 FILLCELL_X32 FILLER_251_1328 ();
 FILLCELL_X32 FILLER_251_1360 ();
 FILLCELL_X32 FILLER_251_1392 ();
 FILLCELL_X32 FILLER_251_1424 ();
 FILLCELL_X32 FILLER_251_1456 ();
 FILLCELL_X32 FILLER_251_1488 ();
 FILLCELL_X32 FILLER_251_1520 ();
 FILLCELL_X32 FILLER_251_1552 ();
 FILLCELL_X32 FILLER_251_1584 ();
 FILLCELL_X32 FILLER_251_1616 ();
 FILLCELL_X32 FILLER_251_1648 ();
 FILLCELL_X32 FILLER_251_1680 ();
 FILLCELL_X32 FILLER_251_1712 ();
 FILLCELL_X32 FILLER_251_1744 ();
 FILLCELL_X32 FILLER_251_1776 ();
 FILLCELL_X32 FILLER_251_1808 ();
 FILLCELL_X32 FILLER_251_1840 ();
 FILLCELL_X32 FILLER_251_1872 ();
 FILLCELL_X32 FILLER_251_1904 ();
 FILLCELL_X32 FILLER_251_1936 ();
 FILLCELL_X32 FILLER_251_1968 ();
 FILLCELL_X32 FILLER_251_2000 ();
 FILLCELL_X32 FILLER_251_2032 ();
 FILLCELL_X32 FILLER_251_2064 ();
 FILLCELL_X32 FILLER_251_2096 ();
 FILLCELL_X32 FILLER_251_2128 ();
 FILLCELL_X32 FILLER_251_2160 ();
 FILLCELL_X32 FILLER_251_2192 ();
 FILLCELL_X32 FILLER_251_2224 ();
 FILLCELL_X32 FILLER_251_2256 ();
 FILLCELL_X32 FILLER_251_2288 ();
 FILLCELL_X32 FILLER_251_2320 ();
 FILLCELL_X32 FILLER_251_2352 ();
 FILLCELL_X32 FILLER_251_2384 ();
 FILLCELL_X16 FILLER_251_2416 ();
 FILLCELL_X4 FILLER_251_2432 ();
 FILLCELL_X32 FILLER_252_1 ();
 FILLCELL_X32 FILLER_252_33 ();
 FILLCELL_X32 FILLER_252_65 ();
 FILLCELL_X32 FILLER_252_97 ();
 FILLCELL_X32 FILLER_252_129 ();
 FILLCELL_X32 FILLER_252_161 ();
 FILLCELL_X32 FILLER_252_193 ();
 FILLCELL_X32 FILLER_252_225 ();
 FILLCELL_X32 FILLER_252_257 ();
 FILLCELL_X32 FILLER_252_289 ();
 FILLCELL_X32 FILLER_252_321 ();
 FILLCELL_X32 FILLER_252_353 ();
 FILLCELL_X32 FILLER_252_385 ();
 FILLCELL_X32 FILLER_252_417 ();
 FILLCELL_X32 FILLER_252_449 ();
 FILLCELL_X32 FILLER_252_481 ();
 FILLCELL_X32 FILLER_252_513 ();
 FILLCELL_X32 FILLER_252_545 ();
 FILLCELL_X32 FILLER_252_577 ();
 FILLCELL_X16 FILLER_252_609 ();
 FILLCELL_X4 FILLER_252_625 ();
 FILLCELL_X2 FILLER_252_629 ();
 FILLCELL_X32 FILLER_252_632 ();
 FILLCELL_X32 FILLER_252_664 ();
 FILLCELL_X32 FILLER_252_696 ();
 FILLCELL_X32 FILLER_252_728 ();
 FILLCELL_X32 FILLER_252_760 ();
 FILLCELL_X32 FILLER_252_792 ();
 FILLCELL_X32 FILLER_252_824 ();
 FILLCELL_X32 FILLER_252_856 ();
 FILLCELL_X32 FILLER_252_888 ();
 FILLCELL_X32 FILLER_252_920 ();
 FILLCELL_X32 FILLER_252_952 ();
 FILLCELL_X32 FILLER_252_984 ();
 FILLCELL_X32 FILLER_252_1016 ();
 FILLCELL_X32 FILLER_252_1048 ();
 FILLCELL_X32 FILLER_252_1080 ();
 FILLCELL_X32 FILLER_252_1112 ();
 FILLCELL_X32 FILLER_252_1144 ();
 FILLCELL_X32 FILLER_252_1176 ();
 FILLCELL_X32 FILLER_252_1208 ();
 FILLCELL_X32 FILLER_252_1240 ();
 FILLCELL_X32 FILLER_252_1272 ();
 FILLCELL_X32 FILLER_252_1304 ();
 FILLCELL_X32 FILLER_252_1336 ();
 FILLCELL_X32 FILLER_252_1368 ();
 FILLCELL_X32 FILLER_252_1400 ();
 FILLCELL_X32 FILLER_252_1432 ();
 FILLCELL_X32 FILLER_252_1464 ();
 FILLCELL_X32 FILLER_252_1496 ();
 FILLCELL_X32 FILLER_252_1528 ();
 FILLCELL_X32 FILLER_252_1560 ();
 FILLCELL_X32 FILLER_252_1592 ();
 FILLCELL_X32 FILLER_252_1624 ();
 FILLCELL_X32 FILLER_252_1656 ();
 FILLCELL_X32 FILLER_252_1688 ();
 FILLCELL_X32 FILLER_252_1720 ();
 FILLCELL_X32 FILLER_252_1752 ();
 FILLCELL_X32 FILLER_252_1784 ();
 FILLCELL_X32 FILLER_252_1816 ();
 FILLCELL_X32 FILLER_252_1848 ();
 FILLCELL_X8 FILLER_252_1880 ();
 FILLCELL_X4 FILLER_252_1888 ();
 FILLCELL_X2 FILLER_252_1892 ();
 FILLCELL_X32 FILLER_252_1895 ();
 FILLCELL_X32 FILLER_252_1927 ();
 FILLCELL_X32 FILLER_252_1959 ();
 FILLCELL_X32 FILLER_252_1991 ();
 FILLCELL_X32 FILLER_252_2023 ();
 FILLCELL_X32 FILLER_252_2055 ();
 FILLCELL_X32 FILLER_252_2087 ();
 FILLCELL_X32 FILLER_252_2119 ();
 FILLCELL_X32 FILLER_252_2151 ();
 FILLCELL_X32 FILLER_252_2183 ();
 FILLCELL_X32 FILLER_252_2215 ();
 FILLCELL_X32 FILLER_252_2247 ();
 FILLCELL_X32 FILLER_252_2279 ();
 FILLCELL_X32 FILLER_252_2311 ();
 FILLCELL_X32 FILLER_252_2343 ();
 FILLCELL_X32 FILLER_252_2375 ();
 FILLCELL_X16 FILLER_252_2407 ();
 FILLCELL_X8 FILLER_252_2423 ();
 FILLCELL_X4 FILLER_252_2431 ();
 FILLCELL_X1 FILLER_252_2435 ();
 FILLCELL_X32 FILLER_253_1 ();
 FILLCELL_X32 FILLER_253_33 ();
 FILLCELL_X32 FILLER_253_65 ();
 FILLCELL_X32 FILLER_253_97 ();
 FILLCELL_X32 FILLER_253_129 ();
 FILLCELL_X32 FILLER_253_161 ();
 FILLCELL_X32 FILLER_253_193 ();
 FILLCELL_X32 FILLER_253_225 ();
 FILLCELL_X32 FILLER_253_257 ();
 FILLCELL_X32 FILLER_253_289 ();
 FILLCELL_X32 FILLER_253_321 ();
 FILLCELL_X32 FILLER_253_353 ();
 FILLCELL_X32 FILLER_253_385 ();
 FILLCELL_X32 FILLER_253_417 ();
 FILLCELL_X32 FILLER_253_449 ();
 FILLCELL_X32 FILLER_253_481 ();
 FILLCELL_X32 FILLER_253_513 ();
 FILLCELL_X32 FILLER_253_545 ();
 FILLCELL_X32 FILLER_253_577 ();
 FILLCELL_X32 FILLER_253_609 ();
 FILLCELL_X32 FILLER_253_641 ();
 FILLCELL_X32 FILLER_253_673 ();
 FILLCELL_X32 FILLER_253_705 ();
 FILLCELL_X32 FILLER_253_737 ();
 FILLCELL_X32 FILLER_253_769 ();
 FILLCELL_X32 FILLER_253_801 ();
 FILLCELL_X32 FILLER_253_833 ();
 FILLCELL_X32 FILLER_253_865 ();
 FILLCELL_X32 FILLER_253_897 ();
 FILLCELL_X32 FILLER_253_929 ();
 FILLCELL_X32 FILLER_253_961 ();
 FILLCELL_X32 FILLER_253_993 ();
 FILLCELL_X32 FILLER_253_1025 ();
 FILLCELL_X32 FILLER_253_1057 ();
 FILLCELL_X32 FILLER_253_1089 ();
 FILLCELL_X32 FILLER_253_1121 ();
 FILLCELL_X32 FILLER_253_1153 ();
 FILLCELL_X32 FILLER_253_1185 ();
 FILLCELL_X32 FILLER_253_1217 ();
 FILLCELL_X8 FILLER_253_1249 ();
 FILLCELL_X4 FILLER_253_1257 ();
 FILLCELL_X2 FILLER_253_1261 ();
 FILLCELL_X32 FILLER_253_1264 ();
 FILLCELL_X32 FILLER_253_1296 ();
 FILLCELL_X32 FILLER_253_1328 ();
 FILLCELL_X32 FILLER_253_1360 ();
 FILLCELL_X32 FILLER_253_1392 ();
 FILLCELL_X32 FILLER_253_1424 ();
 FILLCELL_X32 FILLER_253_1456 ();
 FILLCELL_X32 FILLER_253_1488 ();
 FILLCELL_X32 FILLER_253_1520 ();
 FILLCELL_X32 FILLER_253_1552 ();
 FILLCELL_X32 FILLER_253_1584 ();
 FILLCELL_X32 FILLER_253_1616 ();
 FILLCELL_X32 FILLER_253_1648 ();
 FILLCELL_X32 FILLER_253_1680 ();
 FILLCELL_X32 FILLER_253_1712 ();
 FILLCELL_X32 FILLER_253_1744 ();
 FILLCELL_X32 FILLER_253_1776 ();
 FILLCELL_X32 FILLER_253_1808 ();
 FILLCELL_X32 FILLER_253_1840 ();
 FILLCELL_X32 FILLER_253_1872 ();
 FILLCELL_X32 FILLER_253_1904 ();
 FILLCELL_X32 FILLER_253_1936 ();
 FILLCELL_X32 FILLER_253_1968 ();
 FILLCELL_X32 FILLER_253_2000 ();
 FILLCELL_X32 FILLER_253_2032 ();
 FILLCELL_X32 FILLER_253_2064 ();
 FILLCELL_X32 FILLER_253_2096 ();
 FILLCELL_X32 FILLER_253_2128 ();
 FILLCELL_X32 FILLER_253_2160 ();
 FILLCELL_X32 FILLER_253_2192 ();
 FILLCELL_X32 FILLER_253_2224 ();
 FILLCELL_X32 FILLER_253_2256 ();
 FILLCELL_X32 FILLER_253_2288 ();
 FILLCELL_X32 FILLER_253_2320 ();
 FILLCELL_X32 FILLER_253_2352 ();
 FILLCELL_X32 FILLER_253_2384 ();
 FILLCELL_X16 FILLER_253_2416 ();
 FILLCELL_X4 FILLER_253_2432 ();
 FILLCELL_X32 FILLER_254_1 ();
 FILLCELL_X32 FILLER_254_33 ();
 FILLCELL_X32 FILLER_254_65 ();
 FILLCELL_X32 FILLER_254_97 ();
 FILLCELL_X32 FILLER_254_129 ();
 FILLCELL_X32 FILLER_254_161 ();
 FILLCELL_X32 FILLER_254_193 ();
 FILLCELL_X32 FILLER_254_225 ();
 FILLCELL_X32 FILLER_254_257 ();
 FILLCELL_X32 FILLER_254_289 ();
 FILLCELL_X32 FILLER_254_321 ();
 FILLCELL_X32 FILLER_254_353 ();
 FILLCELL_X32 FILLER_254_385 ();
 FILLCELL_X32 FILLER_254_417 ();
 FILLCELL_X32 FILLER_254_449 ();
 FILLCELL_X32 FILLER_254_481 ();
 FILLCELL_X32 FILLER_254_513 ();
 FILLCELL_X32 FILLER_254_545 ();
 FILLCELL_X32 FILLER_254_577 ();
 FILLCELL_X16 FILLER_254_609 ();
 FILLCELL_X4 FILLER_254_625 ();
 FILLCELL_X2 FILLER_254_629 ();
 FILLCELL_X32 FILLER_254_632 ();
 FILLCELL_X32 FILLER_254_664 ();
 FILLCELL_X32 FILLER_254_696 ();
 FILLCELL_X32 FILLER_254_728 ();
 FILLCELL_X32 FILLER_254_760 ();
 FILLCELL_X32 FILLER_254_792 ();
 FILLCELL_X32 FILLER_254_824 ();
 FILLCELL_X32 FILLER_254_856 ();
 FILLCELL_X32 FILLER_254_888 ();
 FILLCELL_X32 FILLER_254_920 ();
 FILLCELL_X32 FILLER_254_952 ();
 FILLCELL_X32 FILLER_254_984 ();
 FILLCELL_X32 FILLER_254_1016 ();
 FILLCELL_X32 FILLER_254_1048 ();
 FILLCELL_X32 FILLER_254_1080 ();
 FILLCELL_X32 FILLER_254_1112 ();
 FILLCELL_X32 FILLER_254_1144 ();
 FILLCELL_X32 FILLER_254_1176 ();
 FILLCELL_X32 FILLER_254_1208 ();
 FILLCELL_X32 FILLER_254_1240 ();
 FILLCELL_X32 FILLER_254_1272 ();
 FILLCELL_X32 FILLER_254_1304 ();
 FILLCELL_X32 FILLER_254_1336 ();
 FILLCELL_X32 FILLER_254_1368 ();
 FILLCELL_X32 FILLER_254_1400 ();
 FILLCELL_X32 FILLER_254_1432 ();
 FILLCELL_X32 FILLER_254_1464 ();
 FILLCELL_X32 FILLER_254_1496 ();
 FILLCELL_X32 FILLER_254_1528 ();
 FILLCELL_X32 FILLER_254_1560 ();
 FILLCELL_X32 FILLER_254_1592 ();
 FILLCELL_X32 FILLER_254_1624 ();
 FILLCELL_X32 FILLER_254_1656 ();
 FILLCELL_X32 FILLER_254_1688 ();
 FILLCELL_X32 FILLER_254_1720 ();
 FILLCELL_X32 FILLER_254_1752 ();
 FILLCELL_X32 FILLER_254_1784 ();
 FILLCELL_X32 FILLER_254_1816 ();
 FILLCELL_X32 FILLER_254_1848 ();
 FILLCELL_X8 FILLER_254_1880 ();
 FILLCELL_X4 FILLER_254_1888 ();
 FILLCELL_X2 FILLER_254_1892 ();
 FILLCELL_X32 FILLER_254_1895 ();
 FILLCELL_X32 FILLER_254_1927 ();
 FILLCELL_X32 FILLER_254_1959 ();
 FILLCELL_X32 FILLER_254_1991 ();
 FILLCELL_X32 FILLER_254_2023 ();
 FILLCELL_X32 FILLER_254_2055 ();
 FILLCELL_X32 FILLER_254_2087 ();
 FILLCELL_X32 FILLER_254_2119 ();
 FILLCELL_X32 FILLER_254_2151 ();
 FILLCELL_X32 FILLER_254_2183 ();
 FILLCELL_X32 FILLER_254_2215 ();
 FILLCELL_X32 FILLER_254_2247 ();
 FILLCELL_X32 FILLER_254_2279 ();
 FILLCELL_X32 FILLER_254_2311 ();
 FILLCELL_X32 FILLER_254_2343 ();
 FILLCELL_X32 FILLER_254_2375 ();
 FILLCELL_X16 FILLER_254_2407 ();
 FILLCELL_X8 FILLER_254_2423 ();
 FILLCELL_X4 FILLER_254_2431 ();
 FILLCELL_X1 FILLER_254_2435 ();
 FILLCELL_X32 FILLER_255_1 ();
 FILLCELL_X32 FILLER_255_33 ();
 FILLCELL_X32 FILLER_255_65 ();
 FILLCELL_X32 FILLER_255_97 ();
 FILLCELL_X32 FILLER_255_129 ();
 FILLCELL_X32 FILLER_255_161 ();
 FILLCELL_X32 FILLER_255_193 ();
 FILLCELL_X32 FILLER_255_225 ();
 FILLCELL_X32 FILLER_255_257 ();
 FILLCELL_X32 FILLER_255_289 ();
 FILLCELL_X32 FILLER_255_321 ();
 FILLCELL_X32 FILLER_255_353 ();
 FILLCELL_X32 FILLER_255_385 ();
 FILLCELL_X32 FILLER_255_417 ();
 FILLCELL_X32 FILLER_255_449 ();
 FILLCELL_X32 FILLER_255_481 ();
 FILLCELL_X32 FILLER_255_513 ();
 FILLCELL_X32 FILLER_255_545 ();
 FILLCELL_X32 FILLER_255_577 ();
 FILLCELL_X32 FILLER_255_609 ();
 FILLCELL_X32 FILLER_255_641 ();
 FILLCELL_X32 FILLER_255_673 ();
 FILLCELL_X32 FILLER_255_705 ();
 FILLCELL_X32 FILLER_255_737 ();
 FILLCELL_X32 FILLER_255_769 ();
 FILLCELL_X32 FILLER_255_801 ();
 FILLCELL_X32 FILLER_255_833 ();
 FILLCELL_X32 FILLER_255_865 ();
 FILLCELL_X32 FILLER_255_897 ();
 FILLCELL_X32 FILLER_255_929 ();
 FILLCELL_X32 FILLER_255_961 ();
 FILLCELL_X32 FILLER_255_993 ();
 FILLCELL_X32 FILLER_255_1025 ();
 FILLCELL_X32 FILLER_255_1057 ();
 FILLCELL_X32 FILLER_255_1089 ();
 FILLCELL_X32 FILLER_255_1121 ();
 FILLCELL_X32 FILLER_255_1153 ();
 FILLCELL_X32 FILLER_255_1185 ();
 FILLCELL_X32 FILLER_255_1217 ();
 FILLCELL_X8 FILLER_255_1249 ();
 FILLCELL_X4 FILLER_255_1257 ();
 FILLCELL_X2 FILLER_255_1261 ();
 FILLCELL_X32 FILLER_255_1264 ();
 FILLCELL_X32 FILLER_255_1296 ();
 FILLCELL_X32 FILLER_255_1328 ();
 FILLCELL_X32 FILLER_255_1360 ();
 FILLCELL_X32 FILLER_255_1392 ();
 FILLCELL_X32 FILLER_255_1424 ();
 FILLCELL_X32 FILLER_255_1456 ();
 FILLCELL_X32 FILLER_255_1488 ();
 FILLCELL_X32 FILLER_255_1520 ();
 FILLCELL_X32 FILLER_255_1552 ();
 FILLCELL_X32 FILLER_255_1584 ();
 FILLCELL_X32 FILLER_255_1616 ();
 FILLCELL_X32 FILLER_255_1648 ();
 FILLCELL_X32 FILLER_255_1680 ();
 FILLCELL_X32 FILLER_255_1712 ();
 FILLCELL_X32 FILLER_255_1744 ();
 FILLCELL_X32 FILLER_255_1776 ();
 FILLCELL_X32 FILLER_255_1808 ();
 FILLCELL_X32 FILLER_255_1840 ();
 FILLCELL_X32 FILLER_255_1872 ();
 FILLCELL_X32 FILLER_255_1904 ();
 FILLCELL_X32 FILLER_255_1936 ();
 FILLCELL_X32 FILLER_255_1968 ();
 FILLCELL_X32 FILLER_255_2000 ();
 FILLCELL_X32 FILLER_255_2032 ();
 FILLCELL_X32 FILLER_255_2064 ();
 FILLCELL_X32 FILLER_255_2096 ();
 FILLCELL_X32 FILLER_255_2128 ();
 FILLCELL_X32 FILLER_255_2160 ();
 FILLCELL_X32 FILLER_255_2192 ();
 FILLCELL_X32 FILLER_255_2224 ();
 FILLCELL_X32 FILLER_255_2256 ();
 FILLCELL_X32 FILLER_255_2288 ();
 FILLCELL_X32 FILLER_255_2320 ();
 FILLCELL_X32 FILLER_255_2352 ();
 FILLCELL_X32 FILLER_255_2384 ();
 FILLCELL_X16 FILLER_255_2416 ();
 FILLCELL_X4 FILLER_255_2432 ();
 FILLCELL_X32 FILLER_256_1 ();
 FILLCELL_X32 FILLER_256_33 ();
 FILLCELL_X32 FILLER_256_65 ();
 FILLCELL_X32 FILLER_256_97 ();
 FILLCELL_X32 FILLER_256_129 ();
 FILLCELL_X32 FILLER_256_161 ();
 FILLCELL_X32 FILLER_256_193 ();
 FILLCELL_X32 FILLER_256_225 ();
 FILLCELL_X32 FILLER_256_257 ();
 FILLCELL_X32 FILLER_256_289 ();
 FILLCELL_X32 FILLER_256_321 ();
 FILLCELL_X32 FILLER_256_353 ();
 FILLCELL_X32 FILLER_256_385 ();
 FILLCELL_X32 FILLER_256_417 ();
 FILLCELL_X32 FILLER_256_449 ();
 FILLCELL_X32 FILLER_256_481 ();
 FILLCELL_X32 FILLER_256_513 ();
 FILLCELL_X32 FILLER_256_545 ();
 FILLCELL_X32 FILLER_256_577 ();
 FILLCELL_X16 FILLER_256_609 ();
 FILLCELL_X4 FILLER_256_625 ();
 FILLCELL_X2 FILLER_256_629 ();
 FILLCELL_X32 FILLER_256_632 ();
 FILLCELL_X32 FILLER_256_664 ();
 FILLCELL_X32 FILLER_256_696 ();
 FILLCELL_X32 FILLER_256_728 ();
 FILLCELL_X32 FILLER_256_760 ();
 FILLCELL_X32 FILLER_256_792 ();
 FILLCELL_X32 FILLER_256_824 ();
 FILLCELL_X32 FILLER_256_856 ();
 FILLCELL_X32 FILLER_256_888 ();
 FILLCELL_X32 FILLER_256_920 ();
 FILLCELL_X32 FILLER_256_952 ();
 FILLCELL_X32 FILLER_256_984 ();
 FILLCELL_X32 FILLER_256_1016 ();
 FILLCELL_X32 FILLER_256_1048 ();
 FILLCELL_X32 FILLER_256_1080 ();
 FILLCELL_X32 FILLER_256_1112 ();
 FILLCELL_X32 FILLER_256_1144 ();
 FILLCELL_X32 FILLER_256_1176 ();
 FILLCELL_X32 FILLER_256_1208 ();
 FILLCELL_X32 FILLER_256_1240 ();
 FILLCELL_X32 FILLER_256_1272 ();
 FILLCELL_X32 FILLER_256_1304 ();
 FILLCELL_X32 FILLER_256_1336 ();
 FILLCELL_X32 FILLER_256_1368 ();
 FILLCELL_X32 FILLER_256_1400 ();
 FILLCELL_X32 FILLER_256_1432 ();
 FILLCELL_X32 FILLER_256_1464 ();
 FILLCELL_X32 FILLER_256_1496 ();
 FILLCELL_X32 FILLER_256_1528 ();
 FILLCELL_X32 FILLER_256_1560 ();
 FILLCELL_X32 FILLER_256_1592 ();
 FILLCELL_X32 FILLER_256_1624 ();
 FILLCELL_X32 FILLER_256_1656 ();
 FILLCELL_X32 FILLER_256_1688 ();
 FILLCELL_X32 FILLER_256_1720 ();
 FILLCELL_X32 FILLER_256_1752 ();
 FILLCELL_X32 FILLER_256_1784 ();
 FILLCELL_X32 FILLER_256_1816 ();
 FILLCELL_X32 FILLER_256_1848 ();
 FILLCELL_X8 FILLER_256_1880 ();
 FILLCELL_X4 FILLER_256_1888 ();
 FILLCELL_X2 FILLER_256_1892 ();
 FILLCELL_X32 FILLER_256_1895 ();
 FILLCELL_X32 FILLER_256_1927 ();
 FILLCELL_X32 FILLER_256_1959 ();
 FILLCELL_X32 FILLER_256_1991 ();
 FILLCELL_X32 FILLER_256_2023 ();
 FILLCELL_X32 FILLER_256_2055 ();
 FILLCELL_X32 FILLER_256_2087 ();
 FILLCELL_X32 FILLER_256_2119 ();
 FILLCELL_X32 FILLER_256_2151 ();
 FILLCELL_X32 FILLER_256_2183 ();
 FILLCELL_X32 FILLER_256_2215 ();
 FILLCELL_X32 FILLER_256_2247 ();
 FILLCELL_X32 FILLER_256_2279 ();
 FILLCELL_X32 FILLER_256_2311 ();
 FILLCELL_X32 FILLER_256_2343 ();
 FILLCELL_X32 FILLER_256_2375 ();
 FILLCELL_X16 FILLER_256_2407 ();
 FILLCELL_X8 FILLER_256_2423 ();
 FILLCELL_X4 FILLER_256_2431 ();
 FILLCELL_X1 FILLER_256_2435 ();
 FILLCELL_X32 FILLER_257_1 ();
 FILLCELL_X32 FILLER_257_33 ();
 FILLCELL_X32 FILLER_257_65 ();
 FILLCELL_X32 FILLER_257_97 ();
 FILLCELL_X32 FILLER_257_129 ();
 FILLCELL_X32 FILLER_257_161 ();
 FILLCELL_X32 FILLER_257_193 ();
 FILLCELL_X32 FILLER_257_225 ();
 FILLCELL_X32 FILLER_257_257 ();
 FILLCELL_X32 FILLER_257_289 ();
 FILLCELL_X32 FILLER_257_321 ();
 FILLCELL_X32 FILLER_257_353 ();
 FILLCELL_X32 FILLER_257_385 ();
 FILLCELL_X32 FILLER_257_417 ();
 FILLCELL_X32 FILLER_257_449 ();
 FILLCELL_X32 FILLER_257_481 ();
 FILLCELL_X32 FILLER_257_513 ();
 FILLCELL_X32 FILLER_257_545 ();
 FILLCELL_X32 FILLER_257_577 ();
 FILLCELL_X32 FILLER_257_609 ();
 FILLCELL_X32 FILLER_257_641 ();
 FILLCELL_X32 FILLER_257_673 ();
 FILLCELL_X32 FILLER_257_705 ();
 FILLCELL_X32 FILLER_257_737 ();
 FILLCELL_X32 FILLER_257_769 ();
 FILLCELL_X32 FILLER_257_801 ();
 FILLCELL_X32 FILLER_257_833 ();
 FILLCELL_X32 FILLER_257_865 ();
 FILLCELL_X32 FILLER_257_897 ();
 FILLCELL_X32 FILLER_257_929 ();
 FILLCELL_X32 FILLER_257_961 ();
 FILLCELL_X32 FILLER_257_993 ();
 FILLCELL_X32 FILLER_257_1025 ();
 FILLCELL_X32 FILLER_257_1057 ();
 FILLCELL_X32 FILLER_257_1089 ();
 FILLCELL_X32 FILLER_257_1121 ();
 FILLCELL_X32 FILLER_257_1153 ();
 FILLCELL_X32 FILLER_257_1185 ();
 FILLCELL_X32 FILLER_257_1217 ();
 FILLCELL_X8 FILLER_257_1249 ();
 FILLCELL_X4 FILLER_257_1257 ();
 FILLCELL_X2 FILLER_257_1261 ();
 FILLCELL_X32 FILLER_257_1264 ();
 FILLCELL_X32 FILLER_257_1296 ();
 FILLCELL_X32 FILLER_257_1328 ();
 FILLCELL_X32 FILLER_257_1360 ();
 FILLCELL_X32 FILLER_257_1392 ();
 FILLCELL_X32 FILLER_257_1424 ();
 FILLCELL_X32 FILLER_257_1456 ();
 FILLCELL_X32 FILLER_257_1488 ();
 FILLCELL_X32 FILLER_257_1520 ();
 FILLCELL_X32 FILLER_257_1552 ();
 FILLCELL_X32 FILLER_257_1584 ();
 FILLCELL_X32 FILLER_257_1616 ();
 FILLCELL_X32 FILLER_257_1648 ();
 FILLCELL_X32 FILLER_257_1680 ();
 FILLCELL_X32 FILLER_257_1712 ();
 FILLCELL_X32 FILLER_257_1744 ();
 FILLCELL_X32 FILLER_257_1776 ();
 FILLCELL_X32 FILLER_257_1808 ();
 FILLCELL_X32 FILLER_257_1840 ();
 FILLCELL_X32 FILLER_257_1872 ();
 FILLCELL_X32 FILLER_257_1904 ();
 FILLCELL_X32 FILLER_257_1936 ();
 FILLCELL_X32 FILLER_257_1968 ();
 FILLCELL_X32 FILLER_257_2000 ();
 FILLCELL_X32 FILLER_257_2032 ();
 FILLCELL_X32 FILLER_257_2064 ();
 FILLCELL_X32 FILLER_257_2096 ();
 FILLCELL_X32 FILLER_257_2128 ();
 FILLCELL_X32 FILLER_257_2160 ();
 FILLCELL_X32 FILLER_257_2192 ();
 FILLCELL_X32 FILLER_257_2224 ();
 FILLCELL_X32 FILLER_257_2256 ();
 FILLCELL_X32 FILLER_257_2288 ();
 FILLCELL_X32 FILLER_257_2320 ();
 FILLCELL_X32 FILLER_257_2352 ();
 FILLCELL_X32 FILLER_257_2384 ();
 FILLCELL_X16 FILLER_257_2416 ();
 FILLCELL_X4 FILLER_257_2432 ();
 FILLCELL_X32 FILLER_258_1 ();
 FILLCELL_X32 FILLER_258_33 ();
 FILLCELL_X32 FILLER_258_65 ();
 FILLCELL_X32 FILLER_258_97 ();
 FILLCELL_X32 FILLER_258_129 ();
 FILLCELL_X32 FILLER_258_161 ();
 FILLCELL_X32 FILLER_258_193 ();
 FILLCELL_X32 FILLER_258_225 ();
 FILLCELL_X32 FILLER_258_257 ();
 FILLCELL_X32 FILLER_258_289 ();
 FILLCELL_X32 FILLER_258_321 ();
 FILLCELL_X32 FILLER_258_353 ();
 FILLCELL_X32 FILLER_258_385 ();
 FILLCELL_X32 FILLER_258_417 ();
 FILLCELL_X32 FILLER_258_449 ();
 FILLCELL_X32 FILLER_258_481 ();
 FILLCELL_X32 FILLER_258_513 ();
 FILLCELL_X32 FILLER_258_545 ();
 FILLCELL_X32 FILLER_258_577 ();
 FILLCELL_X16 FILLER_258_609 ();
 FILLCELL_X4 FILLER_258_625 ();
 FILLCELL_X2 FILLER_258_629 ();
 FILLCELL_X32 FILLER_258_632 ();
 FILLCELL_X32 FILLER_258_664 ();
 FILLCELL_X32 FILLER_258_696 ();
 FILLCELL_X32 FILLER_258_728 ();
 FILLCELL_X32 FILLER_258_760 ();
 FILLCELL_X32 FILLER_258_792 ();
 FILLCELL_X32 FILLER_258_824 ();
 FILLCELL_X32 FILLER_258_856 ();
 FILLCELL_X32 FILLER_258_888 ();
 FILLCELL_X32 FILLER_258_920 ();
 FILLCELL_X32 FILLER_258_952 ();
 FILLCELL_X32 FILLER_258_984 ();
 FILLCELL_X32 FILLER_258_1016 ();
 FILLCELL_X32 FILLER_258_1048 ();
 FILLCELL_X32 FILLER_258_1080 ();
 FILLCELL_X32 FILLER_258_1112 ();
 FILLCELL_X32 FILLER_258_1144 ();
 FILLCELL_X32 FILLER_258_1176 ();
 FILLCELL_X32 FILLER_258_1208 ();
 FILLCELL_X32 FILLER_258_1240 ();
 FILLCELL_X32 FILLER_258_1272 ();
 FILLCELL_X32 FILLER_258_1304 ();
 FILLCELL_X32 FILLER_258_1336 ();
 FILLCELL_X32 FILLER_258_1368 ();
 FILLCELL_X32 FILLER_258_1400 ();
 FILLCELL_X32 FILLER_258_1432 ();
 FILLCELL_X32 FILLER_258_1464 ();
 FILLCELL_X32 FILLER_258_1496 ();
 FILLCELL_X32 FILLER_258_1528 ();
 FILLCELL_X32 FILLER_258_1560 ();
 FILLCELL_X32 FILLER_258_1592 ();
 FILLCELL_X32 FILLER_258_1624 ();
 FILLCELL_X32 FILLER_258_1656 ();
 FILLCELL_X32 FILLER_258_1688 ();
 FILLCELL_X32 FILLER_258_1720 ();
 FILLCELL_X32 FILLER_258_1752 ();
 FILLCELL_X32 FILLER_258_1784 ();
 FILLCELL_X32 FILLER_258_1816 ();
 FILLCELL_X32 FILLER_258_1848 ();
 FILLCELL_X8 FILLER_258_1880 ();
 FILLCELL_X4 FILLER_258_1888 ();
 FILLCELL_X2 FILLER_258_1892 ();
 FILLCELL_X32 FILLER_258_1895 ();
 FILLCELL_X32 FILLER_258_1927 ();
 FILLCELL_X32 FILLER_258_1959 ();
 FILLCELL_X32 FILLER_258_1991 ();
 FILLCELL_X32 FILLER_258_2023 ();
 FILLCELL_X32 FILLER_258_2055 ();
 FILLCELL_X32 FILLER_258_2087 ();
 FILLCELL_X32 FILLER_258_2119 ();
 FILLCELL_X32 FILLER_258_2151 ();
 FILLCELL_X32 FILLER_258_2183 ();
 FILLCELL_X32 FILLER_258_2215 ();
 FILLCELL_X32 FILLER_258_2247 ();
 FILLCELL_X32 FILLER_258_2279 ();
 FILLCELL_X32 FILLER_258_2311 ();
 FILLCELL_X32 FILLER_258_2343 ();
 FILLCELL_X32 FILLER_258_2375 ();
 FILLCELL_X16 FILLER_258_2407 ();
 FILLCELL_X8 FILLER_258_2423 ();
 FILLCELL_X4 FILLER_258_2431 ();
 FILLCELL_X1 FILLER_258_2435 ();
 FILLCELL_X32 FILLER_259_1 ();
 FILLCELL_X32 FILLER_259_33 ();
 FILLCELL_X32 FILLER_259_65 ();
 FILLCELL_X32 FILLER_259_97 ();
 FILLCELL_X32 FILLER_259_129 ();
 FILLCELL_X32 FILLER_259_161 ();
 FILLCELL_X32 FILLER_259_193 ();
 FILLCELL_X32 FILLER_259_225 ();
 FILLCELL_X32 FILLER_259_257 ();
 FILLCELL_X32 FILLER_259_289 ();
 FILLCELL_X32 FILLER_259_321 ();
 FILLCELL_X32 FILLER_259_353 ();
 FILLCELL_X32 FILLER_259_385 ();
 FILLCELL_X32 FILLER_259_417 ();
 FILLCELL_X32 FILLER_259_449 ();
 FILLCELL_X32 FILLER_259_481 ();
 FILLCELL_X32 FILLER_259_513 ();
 FILLCELL_X32 FILLER_259_545 ();
 FILLCELL_X32 FILLER_259_577 ();
 FILLCELL_X32 FILLER_259_609 ();
 FILLCELL_X32 FILLER_259_641 ();
 FILLCELL_X32 FILLER_259_673 ();
 FILLCELL_X32 FILLER_259_705 ();
 FILLCELL_X32 FILLER_259_737 ();
 FILLCELL_X32 FILLER_259_769 ();
 FILLCELL_X32 FILLER_259_801 ();
 FILLCELL_X32 FILLER_259_833 ();
 FILLCELL_X32 FILLER_259_865 ();
 FILLCELL_X32 FILLER_259_897 ();
 FILLCELL_X32 FILLER_259_929 ();
 FILLCELL_X32 FILLER_259_961 ();
 FILLCELL_X32 FILLER_259_993 ();
 FILLCELL_X32 FILLER_259_1025 ();
 FILLCELL_X32 FILLER_259_1057 ();
 FILLCELL_X32 FILLER_259_1089 ();
 FILLCELL_X32 FILLER_259_1121 ();
 FILLCELL_X32 FILLER_259_1153 ();
 FILLCELL_X32 FILLER_259_1185 ();
 FILLCELL_X32 FILLER_259_1217 ();
 FILLCELL_X8 FILLER_259_1249 ();
 FILLCELL_X4 FILLER_259_1257 ();
 FILLCELL_X2 FILLER_259_1261 ();
 FILLCELL_X32 FILLER_259_1264 ();
 FILLCELL_X32 FILLER_259_1296 ();
 FILLCELL_X32 FILLER_259_1328 ();
 FILLCELL_X32 FILLER_259_1360 ();
 FILLCELL_X32 FILLER_259_1392 ();
 FILLCELL_X32 FILLER_259_1424 ();
 FILLCELL_X32 FILLER_259_1456 ();
 FILLCELL_X32 FILLER_259_1488 ();
 FILLCELL_X32 FILLER_259_1520 ();
 FILLCELL_X32 FILLER_259_1552 ();
 FILLCELL_X32 FILLER_259_1584 ();
 FILLCELL_X32 FILLER_259_1616 ();
 FILLCELL_X32 FILLER_259_1648 ();
 FILLCELL_X32 FILLER_259_1680 ();
 FILLCELL_X32 FILLER_259_1712 ();
 FILLCELL_X32 FILLER_259_1744 ();
 FILLCELL_X32 FILLER_259_1776 ();
 FILLCELL_X32 FILLER_259_1808 ();
 FILLCELL_X32 FILLER_259_1840 ();
 FILLCELL_X32 FILLER_259_1872 ();
 FILLCELL_X32 FILLER_259_1904 ();
 FILLCELL_X32 FILLER_259_1936 ();
 FILLCELL_X32 FILLER_259_1968 ();
 FILLCELL_X32 FILLER_259_2000 ();
 FILLCELL_X32 FILLER_259_2032 ();
 FILLCELL_X32 FILLER_259_2064 ();
 FILLCELL_X32 FILLER_259_2096 ();
 FILLCELL_X32 FILLER_259_2128 ();
 FILLCELL_X32 FILLER_259_2160 ();
 FILLCELL_X32 FILLER_259_2192 ();
 FILLCELL_X32 FILLER_259_2224 ();
 FILLCELL_X32 FILLER_259_2256 ();
 FILLCELL_X32 FILLER_259_2288 ();
 FILLCELL_X32 FILLER_259_2320 ();
 FILLCELL_X32 FILLER_259_2352 ();
 FILLCELL_X32 FILLER_259_2384 ();
 FILLCELL_X16 FILLER_259_2416 ();
 FILLCELL_X4 FILLER_259_2432 ();
 FILLCELL_X32 FILLER_260_1 ();
 FILLCELL_X32 FILLER_260_33 ();
 FILLCELL_X32 FILLER_260_65 ();
 FILLCELL_X32 FILLER_260_97 ();
 FILLCELL_X32 FILLER_260_129 ();
 FILLCELL_X32 FILLER_260_161 ();
 FILLCELL_X32 FILLER_260_193 ();
 FILLCELL_X32 FILLER_260_225 ();
 FILLCELL_X32 FILLER_260_257 ();
 FILLCELL_X32 FILLER_260_289 ();
 FILLCELL_X32 FILLER_260_321 ();
 FILLCELL_X32 FILLER_260_353 ();
 FILLCELL_X32 FILLER_260_385 ();
 FILLCELL_X32 FILLER_260_417 ();
 FILLCELL_X32 FILLER_260_449 ();
 FILLCELL_X32 FILLER_260_481 ();
 FILLCELL_X32 FILLER_260_513 ();
 FILLCELL_X32 FILLER_260_545 ();
 FILLCELL_X32 FILLER_260_577 ();
 FILLCELL_X16 FILLER_260_609 ();
 FILLCELL_X4 FILLER_260_625 ();
 FILLCELL_X2 FILLER_260_629 ();
 FILLCELL_X32 FILLER_260_632 ();
 FILLCELL_X32 FILLER_260_664 ();
 FILLCELL_X32 FILLER_260_696 ();
 FILLCELL_X32 FILLER_260_728 ();
 FILLCELL_X32 FILLER_260_760 ();
 FILLCELL_X32 FILLER_260_792 ();
 FILLCELL_X32 FILLER_260_824 ();
 FILLCELL_X32 FILLER_260_856 ();
 FILLCELL_X32 FILLER_260_888 ();
 FILLCELL_X32 FILLER_260_920 ();
 FILLCELL_X32 FILLER_260_952 ();
 FILLCELL_X32 FILLER_260_984 ();
 FILLCELL_X32 FILLER_260_1016 ();
 FILLCELL_X32 FILLER_260_1048 ();
 FILLCELL_X32 FILLER_260_1080 ();
 FILLCELL_X32 FILLER_260_1112 ();
 FILLCELL_X32 FILLER_260_1144 ();
 FILLCELL_X32 FILLER_260_1176 ();
 FILLCELL_X32 FILLER_260_1208 ();
 FILLCELL_X32 FILLER_260_1240 ();
 FILLCELL_X32 FILLER_260_1272 ();
 FILLCELL_X32 FILLER_260_1304 ();
 FILLCELL_X32 FILLER_260_1336 ();
 FILLCELL_X32 FILLER_260_1368 ();
 FILLCELL_X32 FILLER_260_1400 ();
 FILLCELL_X32 FILLER_260_1432 ();
 FILLCELL_X32 FILLER_260_1464 ();
 FILLCELL_X32 FILLER_260_1496 ();
 FILLCELL_X32 FILLER_260_1528 ();
 FILLCELL_X32 FILLER_260_1560 ();
 FILLCELL_X32 FILLER_260_1592 ();
 FILLCELL_X32 FILLER_260_1624 ();
 FILLCELL_X32 FILLER_260_1656 ();
 FILLCELL_X32 FILLER_260_1688 ();
 FILLCELL_X32 FILLER_260_1720 ();
 FILLCELL_X32 FILLER_260_1752 ();
 FILLCELL_X32 FILLER_260_1784 ();
 FILLCELL_X32 FILLER_260_1816 ();
 FILLCELL_X32 FILLER_260_1848 ();
 FILLCELL_X8 FILLER_260_1880 ();
 FILLCELL_X4 FILLER_260_1888 ();
 FILLCELL_X2 FILLER_260_1892 ();
 FILLCELL_X32 FILLER_260_1895 ();
 FILLCELL_X32 FILLER_260_1927 ();
 FILLCELL_X32 FILLER_260_1959 ();
 FILLCELL_X32 FILLER_260_1991 ();
 FILLCELL_X32 FILLER_260_2023 ();
 FILLCELL_X32 FILLER_260_2055 ();
 FILLCELL_X32 FILLER_260_2087 ();
 FILLCELL_X32 FILLER_260_2119 ();
 FILLCELL_X32 FILLER_260_2151 ();
 FILLCELL_X32 FILLER_260_2183 ();
 FILLCELL_X32 FILLER_260_2215 ();
 FILLCELL_X32 FILLER_260_2247 ();
 FILLCELL_X32 FILLER_260_2279 ();
 FILLCELL_X32 FILLER_260_2311 ();
 FILLCELL_X32 FILLER_260_2343 ();
 FILLCELL_X32 FILLER_260_2375 ();
 FILLCELL_X16 FILLER_260_2407 ();
 FILLCELL_X8 FILLER_260_2423 ();
 FILLCELL_X4 FILLER_260_2431 ();
 FILLCELL_X1 FILLER_260_2435 ();
 FILLCELL_X32 FILLER_261_1 ();
 FILLCELL_X32 FILLER_261_33 ();
 FILLCELL_X32 FILLER_261_65 ();
 FILLCELL_X32 FILLER_261_97 ();
 FILLCELL_X32 FILLER_261_129 ();
 FILLCELL_X32 FILLER_261_161 ();
 FILLCELL_X32 FILLER_261_193 ();
 FILLCELL_X32 FILLER_261_225 ();
 FILLCELL_X32 FILLER_261_257 ();
 FILLCELL_X32 FILLER_261_289 ();
 FILLCELL_X32 FILLER_261_321 ();
 FILLCELL_X32 FILLER_261_353 ();
 FILLCELL_X32 FILLER_261_385 ();
 FILLCELL_X32 FILLER_261_417 ();
 FILLCELL_X32 FILLER_261_449 ();
 FILLCELL_X32 FILLER_261_481 ();
 FILLCELL_X32 FILLER_261_513 ();
 FILLCELL_X32 FILLER_261_545 ();
 FILLCELL_X32 FILLER_261_577 ();
 FILLCELL_X32 FILLER_261_609 ();
 FILLCELL_X32 FILLER_261_641 ();
 FILLCELL_X32 FILLER_261_673 ();
 FILLCELL_X32 FILLER_261_705 ();
 FILLCELL_X32 FILLER_261_737 ();
 FILLCELL_X32 FILLER_261_769 ();
 FILLCELL_X32 FILLER_261_801 ();
 FILLCELL_X32 FILLER_261_833 ();
 FILLCELL_X32 FILLER_261_865 ();
 FILLCELL_X32 FILLER_261_897 ();
 FILLCELL_X32 FILLER_261_929 ();
 FILLCELL_X32 FILLER_261_961 ();
 FILLCELL_X32 FILLER_261_993 ();
 FILLCELL_X32 FILLER_261_1025 ();
 FILLCELL_X32 FILLER_261_1057 ();
 FILLCELL_X32 FILLER_261_1089 ();
 FILLCELL_X32 FILLER_261_1121 ();
 FILLCELL_X32 FILLER_261_1153 ();
 FILLCELL_X32 FILLER_261_1185 ();
 FILLCELL_X32 FILLER_261_1217 ();
 FILLCELL_X8 FILLER_261_1249 ();
 FILLCELL_X4 FILLER_261_1257 ();
 FILLCELL_X2 FILLER_261_1261 ();
 FILLCELL_X32 FILLER_261_1264 ();
 FILLCELL_X32 FILLER_261_1296 ();
 FILLCELL_X32 FILLER_261_1328 ();
 FILLCELL_X32 FILLER_261_1360 ();
 FILLCELL_X32 FILLER_261_1392 ();
 FILLCELL_X32 FILLER_261_1424 ();
 FILLCELL_X32 FILLER_261_1456 ();
 FILLCELL_X32 FILLER_261_1488 ();
 FILLCELL_X32 FILLER_261_1520 ();
 FILLCELL_X32 FILLER_261_1552 ();
 FILLCELL_X32 FILLER_261_1584 ();
 FILLCELL_X32 FILLER_261_1616 ();
 FILLCELL_X32 FILLER_261_1648 ();
 FILLCELL_X32 FILLER_261_1680 ();
 FILLCELL_X32 FILLER_261_1712 ();
 FILLCELL_X32 FILLER_261_1744 ();
 FILLCELL_X32 FILLER_261_1776 ();
 FILLCELL_X32 FILLER_261_1808 ();
 FILLCELL_X32 FILLER_261_1840 ();
 FILLCELL_X32 FILLER_261_1872 ();
 FILLCELL_X32 FILLER_261_1904 ();
 FILLCELL_X32 FILLER_261_1936 ();
 FILLCELL_X32 FILLER_261_1968 ();
 FILLCELL_X32 FILLER_261_2000 ();
 FILLCELL_X32 FILLER_261_2032 ();
 FILLCELL_X32 FILLER_261_2064 ();
 FILLCELL_X32 FILLER_261_2096 ();
 FILLCELL_X32 FILLER_261_2128 ();
 FILLCELL_X32 FILLER_261_2160 ();
 FILLCELL_X32 FILLER_261_2192 ();
 FILLCELL_X32 FILLER_261_2224 ();
 FILLCELL_X32 FILLER_261_2256 ();
 FILLCELL_X32 FILLER_261_2288 ();
 FILLCELL_X32 FILLER_261_2320 ();
 FILLCELL_X32 FILLER_261_2352 ();
 FILLCELL_X32 FILLER_261_2384 ();
 FILLCELL_X16 FILLER_261_2416 ();
 FILLCELL_X4 FILLER_261_2432 ();
 FILLCELL_X32 FILLER_262_1 ();
 FILLCELL_X32 FILLER_262_33 ();
 FILLCELL_X32 FILLER_262_65 ();
 FILLCELL_X32 FILLER_262_97 ();
 FILLCELL_X32 FILLER_262_129 ();
 FILLCELL_X32 FILLER_262_161 ();
 FILLCELL_X32 FILLER_262_193 ();
 FILLCELL_X32 FILLER_262_225 ();
 FILLCELL_X32 FILLER_262_257 ();
 FILLCELL_X32 FILLER_262_289 ();
 FILLCELL_X32 FILLER_262_321 ();
 FILLCELL_X32 FILLER_262_353 ();
 FILLCELL_X32 FILLER_262_385 ();
 FILLCELL_X32 FILLER_262_417 ();
 FILLCELL_X32 FILLER_262_449 ();
 FILLCELL_X32 FILLER_262_481 ();
 FILLCELL_X32 FILLER_262_513 ();
 FILLCELL_X32 FILLER_262_545 ();
 FILLCELL_X32 FILLER_262_577 ();
 FILLCELL_X16 FILLER_262_609 ();
 FILLCELL_X4 FILLER_262_625 ();
 FILLCELL_X2 FILLER_262_629 ();
 FILLCELL_X32 FILLER_262_632 ();
 FILLCELL_X32 FILLER_262_664 ();
 FILLCELL_X32 FILLER_262_696 ();
 FILLCELL_X32 FILLER_262_728 ();
 FILLCELL_X32 FILLER_262_760 ();
 FILLCELL_X32 FILLER_262_792 ();
 FILLCELL_X32 FILLER_262_824 ();
 FILLCELL_X32 FILLER_262_856 ();
 FILLCELL_X32 FILLER_262_888 ();
 FILLCELL_X32 FILLER_262_920 ();
 FILLCELL_X32 FILLER_262_952 ();
 FILLCELL_X32 FILLER_262_984 ();
 FILLCELL_X32 FILLER_262_1016 ();
 FILLCELL_X32 FILLER_262_1048 ();
 FILLCELL_X32 FILLER_262_1080 ();
 FILLCELL_X32 FILLER_262_1112 ();
 FILLCELL_X32 FILLER_262_1144 ();
 FILLCELL_X32 FILLER_262_1176 ();
 FILLCELL_X32 FILLER_262_1208 ();
 FILLCELL_X32 FILLER_262_1240 ();
 FILLCELL_X32 FILLER_262_1272 ();
 FILLCELL_X32 FILLER_262_1304 ();
 FILLCELL_X32 FILLER_262_1336 ();
 FILLCELL_X32 FILLER_262_1368 ();
 FILLCELL_X32 FILLER_262_1400 ();
 FILLCELL_X32 FILLER_262_1432 ();
 FILLCELL_X32 FILLER_262_1464 ();
 FILLCELL_X32 FILLER_262_1496 ();
 FILLCELL_X32 FILLER_262_1528 ();
 FILLCELL_X32 FILLER_262_1560 ();
 FILLCELL_X32 FILLER_262_1592 ();
 FILLCELL_X32 FILLER_262_1624 ();
 FILLCELL_X32 FILLER_262_1656 ();
 FILLCELL_X32 FILLER_262_1688 ();
 FILLCELL_X32 FILLER_262_1720 ();
 FILLCELL_X32 FILLER_262_1752 ();
 FILLCELL_X32 FILLER_262_1784 ();
 FILLCELL_X32 FILLER_262_1816 ();
 FILLCELL_X32 FILLER_262_1848 ();
 FILLCELL_X8 FILLER_262_1880 ();
 FILLCELL_X4 FILLER_262_1888 ();
 FILLCELL_X2 FILLER_262_1892 ();
 FILLCELL_X32 FILLER_262_1895 ();
 FILLCELL_X32 FILLER_262_1927 ();
 FILLCELL_X32 FILLER_262_1959 ();
 FILLCELL_X32 FILLER_262_1991 ();
 FILLCELL_X32 FILLER_262_2023 ();
 FILLCELL_X32 FILLER_262_2055 ();
 FILLCELL_X32 FILLER_262_2087 ();
 FILLCELL_X32 FILLER_262_2119 ();
 FILLCELL_X32 FILLER_262_2151 ();
 FILLCELL_X32 FILLER_262_2183 ();
 FILLCELL_X32 FILLER_262_2215 ();
 FILLCELL_X32 FILLER_262_2247 ();
 FILLCELL_X32 FILLER_262_2279 ();
 FILLCELL_X32 FILLER_262_2311 ();
 FILLCELL_X32 FILLER_262_2343 ();
 FILLCELL_X32 FILLER_262_2375 ();
 FILLCELL_X16 FILLER_262_2407 ();
 FILLCELL_X8 FILLER_262_2423 ();
 FILLCELL_X4 FILLER_262_2431 ();
 FILLCELL_X1 FILLER_262_2435 ();
 FILLCELL_X32 FILLER_263_1 ();
 FILLCELL_X32 FILLER_263_33 ();
 FILLCELL_X32 FILLER_263_65 ();
 FILLCELL_X32 FILLER_263_97 ();
 FILLCELL_X32 FILLER_263_129 ();
 FILLCELL_X32 FILLER_263_161 ();
 FILLCELL_X32 FILLER_263_193 ();
 FILLCELL_X32 FILLER_263_225 ();
 FILLCELL_X32 FILLER_263_257 ();
 FILLCELL_X32 FILLER_263_289 ();
 FILLCELL_X32 FILLER_263_321 ();
 FILLCELL_X32 FILLER_263_353 ();
 FILLCELL_X32 FILLER_263_385 ();
 FILLCELL_X32 FILLER_263_417 ();
 FILLCELL_X32 FILLER_263_449 ();
 FILLCELL_X32 FILLER_263_481 ();
 FILLCELL_X32 FILLER_263_513 ();
 FILLCELL_X32 FILLER_263_545 ();
 FILLCELL_X32 FILLER_263_577 ();
 FILLCELL_X32 FILLER_263_609 ();
 FILLCELL_X32 FILLER_263_641 ();
 FILLCELL_X32 FILLER_263_673 ();
 FILLCELL_X32 FILLER_263_705 ();
 FILLCELL_X32 FILLER_263_737 ();
 FILLCELL_X32 FILLER_263_769 ();
 FILLCELL_X32 FILLER_263_801 ();
 FILLCELL_X32 FILLER_263_833 ();
 FILLCELL_X32 FILLER_263_865 ();
 FILLCELL_X32 FILLER_263_897 ();
 FILLCELL_X32 FILLER_263_929 ();
 FILLCELL_X32 FILLER_263_961 ();
 FILLCELL_X32 FILLER_263_993 ();
 FILLCELL_X32 FILLER_263_1025 ();
 FILLCELL_X32 FILLER_263_1057 ();
 FILLCELL_X32 FILLER_263_1089 ();
 FILLCELL_X32 FILLER_263_1121 ();
 FILLCELL_X32 FILLER_263_1153 ();
 FILLCELL_X32 FILLER_263_1185 ();
 FILLCELL_X32 FILLER_263_1217 ();
 FILLCELL_X8 FILLER_263_1249 ();
 FILLCELL_X4 FILLER_263_1257 ();
 FILLCELL_X2 FILLER_263_1261 ();
 FILLCELL_X32 FILLER_263_1264 ();
 FILLCELL_X32 FILLER_263_1296 ();
 FILLCELL_X32 FILLER_263_1328 ();
 FILLCELL_X32 FILLER_263_1360 ();
 FILLCELL_X32 FILLER_263_1392 ();
 FILLCELL_X32 FILLER_263_1424 ();
 FILLCELL_X32 FILLER_263_1456 ();
 FILLCELL_X32 FILLER_263_1488 ();
 FILLCELL_X32 FILLER_263_1520 ();
 FILLCELL_X32 FILLER_263_1552 ();
 FILLCELL_X32 FILLER_263_1584 ();
 FILLCELL_X32 FILLER_263_1616 ();
 FILLCELL_X32 FILLER_263_1648 ();
 FILLCELL_X32 FILLER_263_1680 ();
 FILLCELL_X32 FILLER_263_1712 ();
 FILLCELL_X32 FILLER_263_1744 ();
 FILLCELL_X32 FILLER_263_1776 ();
 FILLCELL_X32 FILLER_263_1808 ();
 FILLCELL_X32 FILLER_263_1840 ();
 FILLCELL_X32 FILLER_263_1872 ();
 FILLCELL_X32 FILLER_263_1904 ();
 FILLCELL_X32 FILLER_263_1936 ();
 FILLCELL_X32 FILLER_263_1968 ();
 FILLCELL_X32 FILLER_263_2000 ();
 FILLCELL_X32 FILLER_263_2032 ();
 FILLCELL_X32 FILLER_263_2064 ();
 FILLCELL_X32 FILLER_263_2096 ();
 FILLCELL_X32 FILLER_263_2128 ();
 FILLCELL_X32 FILLER_263_2160 ();
 FILLCELL_X32 FILLER_263_2192 ();
 FILLCELL_X32 FILLER_263_2224 ();
 FILLCELL_X32 FILLER_263_2256 ();
 FILLCELL_X32 FILLER_263_2288 ();
 FILLCELL_X32 FILLER_263_2320 ();
 FILLCELL_X32 FILLER_263_2352 ();
 FILLCELL_X32 FILLER_263_2384 ();
 FILLCELL_X16 FILLER_263_2416 ();
 FILLCELL_X4 FILLER_263_2432 ();
 FILLCELL_X32 FILLER_264_1 ();
 FILLCELL_X32 FILLER_264_33 ();
 FILLCELL_X32 FILLER_264_65 ();
 FILLCELL_X32 FILLER_264_97 ();
 FILLCELL_X32 FILLER_264_129 ();
 FILLCELL_X32 FILLER_264_161 ();
 FILLCELL_X32 FILLER_264_193 ();
 FILLCELL_X32 FILLER_264_225 ();
 FILLCELL_X32 FILLER_264_257 ();
 FILLCELL_X32 FILLER_264_289 ();
 FILLCELL_X32 FILLER_264_321 ();
 FILLCELL_X32 FILLER_264_353 ();
 FILLCELL_X32 FILLER_264_385 ();
 FILLCELL_X32 FILLER_264_417 ();
 FILLCELL_X32 FILLER_264_449 ();
 FILLCELL_X32 FILLER_264_481 ();
 FILLCELL_X32 FILLER_264_513 ();
 FILLCELL_X32 FILLER_264_545 ();
 FILLCELL_X32 FILLER_264_577 ();
 FILLCELL_X16 FILLER_264_609 ();
 FILLCELL_X4 FILLER_264_625 ();
 FILLCELL_X2 FILLER_264_629 ();
 FILLCELL_X32 FILLER_264_632 ();
 FILLCELL_X32 FILLER_264_664 ();
 FILLCELL_X32 FILLER_264_696 ();
 FILLCELL_X32 FILLER_264_728 ();
 FILLCELL_X32 FILLER_264_760 ();
 FILLCELL_X32 FILLER_264_792 ();
 FILLCELL_X32 FILLER_264_824 ();
 FILLCELL_X32 FILLER_264_856 ();
 FILLCELL_X32 FILLER_264_888 ();
 FILLCELL_X32 FILLER_264_920 ();
 FILLCELL_X32 FILLER_264_952 ();
 FILLCELL_X32 FILLER_264_984 ();
 FILLCELL_X32 FILLER_264_1016 ();
 FILLCELL_X32 FILLER_264_1048 ();
 FILLCELL_X32 FILLER_264_1080 ();
 FILLCELL_X32 FILLER_264_1112 ();
 FILLCELL_X32 FILLER_264_1144 ();
 FILLCELL_X32 FILLER_264_1176 ();
 FILLCELL_X32 FILLER_264_1208 ();
 FILLCELL_X32 FILLER_264_1240 ();
 FILLCELL_X32 FILLER_264_1272 ();
 FILLCELL_X32 FILLER_264_1304 ();
 FILLCELL_X32 FILLER_264_1336 ();
 FILLCELL_X32 FILLER_264_1368 ();
 FILLCELL_X32 FILLER_264_1400 ();
 FILLCELL_X32 FILLER_264_1432 ();
 FILLCELL_X32 FILLER_264_1464 ();
 FILLCELL_X32 FILLER_264_1496 ();
 FILLCELL_X32 FILLER_264_1528 ();
 FILLCELL_X32 FILLER_264_1560 ();
 FILLCELL_X32 FILLER_264_1592 ();
 FILLCELL_X32 FILLER_264_1624 ();
 FILLCELL_X32 FILLER_264_1656 ();
 FILLCELL_X32 FILLER_264_1688 ();
 FILLCELL_X32 FILLER_264_1720 ();
 FILLCELL_X32 FILLER_264_1752 ();
 FILLCELL_X32 FILLER_264_1784 ();
 FILLCELL_X32 FILLER_264_1816 ();
 FILLCELL_X32 FILLER_264_1848 ();
 FILLCELL_X8 FILLER_264_1880 ();
 FILLCELL_X4 FILLER_264_1888 ();
 FILLCELL_X2 FILLER_264_1892 ();
 FILLCELL_X32 FILLER_264_1895 ();
 FILLCELL_X32 FILLER_264_1927 ();
 FILLCELL_X32 FILLER_264_1959 ();
 FILLCELL_X32 FILLER_264_1991 ();
 FILLCELL_X32 FILLER_264_2023 ();
 FILLCELL_X32 FILLER_264_2055 ();
 FILLCELL_X32 FILLER_264_2087 ();
 FILLCELL_X32 FILLER_264_2119 ();
 FILLCELL_X32 FILLER_264_2151 ();
 FILLCELL_X32 FILLER_264_2183 ();
 FILLCELL_X32 FILLER_264_2215 ();
 FILLCELL_X32 FILLER_264_2247 ();
 FILLCELL_X32 FILLER_264_2279 ();
 FILLCELL_X32 FILLER_264_2311 ();
 FILLCELL_X32 FILLER_264_2343 ();
 FILLCELL_X32 FILLER_264_2375 ();
 FILLCELL_X16 FILLER_264_2407 ();
 FILLCELL_X8 FILLER_264_2423 ();
 FILLCELL_X4 FILLER_264_2431 ();
 FILLCELL_X1 FILLER_264_2435 ();
 FILLCELL_X32 FILLER_265_1 ();
 FILLCELL_X32 FILLER_265_33 ();
 FILLCELL_X32 FILLER_265_65 ();
 FILLCELL_X32 FILLER_265_97 ();
 FILLCELL_X32 FILLER_265_129 ();
 FILLCELL_X32 FILLER_265_161 ();
 FILLCELL_X32 FILLER_265_193 ();
 FILLCELL_X32 FILLER_265_225 ();
 FILLCELL_X32 FILLER_265_257 ();
 FILLCELL_X32 FILLER_265_289 ();
 FILLCELL_X32 FILLER_265_321 ();
 FILLCELL_X32 FILLER_265_353 ();
 FILLCELL_X32 FILLER_265_385 ();
 FILLCELL_X32 FILLER_265_417 ();
 FILLCELL_X32 FILLER_265_449 ();
 FILLCELL_X32 FILLER_265_481 ();
 FILLCELL_X32 FILLER_265_513 ();
 FILLCELL_X32 FILLER_265_545 ();
 FILLCELL_X32 FILLER_265_577 ();
 FILLCELL_X32 FILLER_265_609 ();
 FILLCELL_X32 FILLER_265_641 ();
 FILLCELL_X32 FILLER_265_673 ();
 FILLCELL_X32 FILLER_265_705 ();
 FILLCELL_X32 FILLER_265_737 ();
 FILLCELL_X32 FILLER_265_769 ();
 FILLCELL_X32 FILLER_265_801 ();
 FILLCELL_X32 FILLER_265_833 ();
 FILLCELL_X32 FILLER_265_865 ();
 FILLCELL_X32 FILLER_265_897 ();
 FILLCELL_X32 FILLER_265_929 ();
 FILLCELL_X32 FILLER_265_961 ();
 FILLCELL_X32 FILLER_265_993 ();
 FILLCELL_X32 FILLER_265_1025 ();
 FILLCELL_X32 FILLER_265_1057 ();
 FILLCELL_X32 FILLER_265_1089 ();
 FILLCELL_X32 FILLER_265_1121 ();
 FILLCELL_X32 FILLER_265_1153 ();
 FILLCELL_X32 FILLER_265_1185 ();
 FILLCELL_X32 FILLER_265_1217 ();
 FILLCELL_X8 FILLER_265_1249 ();
 FILLCELL_X4 FILLER_265_1257 ();
 FILLCELL_X2 FILLER_265_1261 ();
 FILLCELL_X32 FILLER_265_1264 ();
 FILLCELL_X32 FILLER_265_1296 ();
 FILLCELL_X32 FILLER_265_1328 ();
 FILLCELL_X32 FILLER_265_1360 ();
 FILLCELL_X32 FILLER_265_1392 ();
 FILLCELL_X32 FILLER_265_1424 ();
 FILLCELL_X32 FILLER_265_1456 ();
 FILLCELL_X32 FILLER_265_1488 ();
 FILLCELL_X32 FILLER_265_1520 ();
 FILLCELL_X32 FILLER_265_1552 ();
 FILLCELL_X32 FILLER_265_1584 ();
 FILLCELL_X32 FILLER_265_1616 ();
 FILLCELL_X32 FILLER_265_1648 ();
 FILLCELL_X32 FILLER_265_1680 ();
 FILLCELL_X32 FILLER_265_1712 ();
 FILLCELL_X32 FILLER_265_1744 ();
 FILLCELL_X32 FILLER_265_1776 ();
 FILLCELL_X32 FILLER_265_1808 ();
 FILLCELL_X32 FILLER_265_1840 ();
 FILLCELL_X32 FILLER_265_1872 ();
 FILLCELL_X32 FILLER_265_1904 ();
 FILLCELL_X32 FILLER_265_1936 ();
 FILLCELL_X32 FILLER_265_1968 ();
 FILLCELL_X32 FILLER_265_2000 ();
 FILLCELL_X32 FILLER_265_2032 ();
 FILLCELL_X32 FILLER_265_2064 ();
 FILLCELL_X32 FILLER_265_2096 ();
 FILLCELL_X32 FILLER_265_2128 ();
 FILLCELL_X32 FILLER_265_2160 ();
 FILLCELL_X32 FILLER_265_2192 ();
 FILLCELL_X32 FILLER_265_2224 ();
 FILLCELL_X32 FILLER_265_2256 ();
 FILLCELL_X32 FILLER_265_2288 ();
 FILLCELL_X32 FILLER_265_2320 ();
 FILLCELL_X32 FILLER_265_2352 ();
 FILLCELL_X32 FILLER_265_2384 ();
 FILLCELL_X16 FILLER_265_2416 ();
 FILLCELL_X4 FILLER_265_2432 ();
 FILLCELL_X32 FILLER_266_1 ();
 FILLCELL_X32 FILLER_266_33 ();
 FILLCELL_X32 FILLER_266_65 ();
 FILLCELL_X32 FILLER_266_97 ();
 FILLCELL_X32 FILLER_266_129 ();
 FILLCELL_X32 FILLER_266_161 ();
 FILLCELL_X32 FILLER_266_193 ();
 FILLCELL_X32 FILLER_266_225 ();
 FILLCELL_X32 FILLER_266_257 ();
 FILLCELL_X32 FILLER_266_289 ();
 FILLCELL_X32 FILLER_266_321 ();
 FILLCELL_X32 FILLER_266_353 ();
 FILLCELL_X32 FILLER_266_385 ();
 FILLCELL_X32 FILLER_266_417 ();
 FILLCELL_X32 FILLER_266_449 ();
 FILLCELL_X32 FILLER_266_481 ();
 FILLCELL_X32 FILLER_266_513 ();
 FILLCELL_X32 FILLER_266_545 ();
 FILLCELL_X32 FILLER_266_577 ();
 FILLCELL_X16 FILLER_266_609 ();
 FILLCELL_X4 FILLER_266_625 ();
 FILLCELL_X2 FILLER_266_629 ();
 FILLCELL_X32 FILLER_266_632 ();
 FILLCELL_X32 FILLER_266_664 ();
 FILLCELL_X32 FILLER_266_696 ();
 FILLCELL_X32 FILLER_266_728 ();
 FILLCELL_X32 FILLER_266_760 ();
 FILLCELL_X32 FILLER_266_792 ();
 FILLCELL_X32 FILLER_266_824 ();
 FILLCELL_X32 FILLER_266_856 ();
 FILLCELL_X32 FILLER_266_888 ();
 FILLCELL_X32 FILLER_266_920 ();
 FILLCELL_X32 FILLER_266_952 ();
 FILLCELL_X32 FILLER_266_984 ();
 FILLCELL_X32 FILLER_266_1016 ();
 FILLCELL_X32 FILLER_266_1048 ();
 FILLCELL_X32 FILLER_266_1080 ();
 FILLCELL_X32 FILLER_266_1112 ();
 FILLCELL_X32 FILLER_266_1144 ();
 FILLCELL_X32 FILLER_266_1176 ();
 FILLCELL_X32 FILLER_266_1208 ();
 FILLCELL_X32 FILLER_266_1240 ();
 FILLCELL_X32 FILLER_266_1272 ();
 FILLCELL_X32 FILLER_266_1304 ();
 FILLCELL_X32 FILLER_266_1336 ();
 FILLCELL_X32 FILLER_266_1368 ();
 FILLCELL_X32 FILLER_266_1400 ();
 FILLCELL_X32 FILLER_266_1432 ();
 FILLCELL_X32 FILLER_266_1464 ();
 FILLCELL_X32 FILLER_266_1496 ();
 FILLCELL_X32 FILLER_266_1528 ();
 FILLCELL_X32 FILLER_266_1560 ();
 FILLCELL_X32 FILLER_266_1592 ();
 FILLCELL_X32 FILLER_266_1624 ();
 FILLCELL_X32 FILLER_266_1656 ();
 FILLCELL_X32 FILLER_266_1688 ();
 FILLCELL_X32 FILLER_266_1720 ();
 FILLCELL_X32 FILLER_266_1752 ();
 FILLCELL_X32 FILLER_266_1784 ();
 FILLCELL_X32 FILLER_266_1816 ();
 FILLCELL_X32 FILLER_266_1848 ();
 FILLCELL_X8 FILLER_266_1880 ();
 FILLCELL_X4 FILLER_266_1888 ();
 FILLCELL_X2 FILLER_266_1892 ();
 FILLCELL_X32 FILLER_266_1895 ();
 FILLCELL_X32 FILLER_266_1927 ();
 FILLCELL_X32 FILLER_266_1959 ();
 FILLCELL_X32 FILLER_266_1991 ();
 FILLCELL_X32 FILLER_266_2023 ();
 FILLCELL_X32 FILLER_266_2055 ();
 FILLCELL_X32 FILLER_266_2087 ();
 FILLCELL_X32 FILLER_266_2119 ();
 FILLCELL_X32 FILLER_266_2151 ();
 FILLCELL_X32 FILLER_266_2183 ();
 FILLCELL_X32 FILLER_266_2215 ();
 FILLCELL_X32 FILLER_266_2247 ();
 FILLCELL_X32 FILLER_266_2279 ();
 FILLCELL_X32 FILLER_266_2311 ();
 FILLCELL_X32 FILLER_266_2343 ();
 FILLCELL_X32 FILLER_266_2375 ();
 FILLCELL_X16 FILLER_266_2407 ();
 FILLCELL_X8 FILLER_266_2423 ();
 FILLCELL_X4 FILLER_266_2431 ();
 FILLCELL_X1 FILLER_266_2435 ();
 FILLCELL_X32 FILLER_267_1 ();
 FILLCELL_X32 FILLER_267_33 ();
 FILLCELL_X32 FILLER_267_65 ();
 FILLCELL_X32 FILLER_267_97 ();
 FILLCELL_X32 FILLER_267_129 ();
 FILLCELL_X32 FILLER_267_161 ();
 FILLCELL_X32 FILLER_267_193 ();
 FILLCELL_X32 FILLER_267_225 ();
 FILLCELL_X32 FILLER_267_257 ();
 FILLCELL_X32 FILLER_267_289 ();
 FILLCELL_X32 FILLER_267_321 ();
 FILLCELL_X32 FILLER_267_353 ();
 FILLCELL_X32 FILLER_267_385 ();
 FILLCELL_X32 FILLER_267_417 ();
 FILLCELL_X32 FILLER_267_449 ();
 FILLCELL_X32 FILLER_267_481 ();
 FILLCELL_X32 FILLER_267_513 ();
 FILLCELL_X32 FILLER_267_545 ();
 FILLCELL_X32 FILLER_267_577 ();
 FILLCELL_X32 FILLER_267_609 ();
 FILLCELL_X32 FILLER_267_641 ();
 FILLCELL_X32 FILLER_267_673 ();
 FILLCELL_X32 FILLER_267_705 ();
 FILLCELL_X32 FILLER_267_737 ();
 FILLCELL_X32 FILLER_267_769 ();
 FILLCELL_X32 FILLER_267_801 ();
 FILLCELL_X32 FILLER_267_833 ();
 FILLCELL_X32 FILLER_267_865 ();
 FILLCELL_X32 FILLER_267_897 ();
 FILLCELL_X32 FILLER_267_929 ();
 FILLCELL_X32 FILLER_267_961 ();
 FILLCELL_X32 FILLER_267_993 ();
 FILLCELL_X32 FILLER_267_1025 ();
 FILLCELL_X32 FILLER_267_1057 ();
 FILLCELL_X32 FILLER_267_1089 ();
 FILLCELL_X32 FILLER_267_1121 ();
 FILLCELL_X32 FILLER_267_1153 ();
 FILLCELL_X32 FILLER_267_1185 ();
 FILLCELL_X32 FILLER_267_1217 ();
 FILLCELL_X8 FILLER_267_1249 ();
 FILLCELL_X4 FILLER_267_1257 ();
 FILLCELL_X2 FILLER_267_1261 ();
 FILLCELL_X32 FILLER_267_1264 ();
 FILLCELL_X32 FILLER_267_1296 ();
 FILLCELL_X32 FILLER_267_1328 ();
 FILLCELL_X32 FILLER_267_1360 ();
 FILLCELL_X32 FILLER_267_1392 ();
 FILLCELL_X32 FILLER_267_1424 ();
 FILLCELL_X32 FILLER_267_1456 ();
 FILLCELL_X32 FILLER_267_1488 ();
 FILLCELL_X32 FILLER_267_1520 ();
 FILLCELL_X32 FILLER_267_1552 ();
 FILLCELL_X32 FILLER_267_1584 ();
 FILLCELL_X32 FILLER_267_1616 ();
 FILLCELL_X32 FILLER_267_1648 ();
 FILLCELL_X32 FILLER_267_1680 ();
 FILLCELL_X32 FILLER_267_1712 ();
 FILLCELL_X32 FILLER_267_1744 ();
 FILLCELL_X32 FILLER_267_1776 ();
 FILLCELL_X32 FILLER_267_1808 ();
 FILLCELL_X32 FILLER_267_1840 ();
 FILLCELL_X32 FILLER_267_1872 ();
 FILLCELL_X32 FILLER_267_1904 ();
 FILLCELL_X32 FILLER_267_1936 ();
 FILLCELL_X32 FILLER_267_1968 ();
 FILLCELL_X32 FILLER_267_2000 ();
 FILLCELL_X32 FILLER_267_2032 ();
 FILLCELL_X32 FILLER_267_2064 ();
 FILLCELL_X32 FILLER_267_2096 ();
 FILLCELL_X32 FILLER_267_2128 ();
 FILLCELL_X32 FILLER_267_2160 ();
 FILLCELL_X32 FILLER_267_2192 ();
 FILLCELL_X32 FILLER_267_2224 ();
 FILLCELL_X32 FILLER_267_2256 ();
 FILLCELL_X32 FILLER_267_2288 ();
 FILLCELL_X32 FILLER_267_2320 ();
 FILLCELL_X32 FILLER_267_2352 ();
 FILLCELL_X32 FILLER_267_2384 ();
 FILLCELL_X16 FILLER_267_2416 ();
 FILLCELL_X4 FILLER_267_2432 ();
 FILLCELL_X32 FILLER_268_1 ();
 FILLCELL_X32 FILLER_268_33 ();
 FILLCELL_X32 FILLER_268_65 ();
 FILLCELL_X32 FILLER_268_97 ();
 FILLCELL_X32 FILLER_268_129 ();
 FILLCELL_X32 FILLER_268_161 ();
 FILLCELL_X32 FILLER_268_193 ();
 FILLCELL_X32 FILLER_268_225 ();
 FILLCELL_X32 FILLER_268_257 ();
 FILLCELL_X32 FILLER_268_289 ();
 FILLCELL_X32 FILLER_268_321 ();
 FILLCELL_X32 FILLER_268_353 ();
 FILLCELL_X32 FILLER_268_385 ();
 FILLCELL_X32 FILLER_268_417 ();
 FILLCELL_X32 FILLER_268_449 ();
 FILLCELL_X32 FILLER_268_481 ();
 FILLCELL_X32 FILLER_268_513 ();
 FILLCELL_X32 FILLER_268_545 ();
 FILLCELL_X32 FILLER_268_577 ();
 FILLCELL_X16 FILLER_268_609 ();
 FILLCELL_X4 FILLER_268_625 ();
 FILLCELL_X2 FILLER_268_629 ();
 FILLCELL_X32 FILLER_268_632 ();
 FILLCELL_X32 FILLER_268_664 ();
 FILLCELL_X32 FILLER_268_696 ();
 FILLCELL_X32 FILLER_268_728 ();
 FILLCELL_X32 FILLER_268_760 ();
 FILLCELL_X32 FILLER_268_792 ();
 FILLCELL_X32 FILLER_268_824 ();
 FILLCELL_X32 FILLER_268_856 ();
 FILLCELL_X32 FILLER_268_888 ();
 FILLCELL_X32 FILLER_268_920 ();
 FILLCELL_X32 FILLER_268_952 ();
 FILLCELL_X32 FILLER_268_984 ();
 FILLCELL_X32 FILLER_268_1016 ();
 FILLCELL_X32 FILLER_268_1048 ();
 FILLCELL_X32 FILLER_268_1080 ();
 FILLCELL_X32 FILLER_268_1112 ();
 FILLCELL_X32 FILLER_268_1144 ();
 FILLCELL_X32 FILLER_268_1176 ();
 FILLCELL_X32 FILLER_268_1208 ();
 FILLCELL_X32 FILLER_268_1240 ();
 FILLCELL_X32 FILLER_268_1272 ();
 FILLCELL_X32 FILLER_268_1304 ();
 FILLCELL_X32 FILLER_268_1336 ();
 FILLCELL_X32 FILLER_268_1368 ();
 FILLCELL_X32 FILLER_268_1400 ();
 FILLCELL_X32 FILLER_268_1432 ();
 FILLCELL_X32 FILLER_268_1464 ();
 FILLCELL_X32 FILLER_268_1496 ();
 FILLCELL_X32 FILLER_268_1528 ();
 FILLCELL_X32 FILLER_268_1560 ();
 FILLCELL_X32 FILLER_268_1592 ();
 FILLCELL_X32 FILLER_268_1624 ();
 FILLCELL_X32 FILLER_268_1656 ();
 FILLCELL_X32 FILLER_268_1688 ();
 FILLCELL_X32 FILLER_268_1720 ();
 FILLCELL_X32 FILLER_268_1752 ();
 FILLCELL_X32 FILLER_268_1784 ();
 FILLCELL_X32 FILLER_268_1816 ();
 FILLCELL_X32 FILLER_268_1848 ();
 FILLCELL_X8 FILLER_268_1880 ();
 FILLCELL_X4 FILLER_268_1888 ();
 FILLCELL_X2 FILLER_268_1892 ();
 FILLCELL_X32 FILLER_268_1895 ();
 FILLCELL_X32 FILLER_268_1927 ();
 FILLCELL_X32 FILLER_268_1959 ();
 FILLCELL_X32 FILLER_268_1991 ();
 FILLCELL_X32 FILLER_268_2023 ();
 FILLCELL_X32 FILLER_268_2055 ();
 FILLCELL_X32 FILLER_268_2087 ();
 FILLCELL_X32 FILLER_268_2119 ();
 FILLCELL_X32 FILLER_268_2151 ();
 FILLCELL_X32 FILLER_268_2183 ();
 FILLCELL_X32 FILLER_268_2215 ();
 FILLCELL_X32 FILLER_268_2247 ();
 FILLCELL_X32 FILLER_268_2279 ();
 FILLCELL_X32 FILLER_268_2311 ();
 FILLCELL_X32 FILLER_268_2343 ();
 FILLCELL_X32 FILLER_268_2375 ();
 FILLCELL_X16 FILLER_268_2407 ();
 FILLCELL_X8 FILLER_268_2423 ();
 FILLCELL_X4 FILLER_268_2431 ();
 FILLCELL_X1 FILLER_268_2435 ();
 FILLCELL_X32 FILLER_269_1 ();
 FILLCELL_X32 FILLER_269_33 ();
 FILLCELL_X32 FILLER_269_65 ();
 FILLCELL_X32 FILLER_269_97 ();
 FILLCELL_X32 FILLER_269_129 ();
 FILLCELL_X32 FILLER_269_161 ();
 FILLCELL_X32 FILLER_269_193 ();
 FILLCELL_X32 FILLER_269_225 ();
 FILLCELL_X32 FILLER_269_257 ();
 FILLCELL_X32 FILLER_269_289 ();
 FILLCELL_X32 FILLER_269_321 ();
 FILLCELL_X32 FILLER_269_353 ();
 FILLCELL_X32 FILLER_269_385 ();
 FILLCELL_X32 FILLER_269_417 ();
 FILLCELL_X32 FILLER_269_449 ();
 FILLCELL_X32 FILLER_269_481 ();
 FILLCELL_X32 FILLER_269_513 ();
 FILLCELL_X32 FILLER_269_545 ();
 FILLCELL_X32 FILLER_269_577 ();
 FILLCELL_X32 FILLER_269_609 ();
 FILLCELL_X32 FILLER_269_641 ();
 FILLCELL_X32 FILLER_269_673 ();
 FILLCELL_X32 FILLER_269_705 ();
 FILLCELL_X32 FILLER_269_737 ();
 FILLCELL_X32 FILLER_269_769 ();
 FILLCELL_X32 FILLER_269_801 ();
 FILLCELL_X32 FILLER_269_833 ();
 FILLCELL_X32 FILLER_269_865 ();
 FILLCELL_X32 FILLER_269_897 ();
 FILLCELL_X32 FILLER_269_929 ();
 FILLCELL_X32 FILLER_269_961 ();
 FILLCELL_X32 FILLER_269_993 ();
 FILLCELL_X32 FILLER_269_1025 ();
 FILLCELL_X32 FILLER_269_1057 ();
 FILLCELL_X32 FILLER_269_1089 ();
 FILLCELL_X32 FILLER_269_1121 ();
 FILLCELL_X32 FILLER_269_1153 ();
 FILLCELL_X32 FILLER_269_1185 ();
 FILLCELL_X32 FILLER_269_1217 ();
 FILLCELL_X8 FILLER_269_1249 ();
 FILLCELL_X4 FILLER_269_1257 ();
 FILLCELL_X2 FILLER_269_1261 ();
 FILLCELL_X32 FILLER_269_1264 ();
 FILLCELL_X32 FILLER_269_1296 ();
 FILLCELL_X32 FILLER_269_1328 ();
 FILLCELL_X32 FILLER_269_1360 ();
 FILLCELL_X32 FILLER_269_1392 ();
 FILLCELL_X32 FILLER_269_1424 ();
 FILLCELL_X32 FILLER_269_1456 ();
 FILLCELL_X32 FILLER_269_1488 ();
 FILLCELL_X32 FILLER_269_1520 ();
 FILLCELL_X32 FILLER_269_1552 ();
 FILLCELL_X32 FILLER_269_1584 ();
 FILLCELL_X32 FILLER_269_1616 ();
 FILLCELL_X32 FILLER_269_1648 ();
 FILLCELL_X32 FILLER_269_1680 ();
 FILLCELL_X32 FILLER_269_1712 ();
 FILLCELL_X32 FILLER_269_1744 ();
 FILLCELL_X32 FILLER_269_1776 ();
 FILLCELL_X32 FILLER_269_1808 ();
 FILLCELL_X32 FILLER_269_1840 ();
 FILLCELL_X32 FILLER_269_1872 ();
 FILLCELL_X32 FILLER_269_1904 ();
 FILLCELL_X32 FILLER_269_1936 ();
 FILLCELL_X32 FILLER_269_1968 ();
 FILLCELL_X32 FILLER_269_2000 ();
 FILLCELL_X32 FILLER_269_2032 ();
 FILLCELL_X32 FILLER_269_2064 ();
 FILLCELL_X32 FILLER_269_2096 ();
 FILLCELL_X32 FILLER_269_2128 ();
 FILLCELL_X32 FILLER_269_2160 ();
 FILLCELL_X32 FILLER_269_2192 ();
 FILLCELL_X32 FILLER_269_2224 ();
 FILLCELL_X32 FILLER_269_2256 ();
 FILLCELL_X32 FILLER_269_2288 ();
 FILLCELL_X32 FILLER_269_2320 ();
 FILLCELL_X32 FILLER_269_2352 ();
 FILLCELL_X32 FILLER_269_2384 ();
 FILLCELL_X16 FILLER_269_2416 ();
 FILLCELL_X4 FILLER_269_2432 ();
 FILLCELL_X32 FILLER_270_1 ();
 FILLCELL_X32 FILLER_270_33 ();
 FILLCELL_X32 FILLER_270_65 ();
 FILLCELL_X32 FILLER_270_97 ();
 FILLCELL_X32 FILLER_270_129 ();
 FILLCELL_X32 FILLER_270_161 ();
 FILLCELL_X32 FILLER_270_193 ();
 FILLCELL_X32 FILLER_270_225 ();
 FILLCELL_X32 FILLER_270_257 ();
 FILLCELL_X32 FILLER_270_289 ();
 FILLCELL_X32 FILLER_270_321 ();
 FILLCELL_X32 FILLER_270_353 ();
 FILLCELL_X32 FILLER_270_385 ();
 FILLCELL_X32 FILLER_270_417 ();
 FILLCELL_X32 FILLER_270_449 ();
 FILLCELL_X32 FILLER_270_481 ();
 FILLCELL_X32 FILLER_270_513 ();
 FILLCELL_X32 FILLER_270_545 ();
 FILLCELL_X32 FILLER_270_577 ();
 FILLCELL_X16 FILLER_270_609 ();
 FILLCELL_X4 FILLER_270_625 ();
 FILLCELL_X2 FILLER_270_629 ();
 FILLCELL_X32 FILLER_270_632 ();
 FILLCELL_X32 FILLER_270_664 ();
 FILLCELL_X32 FILLER_270_696 ();
 FILLCELL_X32 FILLER_270_728 ();
 FILLCELL_X32 FILLER_270_760 ();
 FILLCELL_X32 FILLER_270_792 ();
 FILLCELL_X32 FILLER_270_824 ();
 FILLCELL_X32 FILLER_270_856 ();
 FILLCELL_X32 FILLER_270_888 ();
 FILLCELL_X32 FILLER_270_920 ();
 FILLCELL_X32 FILLER_270_952 ();
 FILLCELL_X32 FILLER_270_984 ();
 FILLCELL_X32 FILLER_270_1016 ();
 FILLCELL_X32 FILLER_270_1048 ();
 FILLCELL_X32 FILLER_270_1080 ();
 FILLCELL_X32 FILLER_270_1112 ();
 FILLCELL_X32 FILLER_270_1144 ();
 FILLCELL_X32 FILLER_270_1176 ();
 FILLCELL_X32 FILLER_270_1208 ();
 FILLCELL_X32 FILLER_270_1240 ();
 FILLCELL_X32 FILLER_270_1272 ();
 FILLCELL_X32 FILLER_270_1304 ();
 FILLCELL_X32 FILLER_270_1336 ();
 FILLCELL_X32 FILLER_270_1368 ();
 FILLCELL_X32 FILLER_270_1400 ();
 FILLCELL_X32 FILLER_270_1432 ();
 FILLCELL_X32 FILLER_270_1464 ();
 FILLCELL_X32 FILLER_270_1496 ();
 FILLCELL_X32 FILLER_270_1528 ();
 FILLCELL_X32 FILLER_270_1560 ();
 FILLCELL_X32 FILLER_270_1592 ();
 FILLCELL_X32 FILLER_270_1624 ();
 FILLCELL_X32 FILLER_270_1656 ();
 FILLCELL_X32 FILLER_270_1688 ();
 FILLCELL_X32 FILLER_270_1720 ();
 FILLCELL_X32 FILLER_270_1752 ();
 FILLCELL_X32 FILLER_270_1784 ();
 FILLCELL_X32 FILLER_270_1816 ();
 FILLCELL_X32 FILLER_270_1848 ();
 FILLCELL_X8 FILLER_270_1880 ();
 FILLCELL_X4 FILLER_270_1888 ();
 FILLCELL_X2 FILLER_270_1892 ();
 FILLCELL_X32 FILLER_270_1895 ();
 FILLCELL_X32 FILLER_270_1927 ();
 FILLCELL_X32 FILLER_270_1959 ();
 FILLCELL_X32 FILLER_270_1991 ();
 FILLCELL_X32 FILLER_270_2023 ();
 FILLCELL_X32 FILLER_270_2055 ();
 FILLCELL_X32 FILLER_270_2087 ();
 FILLCELL_X32 FILLER_270_2119 ();
 FILLCELL_X32 FILLER_270_2151 ();
 FILLCELL_X32 FILLER_270_2183 ();
 FILLCELL_X32 FILLER_270_2215 ();
 FILLCELL_X32 FILLER_270_2247 ();
 FILLCELL_X32 FILLER_270_2279 ();
 FILLCELL_X32 FILLER_270_2311 ();
 FILLCELL_X32 FILLER_270_2343 ();
 FILLCELL_X32 FILLER_270_2375 ();
 FILLCELL_X16 FILLER_270_2407 ();
 FILLCELL_X8 FILLER_270_2423 ();
 FILLCELL_X4 FILLER_270_2431 ();
 FILLCELL_X1 FILLER_270_2435 ();
 FILLCELL_X32 FILLER_271_1 ();
 FILLCELL_X32 FILLER_271_33 ();
 FILLCELL_X32 FILLER_271_65 ();
 FILLCELL_X32 FILLER_271_97 ();
 FILLCELL_X32 FILLER_271_129 ();
 FILLCELL_X32 FILLER_271_161 ();
 FILLCELL_X32 FILLER_271_193 ();
 FILLCELL_X32 FILLER_271_225 ();
 FILLCELL_X32 FILLER_271_257 ();
 FILLCELL_X32 FILLER_271_289 ();
 FILLCELL_X32 FILLER_271_321 ();
 FILLCELL_X32 FILLER_271_353 ();
 FILLCELL_X32 FILLER_271_385 ();
 FILLCELL_X32 FILLER_271_417 ();
 FILLCELL_X32 FILLER_271_449 ();
 FILLCELL_X32 FILLER_271_481 ();
 FILLCELL_X32 FILLER_271_513 ();
 FILLCELL_X32 FILLER_271_545 ();
 FILLCELL_X32 FILLER_271_577 ();
 FILLCELL_X32 FILLER_271_609 ();
 FILLCELL_X32 FILLER_271_641 ();
 FILLCELL_X32 FILLER_271_673 ();
 FILLCELL_X32 FILLER_271_705 ();
 FILLCELL_X32 FILLER_271_737 ();
 FILLCELL_X32 FILLER_271_769 ();
 FILLCELL_X32 FILLER_271_801 ();
 FILLCELL_X32 FILLER_271_833 ();
 FILLCELL_X32 FILLER_271_865 ();
 FILLCELL_X32 FILLER_271_897 ();
 FILLCELL_X32 FILLER_271_929 ();
 FILLCELL_X32 FILLER_271_961 ();
 FILLCELL_X32 FILLER_271_993 ();
 FILLCELL_X32 FILLER_271_1025 ();
 FILLCELL_X32 FILLER_271_1057 ();
 FILLCELL_X32 FILLER_271_1089 ();
 FILLCELL_X32 FILLER_271_1121 ();
 FILLCELL_X32 FILLER_271_1153 ();
 FILLCELL_X32 FILLER_271_1185 ();
 FILLCELL_X32 FILLER_271_1217 ();
 FILLCELL_X8 FILLER_271_1249 ();
 FILLCELL_X4 FILLER_271_1257 ();
 FILLCELL_X2 FILLER_271_1261 ();
 FILLCELL_X32 FILLER_271_1264 ();
 FILLCELL_X32 FILLER_271_1296 ();
 FILLCELL_X32 FILLER_271_1328 ();
 FILLCELL_X32 FILLER_271_1360 ();
 FILLCELL_X32 FILLER_271_1392 ();
 FILLCELL_X32 FILLER_271_1424 ();
 FILLCELL_X32 FILLER_271_1456 ();
 FILLCELL_X32 FILLER_271_1488 ();
 FILLCELL_X32 FILLER_271_1520 ();
 FILLCELL_X32 FILLER_271_1552 ();
 FILLCELL_X32 FILLER_271_1584 ();
 FILLCELL_X32 FILLER_271_1616 ();
 FILLCELL_X32 FILLER_271_1648 ();
 FILLCELL_X32 FILLER_271_1680 ();
 FILLCELL_X32 FILLER_271_1712 ();
 FILLCELL_X32 FILLER_271_1744 ();
 FILLCELL_X32 FILLER_271_1776 ();
 FILLCELL_X32 FILLER_271_1808 ();
 FILLCELL_X32 FILLER_271_1840 ();
 FILLCELL_X32 FILLER_271_1872 ();
 FILLCELL_X32 FILLER_271_1904 ();
 FILLCELL_X32 FILLER_271_1936 ();
 FILLCELL_X32 FILLER_271_1968 ();
 FILLCELL_X32 FILLER_271_2000 ();
 FILLCELL_X32 FILLER_271_2032 ();
 FILLCELL_X32 FILLER_271_2064 ();
 FILLCELL_X32 FILLER_271_2096 ();
 FILLCELL_X32 FILLER_271_2128 ();
 FILLCELL_X32 FILLER_271_2160 ();
 FILLCELL_X32 FILLER_271_2192 ();
 FILLCELL_X32 FILLER_271_2224 ();
 FILLCELL_X32 FILLER_271_2256 ();
 FILLCELL_X32 FILLER_271_2288 ();
 FILLCELL_X32 FILLER_271_2320 ();
 FILLCELL_X32 FILLER_271_2352 ();
 FILLCELL_X32 FILLER_271_2384 ();
 FILLCELL_X16 FILLER_271_2416 ();
 FILLCELL_X4 FILLER_271_2432 ();
 FILLCELL_X32 FILLER_272_1 ();
 FILLCELL_X32 FILLER_272_33 ();
 FILLCELL_X32 FILLER_272_65 ();
 FILLCELL_X32 FILLER_272_97 ();
 FILLCELL_X32 FILLER_272_129 ();
 FILLCELL_X32 FILLER_272_161 ();
 FILLCELL_X32 FILLER_272_193 ();
 FILLCELL_X32 FILLER_272_225 ();
 FILLCELL_X32 FILLER_272_257 ();
 FILLCELL_X32 FILLER_272_289 ();
 FILLCELL_X32 FILLER_272_321 ();
 FILLCELL_X32 FILLER_272_353 ();
 FILLCELL_X32 FILLER_272_385 ();
 FILLCELL_X32 FILLER_272_417 ();
 FILLCELL_X32 FILLER_272_449 ();
 FILLCELL_X32 FILLER_272_481 ();
 FILLCELL_X32 FILLER_272_513 ();
 FILLCELL_X32 FILLER_272_545 ();
 FILLCELL_X32 FILLER_272_577 ();
 FILLCELL_X16 FILLER_272_609 ();
 FILLCELL_X4 FILLER_272_625 ();
 FILLCELL_X2 FILLER_272_629 ();
 FILLCELL_X32 FILLER_272_632 ();
 FILLCELL_X32 FILLER_272_664 ();
 FILLCELL_X32 FILLER_272_696 ();
 FILLCELL_X32 FILLER_272_728 ();
 FILLCELL_X32 FILLER_272_760 ();
 FILLCELL_X32 FILLER_272_792 ();
 FILLCELL_X32 FILLER_272_824 ();
 FILLCELL_X32 FILLER_272_856 ();
 FILLCELL_X32 FILLER_272_888 ();
 FILLCELL_X32 FILLER_272_920 ();
 FILLCELL_X32 FILLER_272_952 ();
 FILLCELL_X32 FILLER_272_984 ();
 FILLCELL_X32 FILLER_272_1016 ();
 FILLCELL_X32 FILLER_272_1048 ();
 FILLCELL_X32 FILLER_272_1080 ();
 FILLCELL_X32 FILLER_272_1112 ();
 FILLCELL_X32 FILLER_272_1144 ();
 FILLCELL_X32 FILLER_272_1176 ();
 FILLCELL_X32 FILLER_272_1208 ();
 FILLCELL_X32 FILLER_272_1240 ();
 FILLCELL_X32 FILLER_272_1272 ();
 FILLCELL_X32 FILLER_272_1304 ();
 FILLCELL_X32 FILLER_272_1336 ();
 FILLCELL_X32 FILLER_272_1368 ();
 FILLCELL_X32 FILLER_272_1400 ();
 FILLCELL_X32 FILLER_272_1432 ();
 FILLCELL_X32 FILLER_272_1464 ();
 FILLCELL_X32 FILLER_272_1496 ();
 FILLCELL_X32 FILLER_272_1528 ();
 FILLCELL_X32 FILLER_272_1560 ();
 FILLCELL_X32 FILLER_272_1592 ();
 FILLCELL_X32 FILLER_272_1624 ();
 FILLCELL_X32 FILLER_272_1656 ();
 FILLCELL_X32 FILLER_272_1688 ();
 FILLCELL_X32 FILLER_272_1720 ();
 FILLCELL_X32 FILLER_272_1752 ();
 FILLCELL_X32 FILLER_272_1784 ();
 FILLCELL_X32 FILLER_272_1816 ();
 FILLCELL_X32 FILLER_272_1848 ();
 FILLCELL_X8 FILLER_272_1880 ();
 FILLCELL_X4 FILLER_272_1888 ();
 FILLCELL_X2 FILLER_272_1892 ();
 FILLCELL_X32 FILLER_272_1895 ();
 FILLCELL_X32 FILLER_272_1927 ();
 FILLCELL_X32 FILLER_272_1959 ();
 FILLCELL_X32 FILLER_272_1991 ();
 FILLCELL_X32 FILLER_272_2023 ();
 FILLCELL_X32 FILLER_272_2055 ();
 FILLCELL_X32 FILLER_272_2087 ();
 FILLCELL_X32 FILLER_272_2119 ();
 FILLCELL_X32 FILLER_272_2151 ();
 FILLCELL_X32 FILLER_272_2183 ();
 FILLCELL_X32 FILLER_272_2215 ();
 FILLCELL_X32 FILLER_272_2247 ();
 FILLCELL_X32 FILLER_272_2279 ();
 FILLCELL_X32 FILLER_272_2311 ();
 FILLCELL_X32 FILLER_272_2343 ();
 FILLCELL_X32 FILLER_272_2375 ();
 FILLCELL_X16 FILLER_272_2407 ();
 FILLCELL_X8 FILLER_272_2423 ();
 FILLCELL_X4 FILLER_272_2431 ();
 FILLCELL_X1 FILLER_272_2435 ();
 FILLCELL_X32 FILLER_273_1 ();
 FILLCELL_X32 FILLER_273_33 ();
 FILLCELL_X32 FILLER_273_65 ();
 FILLCELL_X32 FILLER_273_97 ();
 FILLCELL_X32 FILLER_273_129 ();
 FILLCELL_X32 FILLER_273_161 ();
 FILLCELL_X32 FILLER_273_193 ();
 FILLCELL_X32 FILLER_273_225 ();
 FILLCELL_X32 FILLER_273_257 ();
 FILLCELL_X32 FILLER_273_289 ();
 FILLCELL_X32 FILLER_273_321 ();
 FILLCELL_X32 FILLER_273_353 ();
 FILLCELL_X32 FILLER_273_385 ();
 FILLCELL_X32 FILLER_273_417 ();
 FILLCELL_X32 FILLER_273_449 ();
 FILLCELL_X32 FILLER_273_481 ();
 FILLCELL_X32 FILLER_273_513 ();
 FILLCELL_X32 FILLER_273_545 ();
 FILLCELL_X32 FILLER_273_577 ();
 FILLCELL_X32 FILLER_273_609 ();
 FILLCELL_X32 FILLER_273_641 ();
 FILLCELL_X32 FILLER_273_673 ();
 FILLCELL_X32 FILLER_273_705 ();
 FILLCELL_X32 FILLER_273_737 ();
 FILLCELL_X32 FILLER_273_769 ();
 FILLCELL_X32 FILLER_273_801 ();
 FILLCELL_X32 FILLER_273_833 ();
 FILLCELL_X32 FILLER_273_865 ();
 FILLCELL_X32 FILLER_273_897 ();
 FILLCELL_X32 FILLER_273_929 ();
 FILLCELL_X32 FILLER_273_961 ();
 FILLCELL_X32 FILLER_273_993 ();
 FILLCELL_X32 FILLER_273_1025 ();
 FILLCELL_X32 FILLER_273_1057 ();
 FILLCELL_X32 FILLER_273_1089 ();
 FILLCELL_X32 FILLER_273_1121 ();
 FILLCELL_X32 FILLER_273_1153 ();
 FILLCELL_X32 FILLER_273_1185 ();
 FILLCELL_X32 FILLER_273_1217 ();
 FILLCELL_X8 FILLER_273_1249 ();
 FILLCELL_X4 FILLER_273_1257 ();
 FILLCELL_X2 FILLER_273_1261 ();
 FILLCELL_X32 FILLER_273_1264 ();
 FILLCELL_X32 FILLER_273_1296 ();
 FILLCELL_X32 FILLER_273_1328 ();
 FILLCELL_X32 FILLER_273_1360 ();
 FILLCELL_X32 FILLER_273_1392 ();
 FILLCELL_X32 FILLER_273_1424 ();
 FILLCELL_X32 FILLER_273_1456 ();
 FILLCELL_X32 FILLER_273_1488 ();
 FILLCELL_X32 FILLER_273_1520 ();
 FILLCELL_X32 FILLER_273_1552 ();
 FILLCELL_X32 FILLER_273_1584 ();
 FILLCELL_X32 FILLER_273_1616 ();
 FILLCELL_X32 FILLER_273_1648 ();
 FILLCELL_X32 FILLER_273_1680 ();
 FILLCELL_X32 FILLER_273_1712 ();
 FILLCELL_X32 FILLER_273_1744 ();
 FILLCELL_X32 FILLER_273_1776 ();
 FILLCELL_X32 FILLER_273_1808 ();
 FILLCELL_X32 FILLER_273_1840 ();
 FILLCELL_X32 FILLER_273_1872 ();
 FILLCELL_X32 FILLER_273_1904 ();
 FILLCELL_X32 FILLER_273_1936 ();
 FILLCELL_X32 FILLER_273_1968 ();
 FILLCELL_X32 FILLER_273_2000 ();
 FILLCELL_X32 FILLER_273_2032 ();
 FILLCELL_X32 FILLER_273_2064 ();
 FILLCELL_X32 FILLER_273_2096 ();
 FILLCELL_X32 FILLER_273_2128 ();
 FILLCELL_X32 FILLER_273_2160 ();
 FILLCELL_X32 FILLER_273_2192 ();
 FILLCELL_X32 FILLER_273_2224 ();
 FILLCELL_X32 FILLER_273_2256 ();
 FILLCELL_X32 FILLER_273_2288 ();
 FILLCELL_X32 FILLER_273_2320 ();
 FILLCELL_X32 FILLER_273_2352 ();
 FILLCELL_X32 FILLER_273_2384 ();
 FILLCELL_X16 FILLER_273_2416 ();
 FILLCELL_X4 FILLER_273_2432 ();
 FILLCELL_X32 FILLER_274_1 ();
 FILLCELL_X32 FILLER_274_33 ();
 FILLCELL_X32 FILLER_274_65 ();
 FILLCELL_X32 FILLER_274_97 ();
 FILLCELL_X32 FILLER_274_129 ();
 FILLCELL_X32 FILLER_274_161 ();
 FILLCELL_X32 FILLER_274_193 ();
 FILLCELL_X32 FILLER_274_225 ();
 FILLCELL_X32 FILLER_274_257 ();
 FILLCELL_X32 FILLER_274_289 ();
 FILLCELL_X32 FILLER_274_321 ();
 FILLCELL_X32 FILLER_274_353 ();
 FILLCELL_X32 FILLER_274_385 ();
 FILLCELL_X32 FILLER_274_417 ();
 FILLCELL_X32 FILLER_274_449 ();
 FILLCELL_X32 FILLER_274_481 ();
 FILLCELL_X32 FILLER_274_513 ();
 FILLCELL_X32 FILLER_274_545 ();
 FILLCELL_X32 FILLER_274_577 ();
 FILLCELL_X16 FILLER_274_609 ();
 FILLCELL_X4 FILLER_274_625 ();
 FILLCELL_X2 FILLER_274_629 ();
 FILLCELL_X32 FILLER_274_632 ();
 FILLCELL_X32 FILLER_274_664 ();
 FILLCELL_X32 FILLER_274_696 ();
 FILLCELL_X32 FILLER_274_728 ();
 FILLCELL_X32 FILLER_274_760 ();
 FILLCELL_X32 FILLER_274_792 ();
 FILLCELL_X32 FILLER_274_824 ();
 FILLCELL_X32 FILLER_274_856 ();
 FILLCELL_X32 FILLER_274_888 ();
 FILLCELL_X32 FILLER_274_920 ();
 FILLCELL_X32 FILLER_274_952 ();
 FILLCELL_X32 FILLER_274_984 ();
 FILLCELL_X32 FILLER_274_1016 ();
 FILLCELL_X32 FILLER_274_1048 ();
 FILLCELL_X32 FILLER_274_1080 ();
 FILLCELL_X32 FILLER_274_1112 ();
 FILLCELL_X32 FILLER_274_1144 ();
 FILLCELL_X32 FILLER_274_1176 ();
 FILLCELL_X32 FILLER_274_1208 ();
 FILLCELL_X32 FILLER_274_1240 ();
 FILLCELL_X32 FILLER_274_1272 ();
 FILLCELL_X32 FILLER_274_1304 ();
 FILLCELL_X32 FILLER_274_1336 ();
 FILLCELL_X32 FILLER_274_1368 ();
 FILLCELL_X32 FILLER_274_1400 ();
 FILLCELL_X32 FILLER_274_1432 ();
 FILLCELL_X32 FILLER_274_1464 ();
 FILLCELL_X32 FILLER_274_1496 ();
 FILLCELL_X32 FILLER_274_1528 ();
 FILLCELL_X32 FILLER_274_1560 ();
 FILLCELL_X32 FILLER_274_1592 ();
 FILLCELL_X32 FILLER_274_1624 ();
 FILLCELL_X32 FILLER_274_1656 ();
 FILLCELL_X32 FILLER_274_1688 ();
 FILLCELL_X32 FILLER_274_1720 ();
 FILLCELL_X32 FILLER_274_1752 ();
 FILLCELL_X32 FILLER_274_1784 ();
 FILLCELL_X32 FILLER_274_1816 ();
 FILLCELL_X32 FILLER_274_1848 ();
 FILLCELL_X8 FILLER_274_1880 ();
 FILLCELL_X4 FILLER_274_1888 ();
 FILLCELL_X2 FILLER_274_1892 ();
 FILLCELL_X32 FILLER_274_1895 ();
 FILLCELL_X32 FILLER_274_1927 ();
 FILLCELL_X32 FILLER_274_1959 ();
 FILLCELL_X32 FILLER_274_1991 ();
 FILLCELL_X32 FILLER_274_2023 ();
 FILLCELL_X32 FILLER_274_2055 ();
 FILLCELL_X32 FILLER_274_2087 ();
 FILLCELL_X32 FILLER_274_2119 ();
 FILLCELL_X32 FILLER_274_2151 ();
 FILLCELL_X32 FILLER_274_2183 ();
 FILLCELL_X32 FILLER_274_2215 ();
 FILLCELL_X32 FILLER_274_2247 ();
 FILLCELL_X32 FILLER_274_2279 ();
 FILLCELL_X32 FILLER_274_2311 ();
 FILLCELL_X32 FILLER_274_2343 ();
 FILLCELL_X32 FILLER_274_2375 ();
 FILLCELL_X16 FILLER_274_2407 ();
 FILLCELL_X8 FILLER_274_2423 ();
 FILLCELL_X4 FILLER_274_2431 ();
 FILLCELL_X1 FILLER_274_2435 ();
 FILLCELL_X32 FILLER_275_1 ();
 FILLCELL_X32 FILLER_275_33 ();
 FILLCELL_X32 FILLER_275_65 ();
 FILLCELL_X32 FILLER_275_97 ();
 FILLCELL_X32 FILLER_275_129 ();
 FILLCELL_X32 FILLER_275_161 ();
 FILLCELL_X32 FILLER_275_193 ();
 FILLCELL_X32 FILLER_275_225 ();
 FILLCELL_X32 FILLER_275_257 ();
 FILLCELL_X32 FILLER_275_289 ();
 FILLCELL_X32 FILLER_275_321 ();
 FILLCELL_X32 FILLER_275_353 ();
 FILLCELL_X32 FILLER_275_385 ();
 FILLCELL_X32 FILLER_275_417 ();
 FILLCELL_X32 FILLER_275_449 ();
 FILLCELL_X32 FILLER_275_481 ();
 FILLCELL_X32 FILLER_275_513 ();
 FILLCELL_X32 FILLER_275_545 ();
 FILLCELL_X32 FILLER_275_577 ();
 FILLCELL_X32 FILLER_275_609 ();
 FILLCELL_X32 FILLER_275_641 ();
 FILLCELL_X32 FILLER_275_673 ();
 FILLCELL_X32 FILLER_275_705 ();
 FILLCELL_X32 FILLER_275_737 ();
 FILLCELL_X32 FILLER_275_769 ();
 FILLCELL_X32 FILLER_275_801 ();
 FILLCELL_X32 FILLER_275_833 ();
 FILLCELL_X32 FILLER_275_865 ();
 FILLCELL_X32 FILLER_275_897 ();
 FILLCELL_X32 FILLER_275_929 ();
 FILLCELL_X32 FILLER_275_961 ();
 FILLCELL_X32 FILLER_275_993 ();
 FILLCELL_X32 FILLER_275_1025 ();
 FILLCELL_X32 FILLER_275_1057 ();
 FILLCELL_X32 FILLER_275_1089 ();
 FILLCELL_X32 FILLER_275_1121 ();
 FILLCELL_X32 FILLER_275_1153 ();
 FILLCELL_X32 FILLER_275_1185 ();
 FILLCELL_X32 FILLER_275_1217 ();
 FILLCELL_X8 FILLER_275_1249 ();
 FILLCELL_X4 FILLER_275_1257 ();
 FILLCELL_X2 FILLER_275_1261 ();
 FILLCELL_X32 FILLER_275_1264 ();
 FILLCELL_X32 FILLER_275_1296 ();
 FILLCELL_X32 FILLER_275_1328 ();
 FILLCELL_X32 FILLER_275_1360 ();
 FILLCELL_X32 FILLER_275_1392 ();
 FILLCELL_X32 FILLER_275_1424 ();
 FILLCELL_X32 FILLER_275_1456 ();
 FILLCELL_X32 FILLER_275_1488 ();
 FILLCELL_X32 FILLER_275_1520 ();
 FILLCELL_X32 FILLER_275_1552 ();
 FILLCELL_X32 FILLER_275_1584 ();
 FILLCELL_X32 FILLER_275_1616 ();
 FILLCELL_X32 FILLER_275_1648 ();
 FILLCELL_X32 FILLER_275_1680 ();
 FILLCELL_X32 FILLER_275_1712 ();
 FILLCELL_X32 FILLER_275_1744 ();
 FILLCELL_X32 FILLER_275_1776 ();
 FILLCELL_X32 FILLER_275_1808 ();
 FILLCELL_X32 FILLER_275_1840 ();
 FILLCELL_X32 FILLER_275_1872 ();
 FILLCELL_X32 FILLER_275_1904 ();
 FILLCELL_X32 FILLER_275_1936 ();
 FILLCELL_X32 FILLER_275_1968 ();
 FILLCELL_X32 FILLER_275_2000 ();
 FILLCELL_X32 FILLER_275_2032 ();
 FILLCELL_X32 FILLER_275_2064 ();
 FILLCELL_X32 FILLER_275_2096 ();
 FILLCELL_X32 FILLER_275_2128 ();
 FILLCELL_X32 FILLER_275_2160 ();
 FILLCELL_X32 FILLER_275_2192 ();
 FILLCELL_X32 FILLER_275_2224 ();
 FILLCELL_X32 FILLER_275_2256 ();
 FILLCELL_X32 FILLER_275_2288 ();
 FILLCELL_X32 FILLER_275_2320 ();
 FILLCELL_X32 FILLER_275_2352 ();
 FILLCELL_X32 FILLER_275_2384 ();
 FILLCELL_X16 FILLER_275_2416 ();
 FILLCELL_X4 FILLER_275_2432 ();
 FILLCELL_X32 FILLER_276_1 ();
 FILLCELL_X32 FILLER_276_33 ();
 FILLCELL_X32 FILLER_276_65 ();
 FILLCELL_X32 FILLER_276_97 ();
 FILLCELL_X32 FILLER_276_129 ();
 FILLCELL_X32 FILLER_276_161 ();
 FILLCELL_X32 FILLER_276_193 ();
 FILLCELL_X32 FILLER_276_225 ();
 FILLCELL_X32 FILLER_276_257 ();
 FILLCELL_X32 FILLER_276_289 ();
 FILLCELL_X32 FILLER_276_321 ();
 FILLCELL_X32 FILLER_276_353 ();
 FILLCELL_X32 FILLER_276_385 ();
 FILLCELL_X32 FILLER_276_417 ();
 FILLCELL_X32 FILLER_276_449 ();
 FILLCELL_X32 FILLER_276_481 ();
 FILLCELL_X32 FILLER_276_513 ();
 FILLCELL_X32 FILLER_276_545 ();
 FILLCELL_X32 FILLER_276_577 ();
 FILLCELL_X16 FILLER_276_609 ();
 FILLCELL_X4 FILLER_276_625 ();
 FILLCELL_X2 FILLER_276_629 ();
 FILLCELL_X32 FILLER_276_632 ();
 FILLCELL_X32 FILLER_276_664 ();
 FILLCELL_X32 FILLER_276_696 ();
 FILLCELL_X32 FILLER_276_728 ();
 FILLCELL_X32 FILLER_276_760 ();
 FILLCELL_X32 FILLER_276_792 ();
 FILLCELL_X32 FILLER_276_824 ();
 FILLCELL_X32 FILLER_276_856 ();
 FILLCELL_X32 FILLER_276_888 ();
 FILLCELL_X32 FILLER_276_920 ();
 FILLCELL_X32 FILLER_276_952 ();
 FILLCELL_X32 FILLER_276_984 ();
 FILLCELL_X32 FILLER_276_1016 ();
 FILLCELL_X32 FILLER_276_1048 ();
 FILLCELL_X32 FILLER_276_1080 ();
 FILLCELL_X32 FILLER_276_1112 ();
 FILLCELL_X32 FILLER_276_1144 ();
 FILLCELL_X32 FILLER_276_1176 ();
 FILLCELL_X32 FILLER_276_1208 ();
 FILLCELL_X32 FILLER_276_1240 ();
 FILLCELL_X32 FILLER_276_1272 ();
 FILLCELL_X32 FILLER_276_1304 ();
 FILLCELL_X32 FILLER_276_1336 ();
 FILLCELL_X32 FILLER_276_1368 ();
 FILLCELL_X32 FILLER_276_1400 ();
 FILLCELL_X32 FILLER_276_1432 ();
 FILLCELL_X32 FILLER_276_1464 ();
 FILLCELL_X32 FILLER_276_1496 ();
 FILLCELL_X32 FILLER_276_1528 ();
 FILLCELL_X32 FILLER_276_1560 ();
 FILLCELL_X32 FILLER_276_1592 ();
 FILLCELL_X32 FILLER_276_1624 ();
 FILLCELL_X32 FILLER_276_1656 ();
 FILLCELL_X32 FILLER_276_1688 ();
 FILLCELL_X32 FILLER_276_1720 ();
 FILLCELL_X32 FILLER_276_1752 ();
 FILLCELL_X32 FILLER_276_1784 ();
 FILLCELL_X32 FILLER_276_1816 ();
 FILLCELL_X32 FILLER_276_1848 ();
 FILLCELL_X8 FILLER_276_1880 ();
 FILLCELL_X4 FILLER_276_1888 ();
 FILLCELL_X2 FILLER_276_1892 ();
 FILLCELL_X32 FILLER_276_1895 ();
 FILLCELL_X32 FILLER_276_1927 ();
 FILLCELL_X32 FILLER_276_1959 ();
 FILLCELL_X32 FILLER_276_1991 ();
 FILLCELL_X32 FILLER_276_2023 ();
 FILLCELL_X32 FILLER_276_2055 ();
 FILLCELL_X32 FILLER_276_2087 ();
 FILLCELL_X32 FILLER_276_2119 ();
 FILLCELL_X32 FILLER_276_2151 ();
 FILLCELL_X32 FILLER_276_2183 ();
 FILLCELL_X32 FILLER_276_2215 ();
 FILLCELL_X32 FILLER_276_2247 ();
 FILLCELL_X32 FILLER_276_2279 ();
 FILLCELL_X32 FILLER_276_2311 ();
 FILLCELL_X32 FILLER_276_2343 ();
 FILLCELL_X32 FILLER_276_2375 ();
 FILLCELL_X16 FILLER_276_2407 ();
 FILLCELL_X8 FILLER_276_2423 ();
 FILLCELL_X4 FILLER_276_2431 ();
 FILLCELL_X1 FILLER_276_2435 ();
 FILLCELL_X32 FILLER_277_1 ();
 FILLCELL_X32 FILLER_277_33 ();
 FILLCELL_X32 FILLER_277_65 ();
 FILLCELL_X32 FILLER_277_97 ();
 FILLCELL_X32 FILLER_277_129 ();
 FILLCELL_X32 FILLER_277_161 ();
 FILLCELL_X32 FILLER_277_193 ();
 FILLCELL_X32 FILLER_277_225 ();
 FILLCELL_X32 FILLER_277_257 ();
 FILLCELL_X32 FILLER_277_289 ();
 FILLCELL_X32 FILLER_277_321 ();
 FILLCELL_X32 FILLER_277_353 ();
 FILLCELL_X32 FILLER_277_385 ();
 FILLCELL_X32 FILLER_277_417 ();
 FILLCELL_X32 FILLER_277_449 ();
 FILLCELL_X32 FILLER_277_481 ();
 FILLCELL_X32 FILLER_277_513 ();
 FILLCELL_X32 FILLER_277_545 ();
 FILLCELL_X32 FILLER_277_577 ();
 FILLCELL_X32 FILLER_277_609 ();
 FILLCELL_X32 FILLER_277_641 ();
 FILLCELL_X32 FILLER_277_673 ();
 FILLCELL_X32 FILLER_277_705 ();
 FILLCELL_X32 FILLER_277_737 ();
 FILLCELL_X32 FILLER_277_769 ();
 FILLCELL_X32 FILLER_277_801 ();
 FILLCELL_X32 FILLER_277_833 ();
 FILLCELL_X32 FILLER_277_865 ();
 FILLCELL_X32 FILLER_277_897 ();
 FILLCELL_X32 FILLER_277_929 ();
 FILLCELL_X32 FILLER_277_961 ();
 FILLCELL_X32 FILLER_277_993 ();
 FILLCELL_X32 FILLER_277_1025 ();
 FILLCELL_X32 FILLER_277_1057 ();
 FILLCELL_X32 FILLER_277_1089 ();
 FILLCELL_X32 FILLER_277_1121 ();
 FILLCELL_X32 FILLER_277_1153 ();
 FILLCELL_X32 FILLER_277_1185 ();
 FILLCELL_X32 FILLER_277_1217 ();
 FILLCELL_X8 FILLER_277_1249 ();
 FILLCELL_X4 FILLER_277_1257 ();
 FILLCELL_X2 FILLER_277_1261 ();
 FILLCELL_X32 FILLER_277_1264 ();
 FILLCELL_X32 FILLER_277_1296 ();
 FILLCELL_X32 FILLER_277_1328 ();
 FILLCELL_X32 FILLER_277_1360 ();
 FILLCELL_X32 FILLER_277_1392 ();
 FILLCELL_X32 FILLER_277_1424 ();
 FILLCELL_X32 FILLER_277_1456 ();
 FILLCELL_X32 FILLER_277_1488 ();
 FILLCELL_X32 FILLER_277_1520 ();
 FILLCELL_X32 FILLER_277_1552 ();
 FILLCELL_X32 FILLER_277_1584 ();
 FILLCELL_X32 FILLER_277_1616 ();
 FILLCELL_X32 FILLER_277_1648 ();
 FILLCELL_X32 FILLER_277_1680 ();
 FILLCELL_X32 FILLER_277_1712 ();
 FILLCELL_X32 FILLER_277_1744 ();
 FILLCELL_X32 FILLER_277_1776 ();
 FILLCELL_X32 FILLER_277_1808 ();
 FILLCELL_X32 FILLER_277_1840 ();
 FILLCELL_X32 FILLER_277_1872 ();
 FILLCELL_X32 FILLER_277_1904 ();
 FILLCELL_X32 FILLER_277_1936 ();
 FILLCELL_X32 FILLER_277_1968 ();
 FILLCELL_X32 FILLER_277_2000 ();
 FILLCELL_X32 FILLER_277_2032 ();
 FILLCELL_X32 FILLER_277_2064 ();
 FILLCELL_X32 FILLER_277_2096 ();
 FILLCELL_X32 FILLER_277_2128 ();
 FILLCELL_X32 FILLER_277_2160 ();
 FILLCELL_X32 FILLER_277_2192 ();
 FILLCELL_X32 FILLER_277_2224 ();
 FILLCELL_X32 FILLER_277_2256 ();
 FILLCELL_X32 FILLER_277_2288 ();
 FILLCELL_X32 FILLER_277_2320 ();
 FILLCELL_X32 FILLER_277_2352 ();
 FILLCELL_X32 FILLER_277_2384 ();
 FILLCELL_X16 FILLER_277_2416 ();
 FILLCELL_X4 FILLER_277_2432 ();
 FILLCELL_X32 FILLER_278_1 ();
 FILLCELL_X32 FILLER_278_33 ();
 FILLCELL_X32 FILLER_278_65 ();
 FILLCELL_X32 FILLER_278_97 ();
 FILLCELL_X32 FILLER_278_129 ();
 FILLCELL_X32 FILLER_278_161 ();
 FILLCELL_X32 FILLER_278_193 ();
 FILLCELL_X32 FILLER_278_225 ();
 FILLCELL_X32 FILLER_278_257 ();
 FILLCELL_X32 FILLER_278_289 ();
 FILLCELL_X32 FILLER_278_321 ();
 FILLCELL_X32 FILLER_278_353 ();
 FILLCELL_X32 FILLER_278_385 ();
 FILLCELL_X32 FILLER_278_417 ();
 FILLCELL_X32 FILLER_278_449 ();
 FILLCELL_X32 FILLER_278_481 ();
 FILLCELL_X32 FILLER_278_513 ();
 FILLCELL_X32 FILLER_278_545 ();
 FILLCELL_X32 FILLER_278_577 ();
 FILLCELL_X16 FILLER_278_609 ();
 FILLCELL_X4 FILLER_278_625 ();
 FILLCELL_X2 FILLER_278_629 ();
 FILLCELL_X32 FILLER_278_632 ();
 FILLCELL_X32 FILLER_278_664 ();
 FILLCELL_X32 FILLER_278_696 ();
 FILLCELL_X32 FILLER_278_728 ();
 FILLCELL_X32 FILLER_278_760 ();
 FILLCELL_X32 FILLER_278_792 ();
 FILLCELL_X32 FILLER_278_824 ();
 FILLCELL_X32 FILLER_278_856 ();
 FILLCELL_X32 FILLER_278_888 ();
 FILLCELL_X32 FILLER_278_920 ();
 FILLCELL_X32 FILLER_278_952 ();
 FILLCELL_X32 FILLER_278_984 ();
 FILLCELL_X32 FILLER_278_1016 ();
 FILLCELL_X32 FILLER_278_1048 ();
 FILLCELL_X32 FILLER_278_1080 ();
 FILLCELL_X32 FILLER_278_1112 ();
 FILLCELL_X32 FILLER_278_1144 ();
 FILLCELL_X32 FILLER_278_1176 ();
 FILLCELL_X32 FILLER_278_1208 ();
 FILLCELL_X32 FILLER_278_1240 ();
 FILLCELL_X32 FILLER_278_1272 ();
 FILLCELL_X32 FILLER_278_1304 ();
 FILLCELL_X32 FILLER_278_1336 ();
 FILLCELL_X32 FILLER_278_1368 ();
 FILLCELL_X32 FILLER_278_1400 ();
 FILLCELL_X32 FILLER_278_1432 ();
 FILLCELL_X32 FILLER_278_1464 ();
 FILLCELL_X32 FILLER_278_1496 ();
 FILLCELL_X32 FILLER_278_1528 ();
 FILLCELL_X32 FILLER_278_1560 ();
 FILLCELL_X32 FILLER_278_1592 ();
 FILLCELL_X32 FILLER_278_1624 ();
 FILLCELL_X32 FILLER_278_1656 ();
 FILLCELL_X32 FILLER_278_1688 ();
 FILLCELL_X32 FILLER_278_1720 ();
 FILLCELL_X32 FILLER_278_1752 ();
 FILLCELL_X32 FILLER_278_1784 ();
 FILLCELL_X32 FILLER_278_1816 ();
 FILLCELL_X32 FILLER_278_1848 ();
 FILLCELL_X8 FILLER_278_1880 ();
 FILLCELL_X4 FILLER_278_1888 ();
 FILLCELL_X2 FILLER_278_1892 ();
 FILLCELL_X32 FILLER_278_1895 ();
 FILLCELL_X32 FILLER_278_1927 ();
 FILLCELL_X32 FILLER_278_1959 ();
 FILLCELL_X32 FILLER_278_1991 ();
 FILLCELL_X32 FILLER_278_2023 ();
 FILLCELL_X32 FILLER_278_2055 ();
 FILLCELL_X32 FILLER_278_2087 ();
 FILLCELL_X32 FILLER_278_2119 ();
 FILLCELL_X32 FILLER_278_2151 ();
 FILLCELL_X32 FILLER_278_2183 ();
 FILLCELL_X32 FILLER_278_2215 ();
 FILLCELL_X32 FILLER_278_2247 ();
 FILLCELL_X32 FILLER_278_2279 ();
 FILLCELL_X32 FILLER_278_2311 ();
 FILLCELL_X32 FILLER_278_2343 ();
 FILLCELL_X32 FILLER_278_2375 ();
 FILLCELL_X16 FILLER_278_2407 ();
 FILLCELL_X8 FILLER_278_2423 ();
 FILLCELL_X4 FILLER_278_2431 ();
 FILLCELL_X1 FILLER_278_2435 ();
 FILLCELL_X32 FILLER_279_1 ();
 FILLCELL_X32 FILLER_279_33 ();
 FILLCELL_X32 FILLER_279_65 ();
 FILLCELL_X32 FILLER_279_97 ();
 FILLCELL_X32 FILLER_279_129 ();
 FILLCELL_X32 FILLER_279_161 ();
 FILLCELL_X32 FILLER_279_193 ();
 FILLCELL_X32 FILLER_279_225 ();
 FILLCELL_X32 FILLER_279_257 ();
 FILLCELL_X32 FILLER_279_289 ();
 FILLCELL_X32 FILLER_279_321 ();
 FILLCELL_X32 FILLER_279_353 ();
 FILLCELL_X32 FILLER_279_385 ();
 FILLCELL_X32 FILLER_279_417 ();
 FILLCELL_X32 FILLER_279_449 ();
 FILLCELL_X32 FILLER_279_481 ();
 FILLCELL_X32 FILLER_279_513 ();
 FILLCELL_X32 FILLER_279_545 ();
 FILLCELL_X32 FILLER_279_577 ();
 FILLCELL_X32 FILLER_279_609 ();
 FILLCELL_X32 FILLER_279_641 ();
 FILLCELL_X32 FILLER_279_673 ();
 FILLCELL_X32 FILLER_279_705 ();
 FILLCELL_X32 FILLER_279_737 ();
 FILLCELL_X32 FILLER_279_769 ();
 FILLCELL_X32 FILLER_279_801 ();
 FILLCELL_X32 FILLER_279_833 ();
 FILLCELL_X32 FILLER_279_865 ();
 FILLCELL_X32 FILLER_279_897 ();
 FILLCELL_X32 FILLER_279_929 ();
 FILLCELL_X32 FILLER_279_961 ();
 FILLCELL_X32 FILLER_279_993 ();
 FILLCELL_X32 FILLER_279_1025 ();
 FILLCELL_X32 FILLER_279_1057 ();
 FILLCELL_X32 FILLER_279_1089 ();
 FILLCELL_X32 FILLER_279_1121 ();
 FILLCELL_X32 FILLER_279_1153 ();
 FILLCELL_X32 FILLER_279_1185 ();
 FILLCELL_X32 FILLER_279_1217 ();
 FILLCELL_X8 FILLER_279_1249 ();
 FILLCELL_X4 FILLER_279_1257 ();
 FILLCELL_X2 FILLER_279_1261 ();
 FILLCELL_X32 FILLER_279_1264 ();
 FILLCELL_X32 FILLER_279_1296 ();
 FILLCELL_X32 FILLER_279_1328 ();
 FILLCELL_X32 FILLER_279_1360 ();
 FILLCELL_X32 FILLER_279_1392 ();
 FILLCELL_X32 FILLER_279_1424 ();
 FILLCELL_X32 FILLER_279_1456 ();
 FILLCELL_X32 FILLER_279_1488 ();
 FILLCELL_X32 FILLER_279_1520 ();
 FILLCELL_X32 FILLER_279_1552 ();
 FILLCELL_X32 FILLER_279_1584 ();
 FILLCELL_X32 FILLER_279_1616 ();
 FILLCELL_X32 FILLER_279_1648 ();
 FILLCELL_X32 FILLER_279_1680 ();
 FILLCELL_X32 FILLER_279_1712 ();
 FILLCELL_X32 FILLER_279_1744 ();
 FILLCELL_X32 FILLER_279_1776 ();
 FILLCELL_X32 FILLER_279_1808 ();
 FILLCELL_X32 FILLER_279_1840 ();
 FILLCELL_X32 FILLER_279_1872 ();
 FILLCELL_X32 FILLER_279_1904 ();
 FILLCELL_X32 FILLER_279_1936 ();
 FILLCELL_X32 FILLER_279_1968 ();
 FILLCELL_X32 FILLER_279_2000 ();
 FILLCELL_X32 FILLER_279_2032 ();
 FILLCELL_X32 FILLER_279_2064 ();
 FILLCELL_X32 FILLER_279_2096 ();
 FILLCELL_X32 FILLER_279_2128 ();
 FILLCELL_X32 FILLER_279_2160 ();
 FILLCELL_X32 FILLER_279_2192 ();
 FILLCELL_X32 FILLER_279_2224 ();
 FILLCELL_X32 FILLER_279_2256 ();
 FILLCELL_X32 FILLER_279_2288 ();
 FILLCELL_X32 FILLER_279_2320 ();
 FILLCELL_X32 FILLER_279_2352 ();
 FILLCELL_X32 FILLER_279_2384 ();
 FILLCELL_X16 FILLER_279_2416 ();
 FILLCELL_X4 FILLER_279_2432 ();
 FILLCELL_X32 FILLER_280_1 ();
 FILLCELL_X32 FILLER_280_33 ();
 FILLCELL_X32 FILLER_280_65 ();
 FILLCELL_X32 FILLER_280_97 ();
 FILLCELL_X32 FILLER_280_129 ();
 FILLCELL_X32 FILLER_280_161 ();
 FILLCELL_X32 FILLER_280_193 ();
 FILLCELL_X32 FILLER_280_225 ();
 FILLCELL_X32 FILLER_280_257 ();
 FILLCELL_X32 FILLER_280_289 ();
 FILLCELL_X32 FILLER_280_321 ();
 FILLCELL_X32 FILLER_280_353 ();
 FILLCELL_X32 FILLER_280_385 ();
 FILLCELL_X32 FILLER_280_417 ();
 FILLCELL_X32 FILLER_280_449 ();
 FILLCELL_X32 FILLER_280_481 ();
 FILLCELL_X32 FILLER_280_513 ();
 FILLCELL_X32 FILLER_280_545 ();
 FILLCELL_X32 FILLER_280_577 ();
 FILLCELL_X16 FILLER_280_609 ();
 FILLCELL_X4 FILLER_280_625 ();
 FILLCELL_X2 FILLER_280_629 ();
 FILLCELL_X32 FILLER_280_632 ();
 FILLCELL_X32 FILLER_280_664 ();
 FILLCELL_X32 FILLER_280_696 ();
 FILLCELL_X32 FILLER_280_728 ();
 FILLCELL_X32 FILLER_280_760 ();
 FILLCELL_X32 FILLER_280_792 ();
 FILLCELL_X32 FILLER_280_824 ();
 FILLCELL_X32 FILLER_280_856 ();
 FILLCELL_X32 FILLER_280_888 ();
 FILLCELL_X32 FILLER_280_920 ();
 FILLCELL_X32 FILLER_280_952 ();
 FILLCELL_X32 FILLER_280_984 ();
 FILLCELL_X32 FILLER_280_1016 ();
 FILLCELL_X32 FILLER_280_1048 ();
 FILLCELL_X32 FILLER_280_1080 ();
 FILLCELL_X32 FILLER_280_1112 ();
 FILLCELL_X32 FILLER_280_1144 ();
 FILLCELL_X32 FILLER_280_1176 ();
 FILLCELL_X32 FILLER_280_1208 ();
 FILLCELL_X32 FILLER_280_1240 ();
 FILLCELL_X32 FILLER_280_1272 ();
 FILLCELL_X32 FILLER_280_1304 ();
 FILLCELL_X32 FILLER_280_1336 ();
 FILLCELL_X32 FILLER_280_1368 ();
 FILLCELL_X32 FILLER_280_1400 ();
 FILLCELL_X32 FILLER_280_1432 ();
 FILLCELL_X32 FILLER_280_1464 ();
 FILLCELL_X32 FILLER_280_1496 ();
 FILLCELL_X32 FILLER_280_1528 ();
 FILLCELL_X32 FILLER_280_1560 ();
 FILLCELL_X32 FILLER_280_1592 ();
 FILLCELL_X32 FILLER_280_1624 ();
 FILLCELL_X32 FILLER_280_1656 ();
 FILLCELL_X32 FILLER_280_1688 ();
 FILLCELL_X32 FILLER_280_1720 ();
 FILLCELL_X32 FILLER_280_1752 ();
 FILLCELL_X32 FILLER_280_1784 ();
 FILLCELL_X32 FILLER_280_1816 ();
 FILLCELL_X32 FILLER_280_1848 ();
 FILLCELL_X8 FILLER_280_1880 ();
 FILLCELL_X4 FILLER_280_1888 ();
 FILLCELL_X2 FILLER_280_1892 ();
 FILLCELL_X32 FILLER_280_1895 ();
 FILLCELL_X32 FILLER_280_1927 ();
 FILLCELL_X32 FILLER_280_1959 ();
 FILLCELL_X32 FILLER_280_1991 ();
 FILLCELL_X32 FILLER_280_2023 ();
 FILLCELL_X32 FILLER_280_2055 ();
 FILLCELL_X32 FILLER_280_2087 ();
 FILLCELL_X32 FILLER_280_2119 ();
 FILLCELL_X32 FILLER_280_2151 ();
 FILLCELL_X32 FILLER_280_2183 ();
 FILLCELL_X32 FILLER_280_2215 ();
 FILLCELL_X32 FILLER_280_2247 ();
 FILLCELL_X32 FILLER_280_2279 ();
 FILLCELL_X32 FILLER_280_2311 ();
 FILLCELL_X32 FILLER_280_2343 ();
 FILLCELL_X32 FILLER_280_2375 ();
 FILLCELL_X16 FILLER_280_2407 ();
 FILLCELL_X8 FILLER_280_2423 ();
 FILLCELL_X4 FILLER_280_2431 ();
 FILLCELL_X1 FILLER_280_2435 ();
 FILLCELL_X32 FILLER_281_1 ();
 FILLCELL_X32 FILLER_281_33 ();
 FILLCELL_X32 FILLER_281_65 ();
 FILLCELL_X32 FILLER_281_97 ();
 FILLCELL_X32 FILLER_281_129 ();
 FILLCELL_X32 FILLER_281_161 ();
 FILLCELL_X32 FILLER_281_193 ();
 FILLCELL_X32 FILLER_281_225 ();
 FILLCELL_X32 FILLER_281_257 ();
 FILLCELL_X32 FILLER_281_289 ();
 FILLCELL_X32 FILLER_281_321 ();
 FILLCELL_X32 FILLER_281_353 ();
 FILLCELL_X32 FILLER_281_385 ();
 FILLCELL_X32 FILLER_281_417 ();
 FILLCELL_X32 FILLER_281_449 ();
 FILLCELL_X32 FILLER_281_481 ();
 FILLCELL_X32 FILLER_281_513 ();
 FILLCELL_X32 FILLER_281_545 ();
 FILLCELL_X32 FILLER_281_577 ();
 FILLCELL_X32 FILLER_281_609 ();
 FILLCELL_X32 FILLER_281_641 ();
 FILLCELL_X32 FILLER_281_673 ();
 FILLCELL_X32 FILLER_281_705 ();
 FILLCELL_X32 FILLER_281_737 ();
 FILLCELL_X32 FILLER_281_769 ();
 FILLCELL_X32 FILLER_281_801 ();
 FILLCELL_X32 FILLER_281_833 ();
 FILLCELL_X32 FILLER_281_865 ();
 FILLCELL_X32 FILLER_281_897 ();
 FILLCELL_X32 FILLER_281_929 ();
 FILLCELL_X32 FILLER_281_961 ();
 FILLCELL_X32 FILLER_281_993 ();
 FILLCELL_X32 FILLER_281_1025 ();
 FILLCELL_X32 FILLER_281_1057 ();
 FILLCELL_X32 FILLER_281_1089 ();
 FILLCELL_X32 FILLER_281_1121 ();
 FILLCELL_X32 FILLER_281_1153 ();
 FILLCELL_X32 FILLER_281_1185 ();
 FILLCELL_X32 FILLER_281_1217 ();
 FILLCELL_X8 FILLER_281_1249 ();
 FILLCELL_X4 FILLER_281_1257 ();
 FILLCELL_X2 FILLER_281_1261 ();
 FILLCELL_X32 FILLER_281_1264 ();
 FILLCELL_X32 FILLER_281_1296 ();
 FILLCELL_X32 FILLER_281_1328 ();
 FILLCELL_X32 FILLER_281_1360 ();
 FILLCELL_X32 FILLER_281_1392 ();
 FILLCELL_X32 FILLER_281_1424 ();
 FILLCELL_X32 FILLER_281_1456 ();
 FILLCELL_X32 FILLER_281_1488 ();
 FILLCELL_X32 FILLER_281_1520 ();
 FILLCELL_X32 FILLER_281_1552 ();
 FILLCELL_X32 FILLER_281_1584 ();
 FILLCELL_X32 FILLER_281_1616 ();
 FILLCELL_X32 FILLER_281_1648 ();
 FILLCELL_X32 FILLER_281_1680 ();
 FILLCELL_X32 FILLER_281_1712 ();
 FILLCELL_X32 FILLER_281_1744 ();
 FILLCELL_X32 FILLER_281_1776 ();
 FILLCELL_X32 FILLER_281_1808 ();
 FILLCELL_X32 FILLER_281_1840 ();
 FILLCELL_X32 FILLER_281_1872 ();
 FILLCELL_X32 FILLER_281_1904 ();
 FILLCELL_X32 FILLER_281_1936 ();
 FILLCELL_X32 FILLER_281_1968 ();
 FILLCELL_X32 FILLER_281_2000 ();
 FILLCELL_X32 FILLER_281_2032 ();
 FILLCELL_X32 FILLER_281_2064 ();
 FILLCELL_X32 FILLER_281_2096 ();
 FILLCELL_X32 FILLER_281_2128 ();
 FILLCELL_X32 FILLER_281_2160 ();
 FILLCELL_X32 FILLER_281_2192 ();
 FILLCELL_X32 FILLER_281_2224 ();
 FILLCELL_X32 FILLER_281_2256 ();
 FILLCELL_X32 FILLER_281_2288 ();
 FILLCELL_X32 FILLER_281_2320 ();
 FILLCELL_X32 FILLER_281_2352 ();
 FILLCELL_X32 FILLER_281_2384 ();
 FILLCELL_X16 FILLER_281_2416 ();
 FILLCELL_X4 FILLER_281_2432 ();
 FILLCELL_X32 FILLER_282_1 ();
 FILLCELL_X32 FILLER_282_33 ();
 FILLCELL_X32 FILLER_282_65 ();
 FILLCELL_X32 FILLER_282_97 ();
 FILLCELL_X32 FILLER_282_129 ();
 FILLCELL_X32 FILLER_282_161 ();
 FILLCELL_X32 FILLER_282_193 ();
 FILLCELL_X32 FILLER_282_225 ();
 FILLCELL_X32 FILLER_282_257 ();
 FILLCELL_X32 FILLER_282_289 ();
 FILLCELL_X32 FILLER_282_321 ();
 FILLCELL_X32 FILLER_282_353 ();
 FILLCELL_X32 FILLER_282_385 ();
 FILLCELL_X32 FILLER_282_417 ();
 FILLCELL_X32 FILLER_282_449 ();
 FILLCELL_X32 FILLER_282_481 ();
 FILLCELL_X32 FILLER_282_513 ();
 FILLCELL_X32 FILLER_282_545 ();
 FILLCELL_X32 FILLER_282_577 ();
 FILLCELL_X16 FILLER_282_609 ();
 FILLCELL_X4 FILLER_282_625 ();
 FILLCELL_X2 FILLER_282_629 ();
 FILLCELL_X32 FILLER_282_632 ();
 FILLCELL_X32 FILLER_282_664 ();
 FILLCELL_X32 FILLER_282_696 ();
 FILLCELL_X32 FILLER_282_728 ();
 FILLCELL_X32 FILLER_282_760 ();
 FILLCELL_X32 FILLER_282_792 ();
 FILLCELL_X32 FILLER_282_824 ();
 FILLCELL_X32 FILLER_282_856 ();
 FILLCELL_X32 FILLER_282_888 ();
 FILLCELL_X32 FILLER_282_920 ();
 FILLCELL_X32 FILLER_282_952 ();
 FILLCELL_X32 FILLER_282_984 ();
 FILLCELL_X32 FILLER_282_1016 ();
 FILLCELL_X32 FILLER_282_1048 ();
 FILLCELL_X32 FILLER_282_1080 ();
 FILLCELL_X32 FILLER_282_1112 ();
 FILLCELL_X32 FILLER_282_1144 ();
 FILLCELL_X32 FILLER_282_1176 ();
 FILLCELL_X32 FILLER_282_1208 ();
 FILLCELL_X32 FILLER_282_1240 ();
 FILLCELL_X32 FILLER_282_1272 ();
 FILLCELL_X32 FILLER_282_1304 ();
 FILLCELL_X32 FILLER_282_1336 ();
 FILLCELL_X32 FILLER_282_1368 ();
 FILLCELL_X32 FILLER_282_1400 ();
 FILLCELL_X32 FILLER_282_1432 ();
 FILLCELL_X32 FILLER_282_1464 ();
 FILLCELL_X32 FILLER_282_1496 ();
 FILLCELL_X32 FILLER_282_1528 ();
 FILLCELL_X32 FILLER_282_1560 ();
 FILLCELL_X32 FILLER_282_1592 ();
 FILLCELL_X32 FILLER_282_1624 ();
 FILLCELL_X32 FILLER_282_1656 ();
 FILLCELL_X32 FILLER_282_1688 ();
 FILLCELL_X32 FILLER_282_1720 ();
 FILLCELL_X32 FILLER_282_1752 ();
 FILLCELL_X32 FILLER_282_1784 ();
 FILLCELL_X32 FILLER_282_1816 ();
 FILLCELL_X32 FILLER_282_1848 ();
 FILLCELL_X8 FILLER_282_1880 ();
 FILLCELL_X4 FILLER_282_1888 ();
 FILLCELL_X2 FILLER_282_1892 ();
 FILLCELL_X32 FILLER_282_1895 ();
 FILLCELL_X32 FILLER_282_1927 ();
 FILLCELL_X32 FILLER_282_1959 ();
 FILLCELL_X32 FILLER_282_1991 ();
 FILLCELL_X32 FILLER_282_2023 ();
 FILLCELL_X32 FILLER_282_2055 ();
 FILLCELL_X32 FILLER_282_2087 ();
 FILLCELL_X32 FILLER_282_2119 ();
 FILLCELL_X32 FILLER_282_2151 ();
 FILLCELL_X32 FILLER_282_2183 ();
 FILLCELL_X32 FILLER_282_2215 ();
 FILLCELL_X32 FILLER_282_2247 ();
 FILLCELL_X32 FILLER_282_2279 ();
 FILLCELL_X32 FILLER_282_2311 ();
 FILLCELL_X32 FILLER_282_2343 ();
 FILLCELL_X32 FILLER_282_2375 ();
 FILLCELL_X16 FILLER_282_2407 ();
 FILLCELL_X8 FILLER_282_2423 ();
 FILLCELL_X4 FILLER_282_2431 ();
 FILLCELL_X1 FILLER_282_2435 ();
 FILLCELL_X32 FILLER_283_1 ();
 FILLCELL_X32 FILLER_283_33 ();
 FILLCELL_X32 FILLER_283_65 ();
 FILLCELL_X32 FILLER_283_97 ();
 FILLCELL_X32 FILLER_283_129 ();
 FILLCELL_X32 FILLER_283_161 ();
 FILLCELL_X32 FILLER_283_193 ();
 FILLCELL_X32 FILLER_283_225 ();
 FILLCELL_X32 FILLER_283_257 ();
 FILLCELL_X32 FILLER_283_289 ();
 FILLCELL_X32 FILLER_283_321 ();
 FILLCELL_X32 FILLER_283_353 ();
 FILLCELL_X32 FILLER_283_385 ();
 FILLCELL_X32 FILLER_283_417 ();
 FILLCELL_X32 FILLER_283_449 ();
 FILLCELL_X32 FILLER_283_481 ();
 FILLCELL_X32 FILLER_283_513 ();
 FILLCELL_X32 FILLER_283_545 ();
 FILLCELL_X32 FILLER_283_577 ();
 FILLCELL_X32 FILLER_283_609 ();
 FILLCELL_X32 FILLER_283_641 ();
 FILLCELL_X32 FILLER_283_673 ();
 FILLCELL_X32 FILLER_283_705 ();
 FILLCELL_X32 FILLER_283_737 ();
 FILLCELL_X32 FILLER_283_769 ();
 FILLCELL_X32 FILLER_283_801 ();
 FILLCELL_X32 FILLER_283_833 ();
 FILLCELL_X32 FILLER_283_865 ();
 FILLCELL_X32 FILLER_283_897 ();
 FILLCELL_X32 FILLER_283_929 ();
 FILLCELL_X32 FILLER_283_961 ();
 FILLCELL_X32 FILLER_283_993 ();
 FILLCELL_X32 FILLER_283_1025 ();
 FILLCELL_X32 FILLER_283_1057 ();
 FILLCELL_X32 FILLER_283_1089 ();
 FILLCELL_X32 FILLER_283_1121 ();
 FILLCELL_X32 FILLER_283_1153 ();
 FILLCELL_X32 FILLER_283_1185 ();
 FILLCELL_X32 FILLER_283_1217 ();
 FILLCELL_X8 FILLER_283_1249 ();
 FILLCELL_X4 FILLER_283_1257 ();
 FILLCELL_X2 FILLER_283_1261 ();
 FILLCELL_X32 FILLER_283_1264 ();
 FILLCELL_X32 FILLER_283_1296 ();
 FILLCELL_X32 FILLER_283_1328 ();
 FILLCELL_X32 FILLER_283_1360 ();
 FILLCELL_X32 FILLER_283_1392 ();
 FILLCELL_X32 FILLER_283_1424 ();
 FILLCELL_X32 FILLER_283_1456 ();
 FILLCELL_X32 FILLER_283_1488 ();
 FILLCELL_X32 FILLER_283_1520 ();
 FILLCELL_X32 FILLER_283_1552 ();
 FILLCELL_X32 FILLER_283_1584 ();
 FILLCELL_X32 FILLER_283_1616 ();
 FILLCELL_X32 FILLER_283_1648 ();
 FILLCELL_X32 FILLER_283_1680 ();
 FILLCELL_X32 FILLER_283_1712 ();
 FILLCELL_X32 FILLER_283_1744 ();
 FILLCELL_X32 FILLER_283_1776 ();
 FILLCELL_X32 FILLER_283_1808 ();
 FILLCELL_X32 FILLER_283_1840 ();
 FILLCELL_X32 FILLER_283_1872 ();
 FILLCELL_X32 FILLER_283_1904 ();
 FILLCELL_X32 FILLER_283_1936 ();
 FILLCELL_X32 FILLER_283_1968 ();
 FILLCELL_X32 FILLER_283_2000 ();
 FILLCELL_X32 FILLER_283_2032 ();
 FILLCELL_X32 FILLER_283_2064 ();
 FILLCELL_X32 FILLER_283_2096 ();
 FILLCELL_X32 FILLER_283_2128 ();
 FILLCELL_X32 FILLER_283_2160 ();
 FILLCELL_X32 FILLER_283_2192 ();
 FILLCELL_X32 FILLER_283_2224 ();
 FILLCELL_X32 FILLER_283_2256 ();
 FILLCELL_X32 FILLER_283_2288 ();
 FILLCELL_X32 FILLER_283_2320 ();
 FILLCELL_X32 FILLER_283_2352 ();
 FILLCELL_X32 FILLER_283_2384 ();
 FILLCELL_X16 FILLER_283_2416 ();
 FILLCELL_X4 FILLER_283_2432 ();
 FILLCELL_X32 FILLER_284_1 ();
 FILLCELL_X32 FILLER_284_33 ();
 FILLCELL_X32 FILLER_284_65 ();
 FILLCELL_X32 FILLER_284_97 ();
 FILLCELL_X32 FILLER_284_129 ();
 FILLCELL_X32 FILLER_284_161 ();
 FILLCELL_X32 FILLER_284_193 ();
 FILLCELL_X32 FILLER_284_225 ();
 FILLCELL_X32 FILLER_284_257 ();
 FILLCELL_X32 FILLER_284_289 ();
 FILLCELL_X32 FILLER_284_321 ();
 FILLCELL_X32 FILLER_284_353 ();
 FILLCELL_X32 FILLER_284_385 ();
 FILLCELL_X32 FILLER_284_417 ();
 FILLCELL_X32 FILLER_284_449 ();
 FILLCELL_X32 FILLER_284_481 ();
 FILLCELL_X32 FILLER_284_513 ();
 FILLCELL_X32 FILLER_284_545 ();
 FILLCELL_X32 FILLER_284_577 ();
 FILLCELL_X16 FILLER_284_609 ();
 FILLCELL_X4 FILLER_284_625 ();
 FILLCELL_X2 FILLER_284_629 ();
 FILLCELL_X32 FILLER_284_632 ();
 FILLCELL_X32 FILLER_284_664 ();
 FILLCELL_X32 FILLER_284_696 ();
 FILLCELL_X32 FILLER_284_728 ();
 FILLCELL_X32 FILLER_284_760 ();
 FILLCELL_X32 FILLER_284_792 ();
 FILLCELL_X32 FILLER_284_824 ();
 FILLCELL_X32 FILLER_284_856 ();
 FILLCELL_X32 FILLER_284_888 ();
 FILLCELL_X32 FILLER_284_920 ();
 FILLCELL_X32 FILLER_284_952 ();
 FILLCELL_X32 FILLER_284_984 ();
 FILLCELL_X32 FILLER_284_1016 ();
 FILLCELL_X32 FILLER_284_1048 ();
 FILLCELL_X32 FILLER_284_1080 ();
 FILLCELL_X32 FILLER_284_1112 ();
 FILLCELL_X32 FILLER_284_1144 ();
 FILLCELL_X32 FILLER_284_1176 ();
 FILLCELL_X32 FILLER_284_1208 ();
 FILLCELL_X32 FILLER_284_1240 ();
 FILLCELL_X32 FILLER_284_1272 ();
 FILLCELL_X32 FILLER_284_1304 ();
 FILLCELL_X32 FILLER_284_1336 ();
 FILLCELL_X32 FILLER_284_1368 ();
 FILLCELL_X32 FILLER_284_1400 ();
 FILLCELL_X32 FILLER_284_1432 ();
 FILLCELL_X32 FILLER_284_1464 ();
 FILLCELL_X32 FILLER_284_1496 ();
 FILLCELL_X32 FILLER_284_1528 ();
 FILLCELL_X32 FILLER_284_1560 ();
 FILLCELL_X32 FILLER_284_1592 ();
 FILLCELL_X32 FILLER_284_1624 ();
 FILLCELL_X32 FILLER_284_1656 ();
 FILLCELL_X32 FILLER_284_1688 ();
 FILLCELL_X32 FILLER_284_1720 ();
 FILLCELL_X32 FILLER_284_1752 ();
 FILLCELL_X32 FILLER_284_1784 ();
 FILLCELL_X32 FILLER_284_1816 ();
 FILLCELL_X32 FILLER_284_1848 ();
 FILLCELL_X8 FILLER_284_1880 ();
 FILLCELL_X4 FILLER_284_1888 ();
 FILLCELL_X2 FILLER_284_1892 ();
 FILLCELL_X32 FILLER_284_1895 ();
 FILLCELL_X32 FILLER_284_1927 ();
 FILLCELL_X32 FILLER_284_1959 ();
 FILLCELL_X32 FILLER_284_1991 ();
 FILLCELL_X32 FILLER_284_2023 ();
 FILLCELL_X32 FILLER_284_2055 ();
 FILLCELL_X32 FILLER_284_2087 ();
 FILLCELL_X32 FILLER_284_2119 ();
 FILLCELL_X32 FILLER_284_2151 ();
 FILLCELL_X32 FILLER_284_2183 ();
 FILLCELL_X32 FILLER_284_2215 ();
 FILLCELL_X32 FILLER_284_2247 ();
 FILLCELL_X32 FILLER_284_2279 ();
 FILLCELL_X32 FILLER_284_2311 ();
 FILLCELL_X32 FILLER_284_2343 ();
 FILLCELL_X32 FILLER_284_2375 ();
 FILLCELL_X16 FILLER_284_2407 ();
 FILLCELL_X8 FILLER_284_2423 ();
 FILLCELL_X4 FILLER_284_2431 ();
 FILLCELL_X1 FILLER_284_2435 ();
 FILLCELL_X32 FILLER_285_1 ();
 FILLCELL_X32 FILLER_285_33 ();
 FILLCELL_X32 FILLER_285_65 ();
 FILLCELL_X32 FILLER_285_97 ();
 FILLCELL_X32 FILLER_285_129 ();
 FILLCELL_X32 FILLER_285_161 ();
 FILLCELL_X32 FILLER_285_193 ();
 FILLCELL_X32 FILLER_285_225 ();
 FILLCELL_X32 FILLER_285_257 ();
 FILLCELL_X32 FILLER_285_289 ();
 FILLCELL_X32 FILLER_285_321 ();
 FILLCELL_X32 FILLER_285_353 ();
 FILLCELL_X32 FILLER_285_385 ();
 FILLCELL_X32 FILLER_285_417 ();
 FILLCELL_X32 FILLER_285_449 ();
 FILLCELL_X32 FILLER_285_481 ();
 FILLCELL_X32 FILLER_285_513 ();
 FILLCELL_X32 FILLER_285_545 ();
 FILLCELL_X32 FILLER_285_577 ();
 FILLCELL_X32 FILLER_285_609 ();
 FILLCELL_X32 FILLER_285_641 ();
 FILLCELL_X32 FILLER_285_673 ();
 FILLCELL_X32 FILLER_285_705 ();
 FILLCELL_X32 FILLER_285_737 ();
 FILLCELL_X32 FILLER_285_769 ();
 FILLCELL_X32 FILLER_285_801 ();
 FILLCELL_X32 FILLER_285_833 ();
 FILLCELL_X32 FILLER_285_865 ();
 FILLCELL_X32 FILLER_285_897 ();
 FILLCELL_X32 FILLER_285_929 ();
 FILLCELL_X32 FILLER_285_961 ();
 FILLCELL_X32 FILLER_285_993 ();
 FILLCELL_X32 FILLER_285_1025 ();
 FILLCELL_X32 FILLER_285_1057 ();
 FILLCELL_X16 FILLER_285_1089 ();
 FILLCELL_X8 FILLER_285_1105 ();
 FILLCELL_X4 FILLER_285_1113 ();
 FILLCELL_X1 FILLER_285_1117 ();
 FILLCELL_X32 FILLER_285_1121 ();
 FILLCELL_X32 FILLER_285_1153 ();
 FILLCELL_X32 FILLER_285_1185 ();
 FILLCELL_X32 FILLER_285_1217 ();
 FILLCELL_X8 FILLER_285_1249 ();
 FILLCELL_X4 FILLER_285_1257 ();
 FILLCELL_X2 FILLER_285_1261 ();
 FILLCELL_X32 FILLER_285_1264 ();
 FILLCELL_X32 FILLER_285_1296 ();
 FILLCELL_X32 FILLER_285_1328 ();
 FILLCELL_X32 FILLER_285_1360 ();
 FILLCELL_X32 FILLER_285_1392 ();
 FILLCELL_X32 FILLER_285_1424 ();
 FILLCELL_X32 FILLER_285_1456 ();
 FILLCELL_X32 FILLER_285_1488 ();
 FILLCELL_X32 FILLER_285_1520 ();
 FILLCELL_X32 FILLER_285_1552 ();
 FILLCELL_X32 FILLER_285_1584 ();
 FILLCELL_X32 FILLER_285_1616 ();
 FILLCELL_X32 FILLER_285_1648 ();
 FILLCELL_X32 FILLER_285_1680 ();
 FILLCELL_X32 FILLER_285_1712 ();
 FILLCELL_X32 FILLER_285_1744 ();
 FILLCELL_X32 FILLER_285_1776 ();
 FILLCELL_X32 FILLER_285_1808 ();
 FILLCELL_X32 FILLER_285_1840 ();
 FILLCELL_X32 FILLER_285_1872 ();
 FILLCELL_X32 FILLER_285_1904 ();
 FILLCELL_X32 FILLER_285_1936 ();
 FILLCELL_X32 FILLER_285_1968 ();
 FILLCELL_X32 FILLER_285_2000 ();
 FILLCELL_X32 FILLER_285_2032 ();
 FILLCELL_X32 FILLER_285_2064 ();
 FILLCELL_X32 FILLER_285_2096 ();
 FILLCELL_X32 FILLER_285_2128 ();
 FILLCELL_X32 FILLER_285_2160 ();
 FILLCELL_X32 FILLER_285_2192 ();
 FILLCELL_X32 FILLER_285_2224 ();
 FILLCELL_X32 FILLER_285_2256 ();
 FILLCELL_X32 FILLER_285_2288 ();
 FILLCELL_X32 FILLER_285_2320 ();
 FILLCELL_X32 FILLER_285_2352 ();
 FILLCELL_X32 FILLER_285_2384 ();
 FILLCELL_X16 FILLER_285_2416 ();
 FILLCELL_X4 FILLER_285_2432 ();
 FILLCELL_X32 FILLER_286_1 ();
 FILLCELL_X32 FILLER_286_33 ();
 FILLCELL_X32 FILLER_286_65 ();
 FILLCELL_X32 FILLER_286_97 ();
 FILLCELL_X32 FILLER_286_129 ();
 FILLCELL_X32 FILLER_286_161 ();
 FILLCELL_X32 FILLER_286_193 ();
 FILLCELL_X32 FILLER_286_225 ();
 FILLCELL_X32 FILLER_286_257 ();
 FILLCELL_X32 FILLER_286_289 ();
 FILLCELL_X32 FILLER_286_321 ();
 FILLCELL_X32 FILLER_286_353 ();
 FILLCELL_X32 FILLER_286_385 ();
 FILLCELL_X32 FILLER_286_417 ();
 FILLCELL_X32 FILLER_286_449 ();
 FILLCELL_X32 FILLER_286_481 ();
 FILLCELL_X32 FILLER_286_513 ();
 FILLCELL_X32 FILLER_286_545 ();
 FILLCELL_X32 FILLER_286_577 ();
 FILLCELL_X16 FILLER_286_609 ();
 FILLCELL_X4 FILLER_286_625 ();
 FILLCELL_X2 FILLER_286_629 ();
 FILLCELL_X32 FILLER_286_632 ();
 FILLCELL_X32 FILLER_286_664 ();
 FILLCELL_X32 FILLER_286_696 ();
 FILLCELL_X32 FILLER_286_728 ();
 FILLCELL_X32 FILLER_286_760 ();
 FILLCELL_X32 FILLER_286_792 ();
 FILLCELL_X32 FILLER_286_824 ();
 FILLCELL_X32 FILLER_286_856 ();
 FILLCELL_X32 FILLER_286_888 ();
 FILLCELL_X32 FILLER_286_920 ();
 FILLCELL_X32 FILLER_286_952 ();
 FILLCELL_X32 FILLER_286_984 ();
 FILLCELL_X32 FILLER_286_1016 ();
 FILLCELL_X32 FILLER_286_1048 ();
 FILLCELL_X2 FILLER_286_1080 ();
 FILLCELL_X1 FILLER_286_1082 ();
 FILLCELL_X4 FILLER_286_1086 ();
 FILLCELL_X1 FILLER_286_1090 ();
 FILLCELL_X2 FILLER_286_1105 ();
 FILLCELL_X2 FILLER_286_1110 ();
 FILLCELL_X1 FILLER_286_1112 ();
 FILLCELL_X1 FILLER_286_1131 ();
 FILLCELL_X16 FILLER_286_1135 ();
 FILLCELL_X4 FILLER_286_1151 ();
 FILLCELL_X2 FILLER_286_1155 ();
 FILLCELL_X1 FILLER_286_1157 ();
 FILLCELL_X32 FILLER_286_1165 ();
 FILLCELL_X32 FILLER_286_1197 ();
 FILLCELL_X32 FILLER_286_1229 ();
 FILLCELL_X32 FILLER_286_1261 ();
 FILLCELL_X32 FILLER_286_1293 ();
 FILLCELL_X32 FILLER_286_1325 ();
 FILLCELL_X32 FILLER_286_1357 ();
 FILLCELL_X32 FILLER_286_1389 ();
 FILLCELL_X32 FILLER_286_1421 ();
 FILLCELL_X32 FILLER_286_1453 ();
 FILLCELL_X32 FILLER_286_1485 ();
 FILLCELL_X32 FILLER_286_1517 ();
 FILLCELL_X32 FILLER_286_1549 ();
 FILLCELL_X32 FILLER_286_1581 ();
 FILLCELL_X32 FILLER_286_1613 ();
 FILLCELL_X32 FILLER_286_1645 ();
 FILLCELL_X32 FILLER_286_1677 ();
 FILLCELL_X32 FILLER_286_1709 ();
 FILLCELL_X32 FILLER_286_1741 ();
 FILLCELL_X32 FILLER_286_1773 ();
 FILLCELL_X32 FILLER_286_1805 ();
 FILLCELL_X32 FILLER_286_1837 ();
 FILLCELL_X16 FILLER_286_1869 ();
 FILLCELL_X8 FILLER_286_1885 ();
 FILLCELL_X1 FILLER_286_1893 ();
 FILLCELL_X32 FILLER_286_1895 ();
 FILLCELL_X32 FILLER_286_1927 ();
 FILLCELL_X32 FILLER_286_1959 ();
 FILLCELL_X32 FILLER_286_1991 ();
 FILLCELL_X32 FILLER_286_2023 ();
 FILLCELL_X32 FILLER_286_2055 ();
 FILLCELL_X32 FILLER_286_2087 ();
 FILLCELL_X32 FILLER_286_2119 ();
 FILLCELL_X32 FILLER_286_2151 ();
 FILLCELL_X32 FILLER_286_2183 ();
 FILLCELL_X32 FILLER_286_2215 ();
 FILLCELL_X32 FILLER_286_2247 ();
 FILLCELL_X32 FILLER_286_2279 ();
 FILLCELL_X32 FILLER_286_2311 ();
 FILLCELL_X32 FILLER_286_2343 ();
 FILLCELL_X32 FILLER_286_2375 ();
 FILLCELL_X16 FILLER_286_2407 ();
 FILLCELL_X8 FILLER_286_2423 ();
 FILLCELL_X4 FILLER_286_2431 ();
 FILLCELL_X1 FILLER_286_2435 ();
 FILLCELL_X32 FILLER_287_1 ();
 FILLCELL_X32 FILLER_287_33 ();
 FILLCELL_X32 FILLER_287_65 ();
 FILLCELL_X32 FILLER_287_97 ();
 FILLCELL_X32 FILLER_287_129 ();
 FILLCELL_X32 FILLER_287_161 ();
 FILLCELL_X32 FILLER_287_193 ();
 FILLCELL_X32 FILLER_287_225 ();
 FILLCELL_X32 FILLER_287_257 ();
 FILLCELL_X32 FILLER_287_289 ();
 FILLCELL_X32 FILLER_287_321 ();
 FILLCELL_X32 FILLER_287_353 ();
 FILLCELL_X32 FILLER_287_385 ();
 FILLCELL_X32 FILLER_287_417 ();
 FILLCELL_X32 FILLER_287_449 ();
 FILLCELL_X32 FILLER_287_481 ();
 FILLCELL_X32 FILLER_287_513 ();
 FILLCELL_X32 FILLER_287_545 ();
 FILLCELL_X32 FILLER_287_577 ();
 FILLCELL_X32 FILLER_287_609 ();
 FILLCELL_X32 FILLER_287_641 ();
 FILLCELL_X32 FILLER_287_673 ();
 FILLCELL_X32 FILLER_287_705 ();
 FILLCELL_X32 FILLER_287_737 ();
 FILLCELL_X32 FILLER_287_769 ();
 FILLCELL_X32 FILLER_287_801 ();
 FILLCELL_X32 FILLER_287_833 ();
 FILLCELL_X32 FILLER_287_865 ();
 FILLCELL_X32 FILLER_287_897 ();
 FILLCELL_X32 FILLER_287_929 ();
 FILLCELL_X32 FILLER_287_961 ();
 FILLCELL_X32 FILLER_287_993 ();
 FILLCELL_X32 FILLER_287_1025 ();
 FILLCELL_X16 FILLER_287_1057 ();
 FILLCELL_X4 FILLER_287_1140 ();
 FILLCELL_X1 FILLER_287_1156 ();
 FILLCELL_X16 FILLER_287_1171 ();
 FILLCELL_X8 FILLER_287_1187 ();
 FILLCELL_X4 FILLER_287_1195 ();
 FILLCELL_X1 FILLER_287_1199 ();
 FILLCELL_X32 FILLER_287_1209 ();
 FILLCELL_X16 FILLER_287_1241 ();
 FILLCELL_X4 FILLER_287_1257 ();
 FILLCELL_X2 FILLER_287_1261 ();
 FILLCELL_X32 FILLER_287_1264 ();
 FILLCELL_X32 FILLER_287_1296 ();
 FILLCELL_X32 FILLER_287_1328 ();
 FILLCELL_X32 FILLER_287_1360 ();
 FILLCELL_X32 FILLER_287_1392 ();
 FILLCELL_X32 FILLER_287_1424 ();
 FILLCELL_X32 FILLER_287_1456 ();
 FILLCELL_X32 FILLER_287_1488 ();
 FILLCELL_X32 FILLER_287_1520 ();
 FILLCELL_X32 FILLER_287_1552 ();
 FILLCELL_X32 FILLER_287_1584 ();
 FILLCELL_X32 FILLER_287_1616 ();
 FILLCELL_X32 FILLER_287_1648 ();
 FILLCELL_X32 FILLER_287_1680 ();
 FILLCELL_X32 FILLER_287_1712 ();
 FILLCELL_X32 FILLER_287_1744 ();
 FILLCELL_X32 FILLER_287_1776 ();
 FILLCELL_X32 FILLER_287_1808 ();
 FILLCELL_X32 FILLER_287_1840 ();
 FILLCELL_X32 FILLER_287_1872 ();
 FILLCELL_X32 FILLER_287_1904 ();
 FILLCELL_X32 FILLER_287_1936 ();
 FILLCELL_X32 FILLER_287_1968 ();
 FILLCELL_X32 FILLER_287_2000 ();
 FILLCELL_X32 FILLER_287_2032 ();
 FILLCELL_X32 FILLER_287_2064 ();
 FILLCELL_X32 FILLER_287_2096 ();
 FILLCELL_X32 FILLER_287_2128 ();
 FILLCELL_X32 FILLER_287_2160 ();
 FILLCELL_X32 FILLER_287_2192 ();
 FILLCELL_X32 FILLER_287_2224 ();
 FILLCELL_X32 FILLER_287_2256 ();
 FILLCELL_X32 FILLER_287_2288 ();
 FILLCELL_X32 FILLER_287_2320 ();
 FILLCELL_X32 FILLER_287_2352 ();
 FILLCELL_X32 FILLER_287_2384 ();
 FILLCELL_X16 FILLER_287_2416 ();
 FILLCELL_X4 FILLER_287_2432 ();
 FILLCELL_X32 FILLER_288_1 ();
 FILLCELL_X32 FILLER_288_33 ();
 FILLCELL_X32 FILLER_288_65 ();
 FILLCELL_X32 FILLER_288_97 ();
 FILLCELL_X32 FILLER_288_129 ();
 FILLCELL_X32 FILLER_288_161 ();
 FILLCELL_X32 FILLER_288_193 ();
 FILLCELL_X32 FILLER_288_225 ();
 FILLCELL_X32 FILLER_288_257 ();
 FILLCELL_X32 FILLER_288_289 ();
 FILLCELL_X32 FILLER_288_321 ();
 FILLCELL_X32 FILLER_288_353 ();
 FILLCELL_X32 FILLER_288_385 ();
 FILLCELL_X32 FILLER_288_417 ();
 FILLCELL_X32 FILLER_288_449 ();
 FILLCELL_X32 FILLER_288_481 ();
 FILLCELL_X32 FILLER_288_513 ();
 FILLCELL_X32 FILLER_288_545 ();
 FILLCELL_X32 FILLER_288_577 ();
 FILLCELL_X16 FILLER_288_609 ();
 FILLCELL_X4 FILLER_288_625 ();
 FILLCELL_X2 FILLER_288_629 ();
 FILLCELL_X32 FILLER_288_632 ();
 FILLCELL_X32 FILLER_288_664 ();
 FILLCELL_X32 FILLER_288_696 ();
 FILLCELL_X32 FILLER_288_728 ();
 FILLCELL_X32 FILLER_288_760 ();
 FILLCELL_X32 FILLER_288_792 ();
 FILLCELL_X32 FILLER_288_824 ();
 FILLCELL_X32 FILLER_288_856 ();
 FILLCELL_X32 FILLER_288_888 ();
 FILLCELL_X32 FILLER_288_920 ();
 FILLCELL_X32 FILLER_288_952 ();
 FILLCELL_X32 FILLER_288_984 ();
 FILLCELL_X32 FILLER_288_1016 ();
 FILLCELL_X8 FILLER_288_1048 ();
 FILLCELL_X4 FILLER_288_1056 ();
 FILLCELL_X4 FILLER_288_1064 ();
 FILLCELL_X1 FILLER_288_1068 ();
 FILLCELL_X2 FILLER_288_1108 ();
 FILLCELL_X8 FILLER_288_1147 ();
 FILLCELL_X8 FILLER_288_1168 ();
 FILLCELL_X4 FILLER_288_1176 ();
 FILLCELL_X1 FILLER_288_1180 ();
 FILLCELL_X32 FILLER_288_1217 ();
 FILLCELL_X32 FILLER_288_1249 ();
 FILLCELL_X32 FILLER_288_1281 ();
 FILLCELL_X32 FILLER_288_1313 ();
 FILLCELL_X32 FILLER_288_1345 ();
 FILLCELL_X32 FILLER_288_1377 ();
 FILLCELL_X32 FILLER_288_1409 ();
 FILLCELL_X32 FILLER_288_1441 ();
 FILLCELL_X32 FILLER_288_1473 ();
 FILLCELL_X32 FILLER_288_1505 ();
 FILLCELL_X32 FILLER_288_1537 ();
 FILLCELL_X32 FILLER_288_1569 ();
 FILLCELL_X32 FILLER_288_1601 ();
 FILLCELL_X32 FILLER_288_1633 ();
 FILLCELL_X32 FILLER_288_1665 ();
 FILLCELL_X32 FILLER_288_1697 ();
 FILLCELL_X32 FILLER_288_1729 ();
 FILLCELL_X32 FILLER_288_1761 ();
 FILLCELL_X32 FILLER_288_1793 ();
 FILLCELL_X32 FILLER_288_1825 ();
 FILLCELL_X32 FILLER_288_1857 ();
 FILLCELL_X4 FILLER_288_1889 ();
 FILLCELL_X1 FILLER_288_1893 ();
 FILLCELL_X32 FILLER_288_1895 ();
 FILLCELL_X32 FILLER_288_1927 ();
 FILLCELL_X32 FILLER_288_1959 ();
 FILLCELL_X32 FILLER_288_1991 ();
 FILLCELL_X32 FILLER_288_2023 ();
 FILLCELL_X32 FILLER_288_2055 ();
 FILLCELL_X32 FILLER_288_2087 ();
 FILLCELL_X32 FILLER_288_2119 ();
 FILLCELL_X32 FILLER_288_2151 ();
 FILLCELL_X32 FILLER_288_2183 ();
 FILLCELL_X32 FILLER_288_2215 ();
 FILLCELL_X32 FILLER_288_2247 ();
 FILLCELL_X32 FILLER_288_2279 ();
 FILLCELL_X32 FILLER_288_2311 ();
 FILLCELL_X32 FILLER_288_2343 ();
 FILLCELL_X32 FILLER_288_2375 ();
 FILLCELL_X16 FILLER_288_2407 ();
 FILLCELL_X8 FILLER_288_2423 ();
 FILLCELL_X4 FILLER_288_2431 ();
 FILLCELL_X1 FILLER_288_2435 ();
 FILLCELL_X32 FILLER_289_1 ();
 FILLCELL_X32 FILLER_289_33 ();
 FILLCELL_X32 FILLER_289_65 ();
 FILLCELL_X32 FILLER_289_97 ();
 FILLCELL_X32 FILLER_289_129 ();
 FILLCELL_X32 FILLER_289_161 ();
 FILLCELL_X32 FILLER_289_193 ();
 FILLCELL_X32 FILLER_289_225 ();
 FILLCELL_X32 FILLER_289_257 ();
 FILLCELL_X32 FILLER_289_289 ();
 FILLCELL_X32 FILLER_289_321 ();
 FILLCELL_X32 FILLER_289_353 ();
 FILLCELL_X32 FILLER_289_385 ();
 FILLCELL_X32 FILLER_289_417 ();
 FILLCELL_X32 FILLER_289_449 ();
 FILLCELL_X32 FILLER_289_481 ();
 FILLCELL_X32 FILLER_289_513 ();
 FILLCELL_X32 FILLER_289_545 ();
 FILLCELL_X32 FILLER_289_577 ();
 FILLCELL_X32 FILLER_289_609 ();
 FILLCELL_X32 FILLER_289_641 ();
 FILLCELL_X32 FILLER_289_673 ();
 FILLCELL_X32 FILLER_289_705 ();
 FILLCELL_X32 FILLER_289_737 ();
 FILLCELL_X32 FILLER_289_769 ();
 FILLCELL_X32 FILLER_289_801 ();
 FILLCELL_X32 FILLER_289_833 ();
 FILLCELL_X32 FILLER_289_865 ();
 FILLCELL_X32 FILLER_289_897 ();
 FILLCELL_X32 FILLER_289_929 ();
 FILLCELL_X32 FILLER_289_961 ();
 FILLCELL_X32 FILLER_289_993 ();
 FILLCELL_X32 FILLER_289_1025 ();
 FILLCELL_X4 FILLER_289_1057 ();
 FILLCELL_X2 FILLER_289_1061 ();
 FILLCELL_X1 FILLER_289_1082 ();
 FILLCELL_X16 FILLER_289_1107 ();
 FILLCELL_X16 FILLER_289_1131 ();
 FILLCELL_X4 FILLER_289_1147 ();
 FILLCELL_X2 FILLER_289_1151 ();
 FILLCELL_X2 FILLER_289_1167 ();
 FILLCELL_X2 FILLER_289_1182 ();
 FILLCELL_X32 FILLER_289_1220 ();
 FILLCELL_X8 FILLER_289_1252 ();
 FILLCELL_X2 FILLER_289_1260 ();
 FILLCELL_X1 FILLER_289_1262 ();
 FILLCELL_X32 FILLER_289_1264 ();
 FILLCELL_X32 FILLER_289_1296 ();
 FILLCELL_X32 FILLER_289_1328 ();
 FILLCELL_X32 FILLER_289_1360 ();
 FILLCELL_X32 FILLER_289_1392 ();
 FILLCELL_X32 FILLER_289_1424 ();
 FILLCELL_X32 FILLER_289_1456 ();
 FILLCELL_X32 FILLER_289_1488 ();
 FILLCELL_X32 FILLER_289_1520 ();
 FILLCELL_X32 FILLER_289_1552 ();
 FILLCELL_X32 FILLER_289_1584 ();
 FILLCELL_X32 FILLER_289_1616 ();
 FILLCELL_X32 FILLER_289_1648 ();
 FILLCELL_X32 FILLER_289_1680 ();
 FILLCELL_X32 FILLER_289_1712 ();
 FILLCELL_X32 FILLER_289_1744 ();
 FILLCELL_X32 FILLER_289_1776 ();
 FILLCELL_X32 FILLER_289_1808 ();
 FILLCELL_X32 FILLER_289_1840 ();
 FILLCELL_X32 FILLER_289_1872 ();
 FILLCELL_X32 FILLER_289_1904 ();
 FILLCELL_X32 FILLER_289_1936 ();
 FILLCELL_X32 FILLER_289_1968 ();
 FILLCELL_X32 FILLER_289_2000 ();
 FILLCELL_X32 FILLER_289_2032 ();
 FILLCELL_X32 FILLER_289_2064 ();
 FILLCELL_X32 FILLER_289_2096 ();
 FILLCELL_X32 FILLER_289_2128 ();
 FILLCELL_X32 FILLER_289_2160 ();
 FILLCELL_X32 FILLER_289_2192 ();
 FILLCELL_X32 FILLER_289_2224 ();
 FILLCELL_X32 FILLER_289_2256 ();
 FILLCELL_X32 FILLER_289_2288 ();
 FILLCELL_X32 FILLER_289_2320 ();
 FILLCELL_X32 FILLER_289_2352 ();
 FILLCELL_X32 FILLER_289_2384 ();
 FILLCELL_X16 FILLER_289_2416 ();
 FILLCELL_X4 FILLER_289_2432 ();
 FILLCELL_X32 FILLER_290_1 ();
 FILLCELL_X32 FILLER_290_33 ();
 FILLCELL_X32 FILLER_290_65 ();
 FILLCELL_X32 FILLER_290_97 ();
 FILLCELL_X32 FILLER_290_129 ();
 FILLCELL_X32 FILLER_290_161 ();
 FILLCELL_X32 FILLER_290_193 ();
 FILLCELL_X32 FILLER_290_225 ();
 FILLCELL_X32 FILLER_290_257 ();
 FILLCELL_X32 FILLER_290_289 ();
 FILLCELL_X32 FILLER_290_321 ();
 FILLCELL_X32 FILLER_290_353 ();
 FILLCELL_X32 FILLER_290_385 ();
 FILLCELL_X32 FILLER_290_417 ();
 FILLCELL_X32 FILLER_290_449 ();
 FILLCELL_X32 FILLER_290_481 ();
 FILLCELL_X32 FILLER_290_513 ();
 FILLCELL_X32 FILLER_290_545 ();
 FILLCELL_X32 FILLER_290_577 ();
 FILLCELL_X16 FILLER_290_609 ();
 FILLCELL_X4 FILLER_290_625 ();
 FILLCELL_X2 FILLER_290_629 ();
 FILLCELL_X32 FILLER_290_632 ();
 FILLCELL_X32 FILLER_290_664 ();
 FILLCELL_X32 FILLER_290_696 ();
 FILLCELL_X32 FILLER_290_728 ();
 FILLCELL_X32 FILLER_290_760 ();
 FILLCELL_X32 FILLER_290_792 ();
 FILLCELL_X32 FILLER_290_824 ();
 FILLCELL_X32 FILLER_290_856 ();
 FILLCELL_X32 FILLER_290_888 ();
 FILLCELL_X32 FILLER_290_920 ();
 FILLCELL_X32 FILLER_290_952 ();
 FILLCELL_X32 FILLER_290_984 ();
 FILLCELL_X32 FILLER_290_1016 ();
 FILLCELL_X16 FILLER_290_1048 ();
 FILLCELL_X1 FILLER_290_1064 ();
 FILLCELL_X2 FILLER_290_1116 ();
 FILLCELL_X1 FILLER_290_1118 ();
 FILLCELL_X8 FILLER_290_1128 ();
 FILLCELL_X2 FILLER_290_1136 ();
 FILLCELL_X16 FILLER_290_1144 ();
 FILLCELL_X2 FILLER_290_1160 ();
 FILLCELL_X2 FILLER_290_1197 ();
 FILLCELL_X32 FILLER_290_1213 ();
 FILLCELL_X32 FILLER_290_1245 ();
 FILLCELL_X32 FILLER_290_1277 ();
 FILLCELL_X32 FILLER_290_1309 ();
 FILLCELL_X32 FILLER_290_1341 ();
 FILLCELL_X32 FILLER_290_1373 ();
 FILLCELL_X32 FILLER_290_1405 ();
 FILLCELL_X32 FILLER_290_1437 ();
 FILLCELL_X32 FILLER_290_1469 ();
 FILLCELL_X32 FILLER_290_1501 ();
 FILLCELL_X32 FILLER_290_1533 ();
 FILLCELL_X32 FILLER_290_1565 ();
 FILLCELL_X32 FILLER_290_1597 ();
 FILLCELL_X32 FILLER_290_1629 ();
 FILLCELL_X32 FILLER_290_1661 ();
 FILLCELL_X32 FILLER_290_1693 ();
 FILLCELL_X32 FILLER_290_1725 ();
 FILLCELL_X32 FILLER_290_1757 ();
 FILLCELL_X32 FILLER_290_1789 ();
 FILLCELL_X32 FILLER_290_1821 ();
 FILLCELL_X32 FILLER_290_1853 ();
 FILLCELL_X8 FILLER_290_1885 ();
 FILLCELL_X1 FILLER_290_1893 ();
 FILLCELL_X32 FILLER_290_1895 ();
 FILLCELL_X32 FILLER_290_1927 ();
 FILLCELL_X32 FILLER_290_1959 ();
 FILLCELL_X32 FILLER_290_1991 ();
 FILLCELL_X32 FILLER_290_2023 ();
 FILLCELL_X32 FILLER_290_2055 ();
 FILLCELL_X32 FILLER_290_2087 ();
 FILLCELL_X32 FILLER_290_2119 ();
 FILLCELL_X32 FILLER_290_2151 ();
 FILLCELL_X32 FILLER_290_2183 ();
 FILLCELL_X32 FILLER_290_2215 ();
 FILLCELL_X32 FILLER_290_2247 ();
 FILLCELL_X32 FILLER_290_2279 ();
 FILLCELL_X32 FILLER_290_2311 ();
 FILLCELL_X32 FILLER_290_2343 ();
 FILLCELL_X32 FILLER_290_2375 ();
 FILLCELL_X16 FILLER_290_2407 ();
 FILLCELL_X8 FILLER_290_2423 ();
 FILLCELL_X4 FILLER_290_2431 ();
 FILLCELL_X1 FILLER_290_2435 ();
 FILLCELL_X32 FILLER_291_1 ();
 FILLCELL_X32 FILLER_291_33 ();
 FILLCELL_X32 FILLER_291_65 ();
 FILLCELL_X32 FILLER_291_97 ();
 FILLCELL_X32 FILLER_291_129 ();
 FILLCELL_X32 FILLER_291_161 ();
 FILLCELL_X32 FILLER_291_193 ();
 FILLCELL_X32 FILLER_291_225 ();
 FILLCELL_X32 FILLER_291_257 ();
 FILLCELL_X32 FILLER_291_289 ();
 FILLCELL_X32 FILLER_291_321 ();
 FILLCELL_X32 FILLER_291_353 ();
 FILLCELL_X32 FILLER_291_385 ();
 FILLCELL_X32 FILLER_291_417 ();
 FILLCELL_X32 FILLER_291_449 ();
 FILLCELL_X32 FILLER_291_481 ();
 FILLCELL_X32 FILLER_291_513 ();
 FILLCELL_X32 FILLER_291_545 ();
 FILLCELL_X32 FILLER_291_577 ();
 FILLCELL_X32 FILLER_291_609 ();
 FILLCELL_X32 FILLER_291_641 ();
 FILLCELL_X32 FILLER_291_673 ();
 FILLCELL_X32 FILLER_291_705 ();
 FILLCELL_X32 FILLER_291_737 ();
 FILLCELL_X32 FILLER_291_769 ();
 FILLCELL_X32 FILLER_291_801 ();
 FILLCELL_X32 FILLER_291_833 ();
 FILLCELL_X32 FILLER_291_865 ();
 FILLCELL_X32 FILLER_291_897 ();
 FILLCELL_X32 FILLER_291_929 ();
 FILLCELL_X32 FILLER_291_961 ();
 FILLCELL_X32 FILLER_291_993 ();
 FILLCELL_X16 FILLER_291_1025 ();
 FILLCELL_X8 FILLER_291_1041 ();
 FILLCELL_X2 FILLER_291_1049 ();
 FILLCELL_X2 FILLER_291_1092 ();
 FILLCELL_X8 FILLER_291_1104 ();
 FILLCELL_X4 FILLER_291_1112 ();
 FILLCELL_X2 FILLER_291_1116 ();
 FILLCELL_X2 FILLER_291_1131 ();
 FILLCELL_X1 FILLER_291_1133 ();
 FILLCELL_X8 FILLER_291_1144 ();
 FILLCELL_X2 FILLER_291_1152 ();
 FILLCELL_X32 FILLER_291_1171 ();
 FILLCELL_X8 FILLER_291_1203 ();
 FILLCELL_X2 FILLER_291_1211 ();
 FILLCELL_X8 FILLER_291_1222 ();
 FILLCELL_X4 FILLER_291_1230 ();
 FILLCELL_X1 FILLER_291_1234 ();
 FILLCELL_X4 FILLER_291_1240 ();
 FILLCELL_X2 FILLER_291_1244 ();
 FILLCELL_X1 FILLER_291_1246 ();
 FILLCELL_X4 FILLER_291_1259 ();
 FILLCELL_X32 FILLER_291_1264 ();
 FILLCELL_X32 FILLER_291_1296 ();
 FILLCELL_X32 FILLER_291_1328 ();
 FILLCELL_X32 FILLER_291_1360 ();
 FILLCELL_X32 FILLER_291_1392 ();
 FILLCELL_X32 FILLER_291_1424 ();
 FILLCELL_X32 FILLER_291_1456 ();
 FILLCELL_X32 FILLER_291_1488 ();
 FILLCELL_X32 FILLER_291_1520 ();
 FILLCELL_X32 FILLER_291_1552 ();
 FILLCELL_X32 FILLER_291_1584 ();
 FILLCELL_X32 FILLER_291_1616 ();
 FILLCELL_X32 FILLER_291_1648 ();
 FILLCELL_X32 FILLER_291_1680 ();
 FILLCELL_X32 FILLER_291_1712 ();
 FILLCELL_X32 FILLER_291_1744 ();
 FILLCELL_X32 FILLER_291_1776 ();
 FILLCELL_X32 FILLER_291_1808 ();
 FILLCELL_X32 FILLER_291_1840 ();
 FILLCELL_X32 FILLER_291_1872 ();
 FILLCELL_X32 FILLER_291_1904 ();
 FILLCELL_X32 FILLER_291_1936 ();
 FILLCELL_X32 FILLER_291_1968 ();
 FILLCELL_X32 FILLER_291_2000 ();
 FILLCELL_X32 FILLER_291_2032 ();
 FILLCELL_X32 FILLER_291_2064 ();
 FILLCELL_X32 FILLER_291_2096 ();
 FILLCELL_X32 FILLER_291_2128 ();
 FILLCELL_X32 FILLER_291_2160 ();
 FILLCELL_X32 FILLER_291_2192 ();
 FILLCELL_X32 FILLER_291_2224 ();
 FILLCELL_X32 FILLER_291_2256 ();
 FILLCELL_X32 FILLER_291_2288 ();
 FILLCELL_X32 FILLER_291_2320 ();
 FILLCELL_X32 FILLER_291_2352 ();
 FILLCELL_X32 FILLER_291_2384 ();
 FILLCELL_X16 FILLER_291_2416 ();
 FILLCELL_X4 FILLER_291_2432 ();
 FILLCELL_X32 FILLER_292_1 ();
 FILLCELL_X32 FILLER_292_33 ();
 FILLCELL_X32 FILLER_292_65 ();
 FILLCELL_X32 FILLER_292_97 ();
 FILLCELL_X32 FILLER_292_129 ();
 FILLCELL_X32 FILLER_292_161 ();
 FILLCELL_X32 FILLER_292_193 ();
 FILLCELL_X32 FILLER_292_225 ();
 FILLCELL_X32 FILLER_292_257 ();
 FILLCELL_X32 FILLER_292_289 ();
 FILLCELL_X32 FILLER_292_321 ();
 FILLCELL_X32 FILLER_292_353 ();
 FILLCELL_X32 FILLER_292_385 ();
 FILLCELL_X32 FILLER_292_417 ();
 FILLCELL_X32 FILLER_292_449 ();
 FILLCELL_X32 FILLER_292_481 ();
 FILLCELL_X32 FILLER_292_513 ();
 FILLCELL_X32 FILLER_292_545 ();
 FILLCELL_X32 FILLER_292_577 ();
 FILLCELL_X16 FILLER_292_609 ();
 FILLCELL_X4 FILLER_292_625 ();
 FILLCELL_X2 FILLER_292_629 ();
 FILLCELL_X32 FILLER_292_632 ();
 FILLCELL_X32 FILLER_292_664 ();
 FILLCELL_X32 FILLER_292_696 ();
 FILLCELL_X32 FILLER_292_728 ();
 FILLCELL_X32 FILLER_292_760 ();
 FILLCELL_X32 FILLER_292_792 ();
 FILLCELL_X32 FILLER_292_824 ();
 FILLCELL_X32 FILLER_292_856 ();
 FILLCELL_X32 FILLER_292_888 ();
 FILLCELL_X32 FILLER_292_920 ();
 FILLCELL_X32 FILLER_292_952 ();
 FILLCELL_X32 FILLER_292_984 ();
 FILLCELL_X1 FILLER_292_1016 ();
 FILLCELL_X16 FILLER_292_1027 ();
 FILLCELL_X8 FILLER_292_1043 ();
 FILLCELL_X8 FILLER_292_1096 ();
 FILLCELL_X2 FILLER_292_1104 ();
 FILLCELL_X1 FILLER_292_1106 ();
 FILLCELL_X1 FILLER_292_1125 ();
 FILLCELL_X4 FILLER_292_1148 ();
 FILLCELL_X2 FILLER_292_1152 ();
 FILLCELL_X1 FILLER_292_1154 ();
 FILLCELL_X8 FILLER_292_1164 ();
 FILLCELL_X2 FILLER_292_1172 ();
 FILLCELL_X32 FILLER_292_1186 ();
 FILLCELL_X4 FILLER_292_1218 ();
 FILLCELL_X2 FILLER_292_1222 ();
 FILLCELL_X8 FILLER_292_1229 ();
 FILLCELL_X4 FILLER_292_1247 ();
 FILLCELL_X32 FILLER_292_1255 ();
 FILLCELL_X32 FILLER_292_1287 ();
 FILLCELL_X32 FILLER_292_1319 ();
 FILLCELL_X32 FILLER_292_1351 ();
 FILLCELL_X32 FILLER_292_1383 ();
 FILLCELL_X32 FILLER_292_1415 ();
 FILLCELL_X32 FILLER_292_1447 ();
 FILLCELL_X32 FILLER_292_1479 ();
 FILLCELL_X32 FILLER_292_1511 ();
 FILLCELL_X32 FILLER_292_1543 ();
 FILLCELL_X32 FILLER_292_1575 ();
 FILLCELL_X32 FILLER_292_1607 ();
 FILLCELL_X32 FILLER_292_1639 ();
 FILLCELL_X32 FILLER_292_1671 ();
 FILLCELL_X32 FILLER_292_1703 ();
 FILLCELL_X32 FILLER_292_1735 ();
 FILLCELL_X32 FILLER_292_1767 ();
 FILLCELL_X32 FILLER_292_1799 ();
 FILLCELL_X32 FILLER_292_1831 ();
 FILLCELL_X16 FILLER_292_1863 ();
 FILLCELL_X8 FILLER_292_1879 ();
 FILLCELL_X4 FILLER_292_1887 ();
 FILLCELL_X2 FILLER_292_1891 ();
 FILLCELL_X1 FILLER_292_1893 ();
 FILLCELL_X32 FILLER_292_1895 ();
 FILLCELL_X32 FILLER_292_1927 ();
 FILLCELL_X32 FILLER_292_1959 ();
 FILLCELL_X32 FILLER_292_1991 ();
 FILLCELL_X32 FILLER_292_2023 ();
 FILLCELL_X32 FILLER_292_2055 ();
 FILLCELL_X32 FILLER_292_2087 ();
 FILLCELL_X32 FILLER_292_2119 ();
 FILLCELL_X32 FILLER_292_2151 ();
 FILLCELL_X32 FILLER_292_2183 ();
 FILLCELL_X32 FILLER_292_2215 ();
 FILLCELL_X32 FILLER_292_2247 ();
 FILLCELL_X32 FILLER_292_2279 ();
 FILLCELL_X32 FILLER_292_2311 ();
 FILLCELL_X32 FILLER_292_2343 ();
 FILLCELL_X32 FILLER_292_2375 ();
 FILLCELL_X16 FILLER_292_2407 ();
 FILLCELL_X8 FILLER_292_2423 ();
 FILLCELL_X4 FILLER_292_2431 ();
 FILLCELL_X1 FILLER_292_2435 ();
 FILLCELL_X32 FILLER_293_1 ();
 FILLCELL_X32 FILLER_293_33 ();
 FILLCELL_X32 FILLER_293_65 ();
 FILLCELL_X32 FILLER_293_97 ();
 FILLCELL_X32 FILLER_293_129 ();
 FILLCELL_X32 FILLER_293_161 ();
 FILLCELL_X32 FILLER_293_193 ();
 FILLCELL_X32 FILLER_293_225 ();
 FILLCELL_X32 FILLER_293_257 ();
 FILLCELL_X32 FILLER_293_289 ();
 FILLCELL_X32 FILLER_293_321 ();
 FILLCELL_X32 FILLER_293_353 ();
 FILLCELL_X32 FILLER_293_385 ();
 FILLCELL_X32 FILLER_293_417 ();
 FILLCELL_X32 FILLER_293_449 ();
 FILLCELL_X32 FILLER_293_481 ();
 FILLCELL_X32 FILLER_293_513 ();
 FILLCELL_X32 FILLER_293_545 ();
 FILLCELL_X32 FILLER_293_577 ();
 FILLCELL_X32 FILLER_293_609 ();
 FILLCELL_X32 FILLER_293_641 ();
 FILLCELL_X32 FILLER_293_673 ();
 FILLCELL_X32 FILLER_293_705 ();
 FILLCELL_X32 FILLER_293_737 ();
 FILLCELL_X32 FILLER_293_769 ();
 FILLCELL_X32 FILLER_293_801 ();
 FILLCELL_X32 FILLER_293_833 ();
 FILLCELL_X32 FILLER_293_865 ();
 FILLCELL_X32 FILLER_293_897 ();
 FILLCELL_X32 FILLER_293_929 ();
 FILLCELL_X32 FILLER_293_961 ();
 FILLCELL_X8 FILLER_293_993 ();
 FILLCELL_X4 FILLER_293_1001 ();
 FILLCELL_X8 FILLER_293_1007 ();
 FILLCELL_X4 FILLER_293_1015 ();
 FILLCELL_X2 FILLER_293_1019 ();
 FILLCELL_X16 FILLER_293_1031 ();
 FILLCELL_X4 FILLER_293_1047 ();
 FILLCELL_X2 FILLER_293_1051 ();
 FILLCELL_X1 FILLER_293_1053 ();
 FILLCELL_X1 FILLER_293_1064 ();
 FILLCELL_X1 FILLER_293_1088 ();
 FILLCELL_X16 FILLER_293_1094 ();
 FILLCELL_X8 FILLER_293_1110 ();
 FILLCELL_X1 FILLER_293_1118 ();
 FILLCELL_X16 FILLER_293_1155 ();
 FILLCELL_X1 FILLER_293_1171 ();
 FILLCELL_X16 FILLER_293_1176 ();
 FILLCELL_X8 FILLER_293_1192 ();
 FILLCELL_X16 FILLER_293_1207 ();
 FILLCELL_X1 FILLER_293_1223 ();
 FILLCELL_X8 FILLER_293_1264 ();
 FILLCELL_X32 FILLER_293_1282 ();
 FILLCELL_X32 FILLER_293_1314 ();
 FILLCELL_X32 FILLER_293_1346 ();
 FILLCELL_X32 FILLER_293_1378 ();
 FILLCELL_X32 FILLER_293_1410 ();
 FILLCELL_X32 FILLER_293_1442 ();
 FILLCELL_X32 FILLER_293_1474 ();
 FILLCELL_X32 FILLER_293_1506 ();
 FILLCELL_X32 FILLER_293_1538 ();
 FILLCELL_X32 FILLER_293_1570 ();
 FILLCELL_X32 FILLER_293_1602 ();
 FILLCELL_X32 FILLER_293_1634 ();
 FILLCELL_X32 FILLER_293_1666 ();
 FILLCELL_X32 FILLER_293_1698 ();
 FILLCELL_X32 FILLER_293_1730 ();
 FILLCELL_X32 FILLER_293_1762 ();
 FILLCELL_X32 FILLER_293_1794 ();
 FILLCELL_X32 FILLER_293_1826 ();
 FILLCELL_X32 FILLER_293_1858 ();
 FILLCELL_X32 FILLER_293_1890 ();
 FILLCELL_X32 FILLER_293_1922 ();
 FILLCELL_X32 FILLER_293_1954 ();
 FILLCELL_X32 FILLER_293_1986 ();
 FILLCELL_X32 FILLER_293_2018 ();
 FILLCELL_X32 FILLER_293_2050 ();
 FILLCELL_X32 FILLER_293_2082 ();
 FILLCELL_X32 FILLER_293_2114 ();
 FILLCELL_X32 FILLER_293_2146 ();
 FILLCELL_X32 FILLER_293_2178 ();
 FILLCELL_X32 FILLER_293_2210 ();
 FILLCELL_X32 FILLER_293_2242 ();
 FILLCELL_X32 FILLER_293_2274 ();
 FILLCELL_X32 FILLER_293_2306 ();
 FILLCELL_X32 FILLER_293_2338 ();
 FILLCELL_X32 FILLER_293_2370 ();
 FILLCELL_X32 FILLER_293_2402 ();
 FILLCELL_X2 FILLER_293_2434 ();
 FILLCELL_X32 FILLER_294_1 ();
 FILLCELL_X32 FILLER_294_33 ();
 FILLCELL_X32 FILLER_294_65 ();
 FILLCELL_X32 FILLER_294_97 ();
 FILLCELL_X32 FILLER_294_129 ();
 FILLCELL_X32 FILLER_294_161 ();
 FILLCELL_X32 FILLER_294_193 ();
 FILLCELL_X32 FILLER_294_225 ();
 FILLCELL_X32 FILLER_294_257 ();
 FILLCELL_X32 FILLER_294_289 ();
 FILLCELL_X32 FILLER_294_321 ();
 FILLCELL_X32 FILLER_294_353 ();
 FILLCELL_X32 FILLER_294_385 ();
 FILLCELL_X32 FILLER_294_417 ();
 FILLCELL_X32 FILLER_294_449 ();
 FILLCELL_X32 FILLER_294_481 ();
 FILLCELL_X32 FILLER_294_513 ();
 FILLCELL_X32 FILLER_294_545 ();
 FILLCELL_X32 FILLER_294_577 ();
 FILLCELL_X16 FILLER_294_609 ();
 FILLCELL_X4 FILLER_294_625 ();
 FILLCELL_X2 FILLER_294_629 ();
 FILLCELL_X32 FILLER_294_632 ();
 FILLCELL_X32 FILLER_294_664 ();
 FILLCELL_X32 FILLER_294_696 ();
 FILLCELL_X32 FILLER_294_728 ();
 FILLCELL_X32 FILLER_294_760 ();
 FILLCELL_X32 FILLER_294_792 ();
 FILLCELL_X32 FILLER_294_824 ();
 FILLCELL_X32 FILLER_294_856 ();
 FILLCELL_X32 FILLER_294_888 ();
 FILLCELL_X32 FILLER_294_920 ();
 FILLCELL_X32 FILLER_294_952 ();
 FILLCELL_X16 FILLER_294_984 ();
 FILLCELL_X8 FILLER_294_1000 ();
 FILLCELL_X4 FILLER_294_1008 ();
 FILLCELL_X1 FILLER_294_1012 ();
 FILLCELL_X16 FILLER_294_1026 ();
 FILLCELL_X2 FILLER_294_1042 ();
 FILLCELL_X1 FILLER_294_1044 ();
 FILLCELL_X2 FILLER_294_1075 ();
 FILLCELL_X4 FILLER_294_1102 ();
 FILLCELL_X2 FILLER_294_1128 ();
 FILLCELL_X4 FILLER_294_1143 ();
 FILLCELL_X8 FILLER_294_1180 ();
 FILLCELL_X1 FILLER_294_1188 ();
 FILLCELL_X16 FILLER_294_1224 ();
 FILLCELL_X4 FILLER_294_1240 ();
 FILLCELL_X2 FILLER_294_1244 ();
 FILLCELL_X1 FILLER_294_1246 ();
 FILLCELL_X32 FILLER_294_1254 ();
 FILLCELL_X32 FILLER_294_1286 ();
 FILLCELL_X32 FILLER_294_1318 ();
 FILLCELL_X32 FILLER_294_1350 ();
 FILLCELL_X32 FILLER_294_1382 ();
 FILLCELL_X32 FILLER_294_1414 ();
 FILLCELL_X32 FILLER_294_1446 ();
 FILLCELL_X32 FILLER_294_1478 ();
 FILLCELL_X32 FILLER_294_1510 ();
 FILLCELL_X32 FILLER_294_1542 ();
 FILLCELL_X32 FILLER_294_1574 ();
 FILLCELL_X32 FILLER_294_1606 ();
 FILLCELL_X32 FILLER_294_1638 ();
 FILLCELL_X32 FILLER_294_1670 ();
 FILLCELL_X32 FILLER_294_1702 ();
 FILLCELL_X32 FILLER_294_1734 ();
 FILLCELL_X32 FILLER_294_1766 ();
 FILLCELL_X32 FILLER_294_1798 ();
 FILLCELL_X32 FILLER_294_1830 ();
 FILLCELL_X32 FILLER_294_1862 ();
 FILLCELL_X32 FILLER_294_1895 ();
 FILLCELL_X32 FILLER_294_1927 ();
 FILLCELL_X32 FILLER_294_1959 ();
 FILLCELL_X32 FILLER_294_1991 ();
 FILLCELL_X32 FILLER_294_2023 ();
 FILLCELL_X32 FILLER_294_2055 ();
 FILLCELL_X32 FILLER_294_2087 ();
 FILLCELL_X32 FILLER_294_2119 ();
 FILLCELL_X32 FILLER_294_2151 ();
 FILLCELL_X32 FILLER_294_2183 ();
 FILLCELL_X32 FILLER_294_2215 ();
 FILLCELL_X32 FILLER_294_2247 ();
 FILLCELL_X32 FILLER_294_2279 ();
 FILLCELL_X32 FILLER_294_2311 ();
 FILLCELL_X32 FILLER_294_2343 ();
 FILLCELL_X32 FILLER_294_2375 ();
 FILLCELL_X16 FILLER_294_2407 ();
 FILLCELL_X8 FILLER_294_2423 ();
 FILLCELL_X4 FILLER_294_2431 ();
 FILLCELL_X1 FILLER_294_2435 ();
 FILLCELL_X32 FILLER_295_1 ();
 FILLCELL_X32 FILLER_295_33 ();
 FILLCELL_X32 FILLER_295_65 ();
 FILLCELL_X32 FILLER_295_97 ();
 FILLCELL_X32 FILLER_295_129 ();
 FILLCELL_X32 FILLER_295_161 ();
 FILLCELL_X32 FILLER_295_193 ();
 FILLCELL_X32 FILLER_295_225 ();
 FILLCELL_X32 FILLER_295_257 ();
 FILLCELL_X32 FILLER_295_289 ();
 FILLCELL_X32 FILLER_295_321 ();
 FILLCELL_X32 FILLER_295_353 ();
 FILLCELL_X32 FILLER_295_385 ();
 FILLCELL_X32 FILLER_295_417 ();
 FILLCELL_X32 FILLER_295_449 ();
 FILLCELL_X32 FILLER_295_481 ();
 FILLCELL_X32 FILLER_295_513 ();
 FILLCELL_X32 FILLER_295_545 ();
 FILLCELL_X32 FILLER_295_577 ();
 FILLCELL_X32 FILLER_295_609 ();
 FILLCELL_X32 FILLER_295_641 ();
 FILLCELL_X32 FILLER_295_673 ();
 FILLCELL_X32 FILLER_295_705 ();
 FILLCELL_X32 FILLER_295_737 ();
 FILLCELL_X32 FILLER_295_769 ();
 FILLCELL_X32 FILLER_295_801 ();
 FILLCELL_X32 FILLER_295_833 ();
 FILLCELL_X32 FILLER_295_865 ();
 FILLCELL_X32 FILLER_295_897 ();
 FILLCELL_X32 FILLER_295_929 ();
 FILLCELL_X16 FILLER_295_961 ();
 FILLCELL_X8 FILLER_295_977 ();
 FILLCELL_X2 FILLER_295_985 ();
 FILLCELL_X1 FILLER_295_987 ();
 FILLCELL_X8 FILLER_295_993 ();
 FILLCELL_X4 FILLER_295_1001 ();
 FILLCELL_X2 FILLER_295_1005 ();
 FILLCELL_X1 FILLER_295_1007 ();
 FILLCELL_X16 FILLER_295_1026 ();
 FILLCELL_X8 FILLER_295_1042 ();
 FILLCELL_X4 FILLER_295_1050 ();
 FILLCELL_X1 FILLER_295_1054 ();
 FILLCELL_X1 FILLER_295_1059 ();
 FILLCELL_X4 FILLER_295_1097 ();
 FILLCELL_X1 FILLER_295_1101 ();
 FILLCELL_X1 FILLER_295_1111 ();
 FILLCELL_X16 FILLER_295_1133 ();
 FILLCELL_X4 FILLER_295_1149 ();
 FILLCELL_X2 FILLER_295_1153 ();
 FILLCELL_X16 FILLER_295_1164 ();
 FILLCELL_X2 FILLER_295_1180 ();
 FILLCELL_X2 FILLER_295_1188 ();
 FILLCELL_X1 FILLER_295_1207 ();
 FILLCELL_X1 FILLER_295_1217 ();
 FILLCELL_X16 FILLER_295_1233 ();
 FILLCELL_X8 FILLER_295_1249 ();
 FILLCELL_X4 FILLER_295_1257 ();
 FILLCELL_X2 FILLER_295_1261 ();
 FILLCELL_X32 FILLER_295_1264 ();
 FILLCELL_X32 FILLER_295_1296 ();
 FILLCELL_X32 FILLER_295_1328 ();
 FILLCELL_X32 FILLER_295_1360 ();
 FILLCELL_X32 FILLER_295_1392 ();
 FILLCELL_X32 FILLER_295_1424 ();
 FILLCELL_X32 FILLER_295_1456 ();
 FILLCELL_X32 FILLER_295_1488 ();
 FILLCELL_X32 FILLER_295_1520 ();
 FILLCELL_X32 FILLER_295_1552 ();
 FILLCELL_X32 FILLER_295_1584 ();
 FILLCELL_X32 FILLER_295_1616 ();
 FILLCELL_X32 FILLER_295_1648 ();
 FILLCELL_X32 FILLER_295_1680 ();
 FILLCELL_X32 FILLER_295_1712 ();
 FILLCELL_X32 FILLER_295_1744 ();
 FILLCELL_X32 FILLER_295_1776 ();
 FILLCELL_X32 FILLER_295_1808 ();
 FILLCELL_X32 FILLER_295_1840 ();
 FILLCELL_X32 FILLER_295_1872 ();
 FILLCELL_X32 FILLER_295_1904 ();
 FILLCELL_X32 FILLER_295_1936 ();
 FILLCELL_X32 FILLER_295_1968 ();
 FILLCELL_X32 FILLER_295_2000 ();
 FILLCELL_X32 FILLER_295_2032 ();
 FILLCELL_X32 FILLER_295_2064 ();
 FILLCELL_X32 FILLER_295_2096 ();
 FILLCELL_X32 FILLER_295_2128 ();
 FILLCELL_X32 FILLER_295_2160 ();
 FILLCELL_X32 FILLER_295_2192 ();
 FILLCELL_X32 FILLER_295_2224 ();
 FILLCELL_X32 FILLER_295_2256 ();
 FILLCELL_X32 FILLER_295_2288 ();
 FILLCELL_X32 FILLER_295_2320 ();
 FILLCELL_X32 FILLER_295_2352 ();
 FILLCELL_X32 FILLER_295_2384 ();
 FILLCELL_X16 FILLER_295_2416 ();
 FILLCELL_X4 FILLER_295_2432 ();
 FILLCELL_X32 FILLER_296_1 ();
 FILLCELL_X32 FILLER_296_33 ();
 FILLCELL_X32 FILLER_296_65 ();
 FILLCELL_X32 FILLER_296_97 ();
 FILLCELL_X32 FILLER_296_129 ();
 FILLCELL_X32 FILLER_296_161 ();
 FILLCELL_X32 FILLER_296_193 ();
 FILLCELL_X32 FILLER_296_225 ();
 FILLCELL_X32 FILLER_296_257 ();
 FILLCELL_X32 FILLER_296_289 ();
 FILLCELL_X32 FILLER_296_321 ();
 FILLCELL_X32 FILLER_296_353 ();
 FILLCELL_X32 FILLER_296_385 ();
 FILLCELL_X32 FILLER_296_417 ();
 FILLCELL_X32 FILLER_296_449 ();
 FILLCELL_X32 FILLER_296_481 ();
 FILLCELL_X32 FILLER_296_513 ();
 FILLCELL_X32 FILLER_296_545 ();
 FILLCELL_X32 FILLER_296_577 ();
 FILLCELL_X16 FILLER_296_609 ();
 FILLCELL_X4 FILLER_296_625 ();
 FILLCELL_X2 FILLER_296_629 ();
 FILLCELL_X32 FILLER_296_632 ();
 FILLCELL_X32 FILLER_296_664 ();
 FILLCELL_X32 FILLER_296_696 ();
 FILLCELL_X32 FILLER_296_728 ();
 FILLCELL_X32 FILLER_296_760 ();
 FILLCELL_X32 FILLER_296_792 ();
 FILLCELL_X32 FILLER_296_824 ();
 FILLCELL_X32 FILLER_296_856 ();
 FILLCELL_X32 FILLER_296_888 ();
 FILLCELL_X32 FILLER_296_920 ();
 FILLCELL_X32 FILLER_296_952 ();
 FILLCELL_X2 FILLER_296_984 ();
 FILLCELL_X1 FILLER_296_986 ();
 FILLCELL_X8 FILLER_296_1003 ();
 FILLCELL_X4 FILLER_296_1011 ();
 FILLCELL_X1 FILLER_296_1015 ();
 FILLCELL_X8 FILLER_296_1023 ();
 FILLCELL_X4 FILLER_296_1031 ();
 FILLCELL_X1 FILLER_296_1035 ();
 FILLCELL_X16 FILLER_296_1046 ();
 FILLCELL_X2 FILLER_296_1062 ();
 FILLCELL_X1 FILLER_296_1064 ();
 FILLCELL_X8 FILLER_296_1078 ();
 FILLCELL_X8 FILLER_296_1099 ();
 FILLCELL_X2 FILLER_296_1112 ();
 FILLCELL_X16 FILLER_296_1145 ();
 FILLCELL_X8 FILLER_296_1161 ();
 FILLCELL_X4 FILLER_296_1169 ();
 FILLCELL_X1 FILLER_296_1173 ();
 FILLCELL_X4 FILLER_296_1181 ();
 FILLCELL_X4 FILLER_296_1189 ();
 FILLCELL_X2 FILLER_296_1193 ();
 FILLCELL_X4 FILLER_296_1199 ();
 FILLCELL_X1 FILLER_296_1207 ();
 FILLCELL_X8 FILLER_296_1228 ();
 FILLCELL_X2 FILLER_296_1236 ();
 FILLCELL_X2 FILLER_296_1277 ();
 FILLCELL_X32 FILLER_296_1289 ();
 FILLCELL_X32 FILLER_296_1321 ();
 FILLCELL_X32 FILLER_296_1353 ();
 FILLCELL_X32 FILLER_296_1385 ();
 FILLCELL_X32 FILLER_296_1417 ();
 FILLCELL_X32 FILLER_296_1449 ();
 FILLCELL_X32 FILLER_296_1481 ();
 FILLCELL_X32 FILLER_296_1513 ();
 FILLCELL_X32 FILLER_296_1545 ();
 FILLCELL_X32 FILLER_296_1577 ();
 FILLCELL_X32 FILLER_296_1609 ();
 FILLCELL_X32 FILLER_296_1641 ();
 FILLCELL_X32 FILLER_296_1673 ();
 FILLCELL_X32 FILLER_296_1705 ();
 FILLCELL_X32 FILLER_296_1737 ();
 FILLCELL_X32 FILLER_296_1769 ();
 FILLCELL_X32 FILLER_296_1801 ();
 FILLCELL_X32 FILLER_296_1833 ();
 FILLCELL_X16 FILLER_296_1865 ();
 FILLCELL_X8 FILLER_296_1881 ();
 FILLCELL_X4 FILLER_296_1889 ();
 FILLCELL_X1 FILLER_296_1893 ();
 FILLCELL_X32 FILLER_296_1895 ();
 FILLCELL_X32 FILLER_296_1927 ();
 FILLCELL_X32 FILLER_296_1959 ();
 FILLCELL_X32 FILLER_296_1991 ();
 FILLCELL_X32 FILLER_296_2023 ();
 FILLCELL_X32 FILLER_296_2055 ();
 FILLCELL_X32 FILLER_296_2087 ();
 FILLCELL_X32 FILLER_296_2119 ();
 FILLCELL_X32 FILLER_296_2151 ();
 FILLCELL_X32 FILLER_296_2183 ();
 FILLCELL_X32 FILLER_296_2215 ();
 FILLCELL_X32 FILLER_296_2247 ();
 FILLCELL_X32 FILLER_296_2279 ();
 FILLCELL_X32 FILLER_296_2311 ();
 FILLCELL_X32 FILLER_296_2343 ();
 FILLCELL_X32 FILLER_296_2375 ();
 FILLCELL_X16 FILLER_296_2407 ();
 FILLCELL_X8 FILLER_296_2423 ();
 FILLCELL_X4 FILLER_296_2431 ();
 FILLCELL_X1 FILLER_296_2435 ();
 FILLCELL_X32 FILLER_297_1 ();
 FILLCELL_X32 FILLER_297_33 ();
 FILLCELL_X32 FILLER_297_65 ();
 FILLCELL_X32 FILLER_297_97 ();
 FILLCELL_X32 FILLER_297_129 ();
 FILLCELL_X32 FILLER_297_161 ();
 FILLCELL_X32 FILLER_297_193 ();
 FILLCELL_X32 FILLER_297_225 ();
 FILLCELL_X32 FILLER_297_257 ();
 FILLCELL_X32 FILLER_297_289 ();
 FILLCELL_X32 FILLER_297_321 ();
 FILLCELL_X32 FILLER_297_353 ();
 FILLCELL_X32 FILLER_297_385 ();
 FILLCELL_X32 FILLER_297_417 ();
 FILLCELL_X32 FILLER_297_449 ();
 FILLCELL_X32 FILLER_297_481 ();
 FILLCELL_X32 FILLER_297_513 ();
 FILLCELL_X32 FILLER_297_545 ();
 FILLCELL_X32 FILLER_297_577 ();
 FILLCELL_X32 FILLER_297_609 ();
 FILLCELL_X32 FILLER_297_641 ();
 FILLCELL_X32 FILLER_297_673 ();
 FILLCELL_X32 FILLER_297_705 ();
 FILLCELL_X32 FILLER_297_737 ();
 FILLCELL_X32 FILLER_297_769 ();
 FILLCELL_X32 FILLER_297_801 ();
 FILLCELL_X32 FILLER_297_833 ();
 FILLCELL_X32 FILLER_297_865 ();
 FILLCELL_X32 FILLER_297_897 ();
 FILLCELL_X32 FILLER_297_929 ();
 FILLCELL_X16 FILLER_297_961 ();
 FILLCELL_X4 FILLER_297_977 ();
 FILLCELL_X1 FILLER_297_1001 ();
 FILLCELL_X8 FILLER_297_1011 ();
 FILLCELL_X4 FILLER_297_1019 ();
 FILLCELL_X1 FILLER_297_1023 ();
 FILLCELL_X2 FILLER_297_1034 ();
 FILLCELL_X1 FILLER_297_1036 ();
 FILLCELL_X32 FILLER_297_1047 ();
 FILLCELL_X4 FILLER_297_1079 ();
 FILLCELL_X1 FILLER_297_1083 ();
 FILLCELL_X16 FILLER_297_1107 ();
 FILLCELL_X2 FILLER_297_1123 ();
 FILLCELL_X8 FILLER_297_1130 ();
 FILLCELL_X2 FILLER_297_1147 ();
 FILLCELL_X16 FILLER_297_1171 ();
 FILLCELL_X4 FILLER_297_1187 ();
 FILLCELL_X2 FILLER_297_1191 ();
 FILLCELL_X16 FILLER_297_1228 ();
 FILLCELL_X8 FILLER_297_1244 ();
 FILLCELL_X2 FILLER_297_1252 ();
 FILLCELL_X1 FILLER_297_1282 ();
 FILLCELL_X32 FILLER_297_1294 ();
 FILLCELL_X32 FILLER_297_1326 ();
 FILLCELL_X32 FILLER_297_1358 ();
 FILLCELL_X32 FILLER_297_1390 ();
 FILLCELL_X32 FILLER_297_1422 ();
 FILLCELL_X32 FILLER_297_1454 ();
 FILLCELL_X32 FILLER_297_1486 ();
 FILLCELL_X32 FILLER_297_1518 ();
 FILLCELL_X32 FILLER_297_1550 ();
 FILLCELL_X32 FILLER_297_1582 ();
 FILLCELL_X32 FILLER_297_1614 ();
 FILLCELL_X32 FILLER_297_1646 ();
 FILLCELL_X32 FILLER_297_1678 ();
 FILLCELL_X32 FILLER_297_1710 ();
 FILLCELL_X32 FILLER_297_1742 ();
 FILLCELL_X32 FILLER_297_1774 ();
 FILLCELL_X32 FILLER_297_1806 ();
 FILLCELL_X32 FILLER_297_1838 ();
 FILLCELL_X32 FILLER_297_1870 ();
 FILLCELL_X32 FILLER_297_1902 ();
 FILLCELL_X32 FILLER_297_1934 ();
 FILLCELL_X32 FILLER_297_1966 ();
 FILLCELL_X32 FILLER_297_1998 ();
 FILLCELL_X32 FILLER_297_2030 ();
 FILLCELL_X32 FILLER_297_2062 ();
 FILLCELL_X32 FILLER_297_2094 ();
 FILLCELL_X32 FILLER_297_2126 ();
 FILLCELL_X32 FILLER_297_2158 ();
 FILLCELL_X32 FILLER_297_2190 ();
 FILLCELL_X32 FILLER_297_2222 ();
 FILLCELL_X32 FILLER_297_2254 ();
 FILLCELL_X32 FILLER_297_2286 ();
 FILLCELL_X32 FILLER_297_2318 ();
 FILLCELL_X32 FILLER_297_2350 ();
 FILLCELL_X32 FILLER_297_2382 ();
 FILLCELL_X16 FILLER_297_2414 ();
 FILLCELL_X4 FILLER_297_2430 ();
 FILLCELL_X2 FILLER_297_2434 ();
 FILLCELL_X32 FILLER_298_1 ();
 FILLCELL_X32 FILLER_298_33 ();
 FILLCELL_X32 FILLER_298_65 ();
 FILLCELL_X32 FILLER_298_97 ();
 FILLCELL_X32 FILLER_298_129 ();
 FILLCELL_X32 FILLER_298_161 ();
 FILLCELL_X32 FILLER_298_193 ();
 FILLCELL_X32 FILLER_298_225 ();
 FILLCELL_X32 FILLER_298_257 ();
 FILLCELL_X32 FILLER_298_289 ();
 FILLCELL_X32 FILLER_298_321 ();
 FILLCELL_X32 FILLER_298_353 ();
 FILLCELL_X32 FILLER_298_385 ();
 FILLCELL_X32 FILLER_298_417 ();
 FILLCELL_X32 FILLER_298_449 ();
 FILLCELL_X32 FILLER_298_481 ();
 FILLCELL_X32 FILLER_298_513 ();
 FILLCELL_X32 FILLER_298_545 ();
 FILLCELL_X32 FILLER_298_577 ();
 FILLCELL_X16 FILLER_298_609 ();
 FILLCELL_X4 FILLER_298_625 ();
 FILLCELL_X2 FILLER_298_629 ();
 FILLCELL_X32 FILLER_298_632 ();
 FILLCELL_X32 FILLER_298_664 ();
 FILLCELL_X32 FILLER_298_696 ();
 FILLCELL_X32 FILLER_298_728 ();
 FILLCELL_X32 FILLER_298_760 ();
 FILLCELL_X32 FILLER_298_792 ();
 FILLCELL_X32 FILLER_298_824 ();
 FILLCELL_X32 FILLER_298_856 ();
 FILLCELL_X32 FILLER_298_888 ();
 FILLCELL_X32 FILLER_298_920 ();
 FILLCELL_X16 FILLER_298_952 ();
 FILLCELL_X8 FILLER_298_968 ();
 FILLCELL_X4 FILLER_298_976 ();
 FILLCELL_X2 FILLER_298_980 ();
 FILLCELL_X1 FILLER_298_982 ();
 FILLCELL_X2 FILLER_298_986 ();
 FILLCELL_X1 FILLER_298_988 ();
 FILLCELL_X8 FILLER_298_1002 ();
 FILLCELL_X2 FILLER_298_1010 ();
 FILLCELL_X16 FILLER_298_1050 ();
 FILLCELL_X8 FILLER_298_1066 ();
 FILLCELL_X2 FILLER_298_1074 ();
 FILLCELL_X1 FILLER_298_1076 ();
 FILLCELL_X4 FILLER_298_1084 ();
 FILLCELL_X1 FILLER_298_1088 ();
 FILLCELL_X16 FILLER_298_1109 ();
 FILLCELL_X16 FILLER_298_1134 ();
 FILLCELL_X8 FILLER_298_1150 ();
 FILLCELL_X4 FILLER_298_1158 ();
 FILLCELL_X4 FILLER_298_1172 ();
 FILLCELL_X2 FILLER_298_1176 ();
 FILLCELL_X1 FILLER_298_1178 ();
 FILLCELL_X8 FILLER_298_1185 ();
 FILLCELL_X2 FILLER_298_1193 ();
 FILLCELL_X1 FILLER_298_1195 ();
 FILLCELL_X4 FILLER_298_1235 ();
 FILLCELL_X2 FILLER_298_1239 ();
 FILLCELL_X1 FILLER_298_1241 ();
 FILLCELL_X4 FILLER_298_1286 ();
 FILLCELL_X1 FILLER_298_1290 ();
 FILLCELL_X32 FILLER_298_1301 ();
 FILLCELL_X32 FILLER_298_1333 ();
 FILLCELL_X32 FILLER_298_1365 ();
 FILLCELL_X32 FILLER_298_1397 ();
 FILLCELL_X32 FILLER_298_1429 ();
 FILLCELL_X32 FILLER_298_1461 ();
 FILLCELL_X32 FILLER_298_1493 ();
 FILLCELL_X32 FILLER_298_1525 ();
 FILLCELL_X32 FILLER_298_1557 ();
 FILLCELL_X32 FILLER_298_1589 ();
 FILLCELL_X32 FILLER_298_1621 ();
 FILLCELL_X32 FILLER_298_1653 ();
 FILLCELL_X32 FILLER_298_1685 ();
 FILLCELL_X32 FILLER_298_1717 ();
 FILLCELL_X32 FILLER_298_1749 ();
 FILLCELL_X32 FILLER_298_1781 ();
 FILLCELL_X32 FILLER_298_1813 ();
 FILLCELL_X32 FILLER_298_1845 ();
 FILLCELL_X16 FILLER_298_1877 ();
 FILLCELL_X1 FILLER_298_1893 ();
 FILLCELL_X32 FILLER_298_1895 ();
 FILLCELL_X32 FILLER_298_1927 ();
 FILLCELL_X32 FILLER_298_1959 ();
 FILLCELL_X32 FILLER_298_1991 ();
 FILLCELL_X32 FILLER_298_2023 ();
 FILLCELL_X32 FILLER_298_2055 ();
 FILLCELL_X32 FILLER_298_2087 ();
 FILLCELL_X32 FILLER_298_2119 ();
 FILLCELL_X32 FILLER_298_2151 ();
 FILLCELL_X32 FILLER_298_2183 ();
 FILLCELL_X32 FILLER_298_2215 ();
 FILLCELL_X32 FILLER_298_2247 ();
 FILLCELL_X32 FILLER_298_2279 ();
 FILLCELL_X32 FILLER_298_2311 ();
 FILLCELL_X32 FILLER_298_2343 ();
 FILLCELL_X32 FILLER_298_2375 ();
 FILLCELL_X16 FILLER_298_2407 ();
 FILLCELL_X8 FILLER_298_2423 ();
 FILLCELL_X4 FILLER_298_2431 ();
 FILLCELL_X1 FILLER_298_2435 ();
 FILLCELL_X32 FILLER_299_1 ();
 FILLCELL_X32 FILLER_299_33 ();
 FILLCELL_X32 FILLER_299_65 ();
 FILLCELL_X32 FILLER_299_97 ();
 FILLCELL_X32 FILLER_299_129 ();
 FILLCELL_X32 FILLER_299_161 ();
 FILLCELL_X32 FILLER_299_193 ();
 FILLCELL_X32 FILLER_299_225 ();
 FILLCELL_X32 FILLER_299_257 ();
 FILLCELL_X32 FILLER_299_289 ();
 FILLCELL_X32 FILLER_299_321 ();
 FILLCELL_X32 FILLER_299_353 ();
 FILLCELL_X32 FILLER_299_385 ();
 FILLCELL_X32 FILLER_299_417 ();
 FILLCELL_X32 FILLER_299_449 ();
 FILLCELL_X32 FILLER_299_481 ();
 FILLCELL_X32 FILLER_299_513 ();
 FILLCELL_X32 FILLER_299_545 ();
 FILLCELL_X32 FILLER_299_577 ();
 FILLCELL_X32 FILLER_299_609 ();
 FILLCELL_X32 FILLER_299_641 ();
 FILLCELL_X32 FILLER_299_673 ();
 FILLCELL_X32 FILLER_299_705 ();
 FILLCELL_X32 FILLER_299_737 ();
 FILLCELL_X32 FILLER_299_769 ();
 FILLCELL_X32 FILLER_299_801 ();
 FILLCELL_X32 FILLER_299_833 ();
 FILLCELL_X32 FILLER_299_865 ();
 FILLCELL_X32 FILLER_299_897 ();
 FILLCELL_X32 FILLER_299_929 ();
 FILLCELL_X16 FILLER_299_961 ();
 FILLCELL_X8 FILLER_299_977 ();
 FILLCELL_X4 FILLER_299_985 ();
 FILLCELL_X8 FILLER_299_992 ();
 FILLCELL_X4 FILLER_299_1000 ();
 FILLCELL_X1 FILLER_299_1008 ();
 FILLCELL_X2 FILLER_299_1022 ();
 FILLCELL_X4 FILLER_299_1028 ();
 FILLCELL_X2 FILLER_299_1032 ();
 FILLCELL_X1 FILLER_299_1034 ();
 FILLCELL_X8 FILLER_299_1048 ();
 FILLCELL_X4 FILLER_299_1056 ();
 FILLCELL_X2 FILLER_299_1060 ();
 FILLCELL_X8 FILLER_299_1069 ();
 FILLCELL_X8 FILLER_299_1084 ();
 FILLCELL_X1 FILLER_299_1092 ();
 FILLCELL_X16 FILLER_299_1107 ();
 FILLCELL_X4 FILLER_299_1123 ();
 FILLCELL_X2 FILLER_299_1130 ();
 FILLCELL_X1 FILLER_299_1132 ();
 FILLCELL_X8 FILLER_299_1136 ();
 FILLCELL_X1 FILLER_299_1144 ();
 FILLCELL_X4 FILLER_299_1150 ();
 FILLCELL_X2 FILLER_299_1154 ();
 FILLCELL_X1 FILLER_299_1156 ();
 FILLCELL_X1 FILLER_299_1162 ();
 FILLCELL_X2 FILLER_299_1170 ();
 FILLCELL_X2 FILLER_299_1208 ();
 FILLCELL_X1 FILLER_299_1217 ();
 FILLCELL_X32 FILLER_299_1225 ();
 FILLCELL_X4 FILLER_299_1257 ();
 FILLCELL_X2 FILLER_299_1261 ();
 FILLCELL_X16 FILLER_299_1264 ();
 FILLCELL_X8 FILLER_299_1280 ();
 FILLCELL_X2 FILLER_299_1288 ();
 FILLCELL_X1 FILLER_299_1290 ();
 FILLCELL_X4 FILLER_299_1295 ();
 FILLCELL_X32 FILLER_299_1302 ();
 FILLCELL_X32 FILLER_299_1334 ();
 FILLCELL_X32 FILLER_299_1366 ();
 FILLCELL_X32 FILLER_299_1398 ();
 FILLCELL_X32 FILLER_299_1430 ();
 FILLCELL_X32 FILLER_299_1462 ();
 FILLCELL_X32 FILLER_299_1494 ();
 FILLCELL_X32 FILLER_299_1526 ();
 FILLCELL_X32 FILLER_299_1558 ();
 FILLCELL_X32 FILLER_299_1590 ();
 FILLCELL_X32 FILLER_299_1622 ();
 FILLCELL_X32 FILLER_299_1654 ();
 FILLCELL_X32 FILLER_299_1686 ();
 FILLCELL_X32 FILLER_299_1718 ();
 FILLCELL_X32 FILLER_299_1750 ();
 FILLCELL_X32 FILLER_299_1782 ();
 FILLCELL_X32 FILLER_299_1814 ();
 FILLCELL_X32 FILLER_299_1846 ();
 FILLCELL_X32 FILLER_299_1878 ();
 FILLCELL_X32 FILLER_299_1910 ();
 FILLCELL_X32 FILLER_299_1942 ();
 FILLCELL_X32 FILLER_299_1974 ();
 FILLCELL_X32 FILLER_299_2006 ();
 FILLCELL_X32 FILLER_299_2038 ();
 FILLCELL_X32 FILLER_299_2070 ();
 FILLCELL_X32 FILLER_299_2102 ();
 FILLCELL_X32 FILLER_299_2134 ();
 FILLCELL_X32 FILLER_299_2166 ();
 FILLCELL_X32 FILLER_299_2198 ();
 FILLCELL_X32 FILLER_299_2230 ();
 FILLCELL_X32 FILLER_299_2262 ();
 FILLCELL_X32 FILLER_299_2294 ();
 FILLCELL_X32 FILLER_299_2326 ();
 FILLCELL_X32 FILLER_299_2358 ();
 FILLCELL_X32 FILLER_299_2390 ();
 FILLCELL_X8 FILLER_299_2422 ();
 FILLCELL_X4 FILLER_299_2430 ();
 FILLCELL_X2 FILLER_299_2434 ();
 FILLCELL_X32 FILLER_300_1 ();
 FILLCELL_X32 FILLER_300_33 ();
 FILLCELL_X32 FILLER_300_65 ();
 FILLCELL_X32 FILLER_300_97 ();
 FILLCELL_X32 FILLER_300_129 ();
 FILLCELL_X32 FILLER_300_161 ();
 FILLCELL_X32 FILLER_300_193 ();
 FILLCELL_X32 FILLER_300_225 ();
 FILLCELL_X32 FILLER_300_257 ();
 FILLCELL_X32 FILLER_300_289 ();
 FILLCELL_X32 FILLER_300_321 ();
 FILLCELL_X32 FILLER_300_353 ();
 FILLCELL_X32 FILLER_300_385 ();
 FILLCELL_X32 FILLER_300_417 ();
 FILLCELL_X32 FILLER_300_449 ();
 FILLCELL_X32 FILLER_300_481 ();
 FILLCELL_X32 FILLER_300_513 ();
 FILLCELL_X32 FILLER_300_545 ();
 FILLCELL_X32 FILLER_300_577 ();
 FILLCELL_X16 FILLER_300_609 ();
 FILLCELL_X4 FILLER_300_625 ();
 FILLCELL_X2 FILLER_300_629 ();
 FILLCELL_X32 FILLER_300_632 ();
 FILLCELL_X32 FILLER_300_664 ();
 FILLCELL_X32 FILLER_300_696 ();
 FILLCELL_X32 FILLER_300_728 ();
 FILLCELL_X32 FILLER_300_760 ();
 FILLCELL_X32 FILLER_300_792 ();
 FILLCELL_X32 FILLER_300_824 ();
 FILLCELL_X32 FILLER_300_856 ();
 FILLCELL_X32 FILLER_300_888 ();
 FILLCELL_X32 FILLER_300_920 ();
 FILLCELL_X32 FILLER_300_952 ();
 FILLCELL_X16 FILLER_300_984 ();
 FILLCELL_X8 FILLER_300_1000 ();
 FILLCELL_X4 FILLER_300_1008 ();
 FILLCELL_X4 FILLER_300_1025 ();
 FILLCELL_X16 FILLER_300_1035 ();
 FILLCELL_X4 FILLER_300_1051 ();
 FILLCELL_X2 FILLER_300_1055 ();
 FILLCELL_X1 FILLER_300_1057 ();
 FILLCELL_X4 FILLER_300_1063 ();
 FILLCELL_X2 FILLER_300_1067 ();
 FILLCELL_X2 FILLER_300_1075 ();
 FILLCELL_X1 FILLER_300_1077 ();
 FILLCELL_X16 FILLER_300_1085 ();
 FILLCELL_X2 FILLER_300_1101 ();
 FILLCELL_X4 FILLER_300_1110 ();
 FILLCELL_X1 FILLER_300_1114 ();
 FILLCELL_X2 FILLER_300_1141 ();
 FILLCELL_X8 FILLER_300_1148 ();
 FILLCELL_X4 FILLER_300_1156 ();
 FILLCELL_X2 FILLER_300_1160 ();
 FILLCELL_X4 FILLER_300_1181 ();
 FILLCELL_X2 FILLER_300_1185 ();
 FILLCELL_X1 FILLER_300_1187 ();
 FILLCELL_X2 FILLER_300_1226 ();
 FILLCELL_X8 FILLER_300_1235 ();
 FILLCELL_X4 FILLER_300_1243 ();
 FILLCELL_X2 FILLER_300_1247 ();
 FILLCELL_X2 FILLER_300_1253 ();
 FILLCELL_X1 FILLER_300_1255 ();
 FILLCELL_X16 FILLER_300_1260 ();
 FILLCELL_X2 FILLER_300_1276 ();
 FILLCELL_X1 FILLER_300_1281 ();
 FILLCELL_X4 FILLER_300_1286 ();
 FILLCELL_X2 FILLER_300_1290 ();
 FILLCELL_X1 FILLER_300_1298 ();
 FILLCELL_X1 FILLER_300_1305 ();
 FILLCELL_X32 FILLER_300_1320 ();
 FILLCELL_X32 FILLER_300_1352 ();
 FILLCELL_X32 FILLER_300_1384 ();
 FILLCELL_X32 FILLER_300_1416 ();
 FILLCELL_X32 FILLER_300_1448 ();
 FILLCELL_X32 FILLER_300_1480 ();
 FILLCELL_X32 FILLER_300_1512 ();
 FILLCELL_X32 FILLER_300_1544 ();
 FILLCELL_X32 FILLER_300_1576 ();
 FILLCELL_X32 FILLER_300_1608 ();
 FILLCELL_X32 FILLER_300_1640 ();
 FILLCELL_X32 FILLER_300_1672 ();
 FILLCELL_X32 FILLER_300_1704 ();
 FILLCELL_X32 FILLER_300_1736 ();
 FILLCELL_X32 FILLER_300_1768 ();
 FILLCELL_X32 FILLER_300_1800 ();
 FILLCELL_X32 FILLER_300_1832 ();
 FILLCELL_X16 FILLER_300_1864 ();
 FILLCELL_X8 FILLER_300_1880 ();
 FILLCELL_X4 FILLER_300_1888 ();
 FILLCELL_X2 FILLER_300_1892 ();
 FILLCELL_X32 FILLER_300_1895 ();
 FILLCELL_X32 FILLER_300_1927 ();
 FILLCELL_X32 FILLER_300_1959 ();
 FILLCELL_X32 FILLER_300_1991 ();
 FILLCELL_X32 FILLER_300_2023 ();
 FILLCELL_X32 FILLER_300_2055 ();
 FILLCELL_X32 FILLER_300_2087 ();
 FILLCELL_X32 FILLER_300_2119 ();
 FILLCELL_X32 FILLER_300_2151 ();
 FILLCELL_X32 FILLER_300_2183 ();
 FILLCELL_X32 FILLER_300_2215 ();
 FILLCELL_X32 FILLER_300_2247 ();
 FILLCELL_X32 FILLER_300_2279 ();
 FILLCELL_X32 FILLER_300_2311 ();
 FILLCELL_X32 FILLER_300_2343 ();
 FILLCELL_X32 FILLER_300_2375 ();
 FILLCELL_X16 FILLER_300_2407 ();
 FILLCELL_X8 FILLER_300_2423 ();
 FILLCELL_X4 FILLER_300_2431 ();
 FILLCELL_X1 FILLER_300_2435 ();
 FILLCELL_X32 FILLER_301_1 ();
 FILLCELL_X32 FILLER_301_33 ();
 FILLCELL_X32 FILLER_301_65 ();
 FILLCELL_X32 FILLER_301_97 ();
 FILLCELL_X32 FILLER_301_129 ();
 FILLCELL_X32 FILLER_301_161 ();
 FILLCELL_X32 FILLER_301_193 ();
 FILLCELL_X32 FILLER_301_225 ();
 FILLCELL_X32 FILLER_301_257 ();
 FILLCELL_X32 FILLER_301_289 ();
 FILLCELL_X32 FILLER_301_321 ();
 FILLCELL_X32 FILLER_301_353 ();
 FILLCELL_X32 FILLER_301_385 ();
 FILLCELL_X32 FILLER_301_417 ();
 FILLCELL_X32 FILLER_301_449 ();
 FILLCELL_X32 FILLER_301_481 ();
 FILLCELL_X32 FILLER_301_513 ();
 FILLCELL_X32 FILLER_301_545 ();
 FILLCELL_X32 FILLER_301_577 ();
 FILLCELL_X32 FILLER_301_609 ();
 FILLCELL_X32 FILLER_301_641 ();
 FILLCELL_X32 FILLER_301_673 ();
 FILLCELL_X32 FILLER_301_705 ();
 FILLCELL_X32 FILLER_301_737 ();
 FILLCELL_X32 FILLER_301_769 ();
 FILLCELL_X32 FILLER_301_801 ();
 FILLCELL_X32 FILLER_301_833 ();
 FILLCELL_X32 FILLER_301_865 ();
 FILLCELL_X32 FILLER_301_897 ();
 FILLCELL_X32 FILLER_301_929 ();
 FILLCELL_X16 FILLER_301_961 ();
 FILLCELL_X8 FILLER_301_977 ();
 FILLCELL_X4 FILLER_301_985 ();
 FILLCELL_X1 FILLER_301_993 ();
 FILLCELL_X32 FILLER_301_1004 ();
 FILLCELL_X16 FILLER_301_1036 ();
 FILLCELL_X8 FILLER_301_1052 ();
 FILLCELL_X8 FILLER_301_1073 ();
 FILLCELL_X4 FILLER_301_1081 ();
 FILLCELL_X1 FILLER_301_1085 ();
 FILLCELL_X16 FILLER_301_1104 ();
 FILLCELL_X1 FILLER_301_1120 ();
 FILLCELL_X8 FILLER_301_1143 ();
 FILLCELL_X2 FILLER_301_1151 ();
 FILLCELL_X1 FILLER_301_1153 ();
 FILLCELL_X8 FILLER_301_1182 ();
 FILLCELL_X4 FILLER_301_1190 ();
 FILLCELL_X2 FILLER_301_1194 ();
 FILLCELL_X1 FILLER_301_1196 ();
 FILLCELL_X1 FILLER_301_1214 ();
 FILLCELL_X4 FILLER_301_1227 ();
 FILLCELL_X1 FILLER_301_1231 ();
 FILLCELL_X8 FILLER_301_1251 ();
 FILLCELL_X4 FILLER_301_1259 ();
 FILLCELL_X1 FILLER_301_1264 ();
 FILLCELL_X32 FILLER_301_1328 ();
 FILLCELL_X32 FILLER_301_1360 ();
 FILLCELL_X32 FILLER_301_1392 ();
 FILLCELL_X32 FILLER_301_1424 ();
 FILLCELL_X32 FILLER_301_1456 ();
 FILLCELL_X32 FILLER_301_1488 ();
 FILLCELL_X32 FILLER_301_1520 ();
 FILLCELL_X32 FILLER_301_1552 ();
 FILLCELL_X32 FILLER_301_1584 ();
 FILLCELL_X32 FILLER_301_1616 ();
 FILLCELL_X32 FILLER_301_1648 ();
 FILLCELL_X32 FILLER_301_1680 ();
 FILLCELL_X32 FILLER_301_1712 ();
 FILLCELL_X32 FILLER_301_1744 ();
 FILLCELL_X32 FILLER_301_1776 ();
 FILLCELL_X32 FILLER_301_1808 ();
 FILLCELL_X32 FILLER_301_1840 ();
 FILLCELL_X32 FILLER_301_1872 ();
 FILLCELL_X32 FILLER_301_1904 ();
 FILLCELL_X32 FILLER_301_1936 ();
 FILLCELL_X32 FILLER_301_1968 ();
 FILLCELL_X32 FILLER_301_2000 ();
 FILLCELL_X32 FILLER_301_2032 ();
 FILLCELL_X32 FILLER_301_2064 ();
 FILLCELL_X32 FILLER_301_2096 ();
 FILLCELL_X32 FILLER_301_2128 ();
 FILLCELL_X32 FILLER_301_2160 ();
 FILLCELL_X32 FILLER_301_2192 ();
 FILLCELL_X32 FILLER_301_2224 ();
 FILLCELL_X32 FILLER_301_2256 ();
 FILLCELL_X32 FILLER_301_2288 ();
 FILLCELL_X32 FILLER_301_2320 ();
 FILLCELL_X32 FILLER_301_2352 ();
 FILLCELL_X32 FILLER_301_2384 ();
 FILLCELL_X16 FILLER_301_2416 ();
 FILLCELL_X4 FILLER_301_2432 ();
 FILLCELL_X32 FILLER_302_1 ();
 FILLCELL_X32 FILLER_302_33 ();
 FILLCELL_X32 FILLER_302_65 ();
 FILLCELL_X32 FILLER_302_97 ();
 FILLCELL_X32 FILLER_302_129 ();
 FILLCELL_X32 FILLER_302_161 ();
 FILLCELL_X32 FILLER_302_193 ();
 FILLCELL_X32 FILLER_302_225 ();
 FILLCELL_X32 FILLER_302_257 ();
 FILLCELL_X32 FILLER_302_289 ();
 FILLCELL_X32 FILLER_302_321 ();
 FILLCELL_X32 FILLER_302_353 ();
 FILLCELL_X32 FILLER_302_385 ();
 FILLCELL_X32 FILLER_302_417 ();
 FILLCELL_X32 FILLER_302_449 ();
 FILLCELL_X32 FILLER_302_481 ();
 FILLCELL_X32 FILLER_302_513 ();
 FILLCELL_X32 FILLER_302_545 ();
 FILLCELL_X32 FILLER_302_577 ();
 FILLCELL_X16 FILLER_302_609 ();
 FILLCELL_X4 FILLER_302_625 ();
 FILLCELL_X2 FILLER_302_629 ();
 FILLCELL_X32 FILLER_302_632 ();
 FILLCELL_X32 FILLER_302_664 ();
 FILLCELL_X32 FILLER_302_696 ();
 FILLCELL_X32 FILLER_302_728 ();
 FILLCELL_X32 FILLER_302_760 ();
 FILLCELL_X32 FILLER_302_792 ();
 FILLCELL_X32 FILLER_302_824 ();
 FILLCELL_X32 FILLER_302_856 ();
 FILLCELL_X32 FILLER_302_888 ();
 FILLCELL_X32 FILLER_302_920 ();
 FILLCELL_X16 FILLER_302_952 ();
 FILLCELL_X8 FILLER_302_968 ();
 FILLCELL_X4 FILLER_302_976 ();
 FILLCELL_X2 FILLER_302_980 ();
 FILLCELL_X32 FILLER_302_1010 ();
 FILLCELL_X8 FILLER_302_1042 ();
 FILLCELL_X1 FILLER_302_1050 ();
 FILLCELL_X1 FILLER_302_1058 ();
 FILLCELL_X2 FILLER_302_1062 ();
 FILLCELL_X1 FILLER_302_1064 ();
 FILLCELL_X1 FILLER_302_1083 ();
 FILLCELL_X1 FILLER_302_1087 ();
 FILLCELL_X16 FILLER_302_1097 ();
 FILLCELL_X8 FILLER_302_1113 ();
 FILLCELL_X4 FILLER_302_1121 ();
 FILLCELL_X2 FILLER_302_1125 ();
 FILLCELL_X1 FILLER_302_1127 ();
 FILLCELL_X4 FILLER_302_1133 ();
 FILLCELL_X1 FILLER_302_1140 ();
 FILLCELL_X4 FILLER_302_1158 ();
 FILLCELL_X2 FILLER_302_1162 ();
 FILLCELL_X1 FILLER_302_1164 ();
 FILLCELL_X2 FILLER_302_1181 ();
 FILLCELL_X1 FILLER_302_1183 ();
 FILLCELL_X4 FILLER_302_1218 ();
 FILLCELL_X2 FILLER_302_1222 ();
 FILLCELL_X1 FILLER_302_1224 ();
 FILLCELL_X8 FILLER_302_1234 ();
 FILLCELL_X2 FILLER_302_1242 ();
 FILLCELL_X1 FILLER_302_1244 ();
 FILLCELL_X2 FILLER_302_1255 ();
 FILLCELL_X4 FILLER_302_1261 ();
 FILLCELL_X2 FILLER_302_1275 ();
 FILLCELL_X1 FILLER_302_1303 ();
 FILLCELL_X32 FILLER_302_1315 ();
 FILLCELL_X32 FILLER_302_1347 ();
 FILLCELL_X32 FILLER_302_1379 ();
 FILLCELL_X32 FILLER_302_1411 ();
 FILLCELL_X32 FILLER_302_1443 ();
 FILLCELL_X32 FILLER_302_1475 ();
 FILLCELL_X32 FILLER_302_1507 ();
 FILLCELL_X32 FILLER_302_1539 ();
 FILLCELL_X32 FILLER_302_1571 ();
 FILLCELL_X32 FILLER_302_1603 ();
 FILLCELL_X32 FILLER_302_1635 ();
 FILLCELL_X32 FILLER_302_1667 ();
 FILLCELL_X32 FILLER_302_1699 ();
 FILLCELL_X32 FILLER_302_1731 ();
 FILLCELL_X32 FILLER_302_1763 ();
 FILLCELL_X32 FILLER_302_1795 ();
 FILLCELL_X32 FILLER_302_1827 ();
 FILLCELL_X32 FILLER_302_1859 ();
 FILLCELL_X2 FILLER_302_1891 ();
 FILLCELL_X1 FILLER_302_1893 ();
 FILLCELL_X32 FILLER_302_1895 ();
 FILLCELL_X32 FILLER_302_1927 ();
 FILLCELL_X32 FILLER_302_1959 ();
 FILLCELL_X32 FILLER_302_1991 ();
 FILLCELL_X32 FILLER_302_2023 ();
 FILLCELL_X32 FILLER_302_2055 ();
 FILLCELL_X32 FILLER_302_2087 ();
 FILLCELL_X32 FILLER_302_2119 ();
 FILLCELL_X32 FILLER_302_2151 ();
 FILLCELL_X32 FILLER_302_2183 ();
 FILLCELL_X32 FILLER_302_2215 ();
 FILLCELL_X32 FILLER_302_2247 ();
 FILLCELL_X32 FILLER_302_2279 ();
 FILLCELL_X32 FILLER_302_2311 ();
 FILLCELL_X32 FILLER_302_2343 ();
 FILLCELL_X32 FILLER_302_2375 ();
 FILLCELL_X16 FILLER_302_2407 ();
 FILLCELL_X8 FILLER_302_2423 ();
 FILLCELL_X4 FILLER_302_2431 ();
 FILLCELL_X1 FILLER_302_2435 ();
 FILLCELL_X32 FILLER_303_1 ();
 FILLCELL_X32 FILLER_303_33 ();
 FILLCELL_X32 FILLER_303_65 ();
 FILLCELL_X32 FILLER_303_97 ();
 FILLCELL_X32 FILLER_303_129 ();
 FILLCELL_X32 FILLER_303_161 ();
 FILLCELL_X32 FILLER_303_193 ();
 FILLCELL_X32 FILLER_303_225 ();
 FILLCELL_X32 FILLER_303_257 ();
 FILLCELL_X32 FILLER_303_289 ();
 FILLCELL_X32 FILLER_303_321 ();
 FILLCELL_X32 FILLER_303_353 ();
 FILLCELL_X32 FILLER_303_385 ();
 FILLCELL_X32 FILLER_303_417 ();
 FILLCELL_X32 FILLER_303_449 ();
 FILLCELL_X32 FILLER_303_481 ();
 FILLCELL_X32 FILLER_303_513 ();
 FILLCELL_X32 FILLER_303_545 ();
 FILLCELL_X32 FILLER_303_577 ();
 FILLCELL_X32 FILLER_303_609 ();
 FILLCELL_X32 FILLER_303_641 ();
 FILLCELL_X32 FILLER_303_673 ();
 FILLCELL_X32 FILLER_303_705 ();
 FILLCELL_X32 FILLER_303_737 ();
 FILLCELL_X32 FILLER_303_769 ();
 FILLCELL_X32 FILLER_303_801 ();
 FILLCELL_X32 FILLER_303_833 ();
 FILLCELL_X32 FILLER_303_865 ();
 FILLCELL_X32 FILLER_303_897 ();
 FILLCELL_X16 FILLER_303_929 ();
 FILLCELL_X8 FILLER_303_945 ();
 FILLCELL_X4 FILLER_303_953 ();
 FILLCELL_X2 FILLER_303_957 ();
 FILLCELL_X1 FILLER_303_959 ();
 FILLCELL_X4 FILLER_303_979 ();
 FILLCELL_X1 FILLER_303_983 ();
 FILLCELL_X2 FILLER_303_988 ();
 FILLCELL_X2 FILLER_303_998 ();
 FILLCELL_X1 FILLER_303_1000 ();
 FILLCELL_X2 FILLER_303_1005 ();
 FILLCELL_X1 FILLER_303_1007 ();
 FILLCELL_X4 FILLER_303_1015 ();
 FILLCELL_X2 FILLER_303_1019 ();
 FILLCELL_X4 FILLER_303_1036 ();
 FILLCELL_X8 FILLER_303_1058 ();
 FILLCELL_X2 FILLER_303_1066 ();
 FILLCELL_X1 FILLER_303_1068 ();
 FILLCELL_X4 FILLER_303_1075 ();
 FILLCELL_X32 FILLER_303_1092 ();
 FILLCELL_X1 FILLER_303_1124 ();
 FILLCELL_X2 FILLER_303_1140 ();
 FILLCELL_X2 FILLER_303_1152 ();
 FILLCELL_X32 FILLER_303_1183 ();
 FILLCELL_X4 FILLER_303_1215 ();
 FILLCELL_X8 FILLER_303_1223 ();
 FILLCELL_X4 FILLER_303_1231 ();
 FILLCELL_X2 FILLER_303_1235 ();
 FILLCELL_X2 FILLER_303_1248 ();
 FILLCELL_X1 FILLER_303_1262 ();
 FILLCELL_X8 FILLER_303_1264 ();
 FILLCELL_X4 FILLER_303_1272 ();
 FILLCELL_X2 FILLER_303_1276 ();
 FILLCELL_X8 FILLER_303_1281 ();
 FILLCELL_X4 FILLER_303_1289 ();
 FILLCELL_X8 FILLER_303_1296 ();
 FILLCELL_X1 FILLER_303_1324 ();
 FILLCELL_X32 FILLER_303_1329 ();
 FILLCELL_X32 FILLER_303_1361 ();
 FILLCELL_X32 FILLER_303_1393 ();
 FILLCELL_X32 FILLER_303_1425 ();
 FILLCELL_X32 FILLER_303_1457 ();
 FILLCELL_X32 FILLER_303_1489 ();
 FILLCELL_X32 FILLER_303_1521 ();
 FILLCELL_X32 FILLER_303_1553 ();
 FILLCELL_X32 FILLER_303_1585 ();
 FILLCELL_X32 FILLER_303_1617 ();
 FILLCELL_X32 FILLER_303_1649 ();
 FILLCELL_X32 FILLER_303_1681 ();
 FILLCELL_X32 FILLER_303_1713 ();
 FILLCELL_X32 FILLER_303_1745 ();
 FILLCELL_X32 FILLER_303_1777 ();
 FILLCELL_X32 FILLER_303_1809 ();
 FILLCELL_X32 FILLER_303_1841 ();
 FILLCELL_X32 FILLER_303_1873 ();
 FILLCELL_X32 FILLER_303_1905 ();
 FILLCELL_X32 FILLER_303_1937 ();
 FILLCELL_X32 FILLER_303_1969 ();
 FILLCELL_X32 FILLER_303_2001 ();
 FILLCELL_X32 FILLER_303_2033 ();
 FILLCELL_X32 FILLER_303_2065 ();
 FILLCELL_X32 FILLER_303_2097 ();
 FILLCELL_X32 FILLER_303_2129 ();
 FILLCELL_X32 FILLER_303_2161 ();
 FILLCELL_X32 FILLER_303_2193 ();
 FILLCELL_X32 FILLER_303_2225 ();
 FILLCELL_X32 FILLER_303_2257 ();
 FILLCELL_X32 FILLER_303_2289 ();
 FILLCELL_X32 FILLER_303_2321 ();
 FILLCELL_X32 FILLER_303_2353 ();
 FILLCELL_X32 FILLER_303_2385 ();
 FILLCELL_X16 FILLER_303_2417 ();
 FILLCELL_X2 FILLER_303_2433 ();
 FILLCELL_X1 FILLER_303_2435 ();
 FILLCELL_X32 FILLER_304_1 ();
 FILLCELL_X32 FILLER_304_33 ();
 FILLCELL_X32 FILLER_304_65 ();
 FILLCELL_X32 FILLER_304_97 ();
 FILLCELL_X32 FILLER_304_129 ();
 FILLCELL_X32 FILLER_304_161 ();
 FILLCELL_X32 FILLER_304_193 ();
 FILLCELL_X32 FILLER_304_225 ();
 FILLCELL_X32 FILLER_304_257 ();
 FILLCELL_X32 FILLER_304_289 ();
 FILLCELL_X32 FILLER_304_321 ();
 FILLCELL_X32 FILLER_304_353 ();
 FILLCELL_X32 FILLER_304_385 ();
 FILLCELL_X32 FILLER_304_417 ();
 FILLCELL_X32 FILLER_304_449 ();
 FILLCELL_X32 FILLER_304_481 ();
 FILLCELL_X32 FILLER_304_513 ();
 FILLCELL_X32 FILLER_304_545 ();
 FILLCELL_X32 FILLER_304_577 ();
 FILLCELL_X16 FILLER_304_609 ();
 FILLCELL_X4 FILLER_304_625 ();
 FILLCELL_X2 FILLER_304_629 ();
 FILLCELL_X32 FILLER_304_632 ();
 FILLCELL_X32 FILLER_304_664 ();
 FILLCELL_X32 FILLER_304_696 ();
 FILLCELL_X32 FILLER_304_728 ();
 FILLCELL_X32 FILLER_304_760 ();
 FILLCELL_X32 FILLER_304_792 ();
 FILLCELL_X32 FILLER_304_824 ();
 FILLCELL_X32 FILLER_304_856 ();
 FILLCELL_X32 FILLER_304_888 ();
 FILLCELL_X32 FILLER_304_920 ();
 FILLCELL_X4 FILLER_304_952 ();
 FILLCELL_X1 FILLER_304_956 ();
 FILLCELL_X16 FILLER_304_959 ();
 FILLCELL_X8 FILLER_304_992 ();
 FILLCELL_X4 FILLER_304_1000 ();
 FILLCELL_X1 FILLER_304_1004 ();
 FILLCELL_X16 FILLER_304_1049 ();
 FILLCELL_X8 FILLER_304_1065 ();
 FILLCELL_X2 FILLER_304_1099 ();
 FILLCELL_X2 FILLER_304_1105 ();
 FILLCELL_X1 FILLER_304_1107 ();
 FILLCELL_X16 FILLER_304_1113 ();
 FILLCELL_X4 FILLER_304_1129 ();
 FILLCELL_X2 FILLER_304_1133 ();
 FILLCELL_X16 FILLER_304_1141 ();
 FILLCELL_X8 FILLER_304_1157 ();
 FILLCELL_X2 FILLER_304_1165 ();
 FILLCELL_X8 FILLER_304_1179 ();
 FILLCELL_X1 FILLER_304_1187 ();
 FILLCELL_X4 FILLER_304_1205 ();
 FILLCELL_X2 FILLER_304_1220 ();
 FILLCELL_X4 FILLER_304_1235 ();
 FILLCELL_X1 FILLER_304_1239 ();
 FILLCELL_X2 FILLER_304_1245 ();
 FILLCELL_X1 FILLER_304_1247 ();
 FILLCELL_X8 FILLER_304_1252 ();
 FILLCELL_X4 FILLER_304_1260 ();
 FILLCELL_X2 FILLER_304_1264 ();
 FILLCELL_X2 FILLER_304_1279 ();
 FILLCELL_X1 FILLER_304_1281 ();
 FILLCELL_X8 FILLER_304_1285 ();
 FILLCELL_X2 FILLER_304_1300 ();
 FILLCELL_X1 FILLER_304_1302 ();
 FILLCELL_X32 FILLER_304_1328 ();
 FILLCELL_X32 FILLER_304_1360 ();
 FILLCELL_X32 FILLER_304_1392 ();
 FILLCELL_X32 FILLER_304_1424 ();
 FILLCELL_X32 FILLER_304_1456 ();
 FILLCELL_X32 FILLER_304_1488 ();
 FILLCELL_X32 FILLER_304_1520 ();
 FILLCELL_X32 FILLER_304_1552 ();
 FILLCELL_X32 FILLER_304_1584 ();
 FILLCELL_X32 FILLER_304_1616 ();
 FILLCELL_X32 FILLER_304_1648 ();
 FILLCELL_X32 FILLER_304_1680 ();
 FILLCELL_X32 FILLER_304_1712 ();
 FILLCELL_X32 FILLER_304_1744 ();
 FILLCELL_X32 FILLER_304_1776 ();
 FILLCELL_X32 FILLER_304_1808 ();
 FILLCELL_X32 FILLER_304_1840 ();
 FILLCELL_X16 FILLER_304_1872 ();
 FILLCELL_X4 FILLER_304_1888 ();
 FILLCELL_X2 FILLER_304_1892 ();
 FILLCELL_X32 FILLER_304_1895 ();
 FILLCELL_X32 FILLER_304_1927 ();
 FILLCELL_X32 FILLER_304_1959 ();
 FILLCELL_X32 FILLER_304_1991 ();
 FILLCELL_X32 FILLER_304_2023 ();
 FILLCELL_X32 FILLER_304_2055 ();
 FILLCELL_X32 FILLER_304_2087 ();
 FILLCELL_X32 FILLER_304_2119 ();
 FILLCELL_X32 FILLER_304_2151 ();
 FILLCELL_X32 FILLER_304_2183 ();
 FILLCELL_X32 FILLER_304_2215 ();
 FILLCELL_X32 FILLER_304_2247 ();
 FILLCELL_X32 FILLER_304_2279 ();
 FILLCELL_X32 FILLER_304_2311 ();
 FILLCELL_X32 FILLER_304_2343 ();
 FILLCELL_X32 FILLER_304_2375 ();
 FILLCELL_X16 FILLER_304_2407 ();
 FILLCELL_X8 FILLER_304_2423 ();
 FILLCELL_X4 FILLER_304_2431 ();
 FILLCELL_X1 FILLER_304_2435 ();
 FILLCELL_X32 FILLER_305_1 ();
 FILLCELL_X32 FILLER_305_33 ();
 FILLCELL_X32 FILLER_305_65 ();
 FILLCELL_X32 FILLER_305_97 ();
 FILLCELL_X32 FILLER_305_129 ();
 FILLCELL_X32 FILLER_305_161 ();
 FILLCELL_X32 FILLER_305_193 ();
 FILLCELL_X32 FILLER_305_225 ();
 FILLCELL_X32 FILLER_305_257 ();
 FILLCELL_X32 FILLER_305_289 ();
 FILLCELL_X32 FILLER_305_321 ();
 FILLCELL_X32 FILLER_305_353 ();
 FILLCELL_X32 FILLER_305_385 ();
 FILLCELL_X32 FILLER_305_417 ();
 FILLCELL_X32 FILLER_305_449 ();
 FILLCELL_X32 FILLER_305_481 ();
 FILLCELL_X32 FILLER_305_513 ();
 FILLCELL_X32 FILLER_305_545 ();
 FILLCELL_X32 FILLER_305_577 ();
 FILLCELL_X32 FILLER_305_609 ();
 FILLCELL_X32 FILLER_305_641 ();
 FILLCELL_X32 FILLER_305_673 ();
 FILLCELL_X32 FILLER_305_705 ();
 FILLCELL_X32 FILLER_305_737 ();
 FILLCELL_X32 FILLER_305_769 ();
 FILLCELL_X32 FILLER_305_801 ();
 FILLCELL_X32 FILLER_305_833 ();
 FILLCELL_X32 FILLER_305_865 ();
 FILLCELL_X32 FILLER_305_897 ();
 FILLCELL_X16 FILLER_305_929 ();
 FILLCELL_X8 FILLER_305_945 ();
 FILLCELL_X1 FILLER_305_953 ();
 FILLCELL_X16 FILLER_305_956 ();
 FILLCELL_X2 FILLER_305_972 ();
 FILLCELL_X16 FILLER_305_988 ();
 FILLCELL_X8 FILLER_305_1004 ();
 FILLCELL_X1 FILLER_305_1012 ();
 FILLCELL_X2 FILLER_305_1018 ();
 FILLCELL_X1 FILLER_305_1020 ();
 FILLCELL_X1 FILLER_305_1038 ();
 FILLCELL_X16 FILLER_305_1053 ();
 FILLCELL_X1 FILLER_305_1069 ();
 FILLCELL_X8 FILLER_305_1072 ();
 FILLCELL_X4 FILLER_305_1080 ();
 FILLCELL_X2 FILLER_305_1084 ();
 FILLCELL_X1 FILLER_305_1088 ();
 FILLCELL_X32 FILLER_305_1100 ();
 FILLCELL_X2 FILLER_305_1132 ();
 FILLCELL_X1 FILLER_305_1134 ();
 FILLCELL_X16 FILLER_305_1144 ();
 FILLCELL_X8 FILLER_305_1160 ();
 FILLCELL_X4 FILLER_305_1168 ();
 FILLCELL_X1 FILLER_305_1172 ();
 FILLCELL_X16 FILLER_305_1195 ();
 FILLCELL_X4 FILLER_305_1211 ();
 FILLCELL_X2 FILLER_305_1215 ();
 FILLCELL_X16 FILLER_305_1230 ();
 FILLCELL_X8 FILLER_305_1246 ();
 FILLCELL_X2 FILLER_305_1254 ();
 FILLCELL_X1 FILLER_305_1256 ();
 FILLCELL_X2 FILLER_305_1260 ();
 FILLCELL_X1 FILLER_305_1262 ();
 FILLCELL_X1 FILLER_305_1264 ();
 FILLCELL_X4 FILLER_305_1268 ();
 FILLCELL_X2 FILLER_305_1272 ();
 FILLCELL_X1 FILLER_305_1274 ();
 FILLCELL_X8 FILLER_305_1278 ();
 FILLCELL_X1 FILLER_305_1286 ();
 FILLCELL_X4 FILLER_305_1297 ();
 FILLCELL_X1 FILLER_305_1301 ();
 FILLCELL_X2 FILLER_305_1320 ();
 FILLCELL_X1 FILLER_305_1322 ();
 FILLCELL_X1 FILLER_305_1326 ();
 FILLCELL_X32 FILLER_305_1339 ();
 FILLCELL_X32 FILLER_305_1371 ();
 FILLCELL_X32 FILLER_305_1403 ();
 FILLCELL_X32 FILLER_305_1435 ();
 FILLCELL_X32 FILLER_305_1467 ();
 FILLCELL_X32 FILLER_305_1499 ();
 FILLCELL_X32 FILLER_305_1531 ();
 FILLCELL_X32 FILLER_305_1563 ();
 FILLCELL_X32 FILLER_305_1595 ();
 FILLCELL_X32 FILLER_305_1627 ();
 FILLCELL_X32 FILLER_305_1659 ();
 FILLCELL_X32 FILLER_305_1691 ();
 FILLCELL_X32 FILLER_305_1723 ();
 FILLCELL_X32 FILLER_305_1755 ();
 FILLCELL_X32 FILLER_305_1787 ();
 FILLCELL_X32 FILLER_305_1819 ();
 FILLCELL_X32 FILLER_305_1851 ();
 FILLCELL_X32 FILLER_305_1883 ();
 FILLCELL_X32 FILLER_305_1915 ();
 FILLCELL_X32 FILLER_305_1947 ();
 FILLCELL_X32 FILLER_305_1979 ();
 FILLCELL_X32 FILLER_305_2011 ();
 FILLCELL_X32 FILLER_305_2043 ();
 FILLCELL_X32 FILLER_305_2075 ();
 FILLCELL_X32 FILLER_305_2107 ();
 FILLCELL_X32 FILLER_305_2139 ();
 FILLCELL_X32 FILLER_305_2171 ();
 FILLCELL_X32 FILLER_305_2203 ();
 FILLCELL_X32 FILLER_305_2235 ();
 FILLCELL_X32 FILLER_305_2267 ();
 FILLCELL_X32 FILLER_305_2299 ();
 FILLCELL_X32 FILLER_305_2331 ();
 FILLCELL_X32 FILLER_305_2363 ();
 FILLCELL_X32 FILLER_305_2395 ();
 FILLCELL_X8 FILLER_305_2427 ();
 FILLCELL_X1 FILLER_305_2435 ();
 FILLCELL_X32 FILLER_306_1 ();
 FILLCELL_X32 FILLER_306_33 ();
 FILLCELL_X32 FILLER_306_65 ();
 FILLCELL_X32 FILLER_306_97 ();
 FILLCELL_X32 FILLER_306_129 ();
 FILLCELL_X32 FILLER_306_161 ();
 FILLCELL_X32 FILLER_306_193 ();
 FILLCELL_X32 FILLER_306_225 ();
 FILLCELL_X32 FILLER_306_257 ();
 FILLCELL_X32 FILLER_306_289 ();
 FILLCELL_X32 FILLER_306_321 ();
 FILLCELL_X32 FILLER_306_353 ();
 FILLCELL_X32 FILLER_306_385 ();
 FILLCELL_X32 FILLER_306_417 ();
 FILLCELL_X32 FILLER_306_449 ();
 FILLCELL_X32 FILLER_306_481 ();
 FILLCELL_X32 FILLER_306_513 ();
 FILLCELL_X32 FILLER_306_545 ();
 FILLCELL_X32 FILLER_306_577 ();
 FILLCELL_X16 FILLER_306_609 ();
 FILLCELL_X4 FILLER_306_625 ();
 FILLCELL_X2 FILLER_306_629 ();
 FILLCELL_X32 FILLER_306_632 ();
 FILLCELL_X32 FILLER_306_664 ();
 FILLCELL_X32 FILLER_306_696 ();
 FILLCELL_X32 FILLER_306_728 ();
 FILLCELL_X32 FILLER_306_760 ();
 FILLCELL_X32 FILLER_306_792 ();
 FILLCELL_X32 FILLER_306_824 ();
 FILLCELL_X32 FILLER_306_856 ();
 FILLCELL_X2 FILLER_306_888 ();
 FILLCELL_X16 FILLER_306_894 ();
 FILLCELL_X4 FILLER_306_910 ();
 FILLCELL_X8 FILLER_306_922 ();
 FILLCELL_X4 FILLER_306_930 ();
 FILLCELL_X1 FILLER_306_934 ();
 FILLCELL_X2 FILLER_306_953 ();
 FILLCELL_X1 FILLER_306_955 ();
 FILLCELL_X32 FILLER_306_966 ();
 FILLCELL_X16 FILLER_306_998 ();
 FILLCELL_X8 FILLER_306_1014 ();
 FILLCELL_X2 FILLER_306_1022 ();
 FILLCELL_X16 FILLER_306_1026 ();
 FILLCELL_X8 FILLER_306_1042 ();
 FILLCELL_X1 FILLER_306_1050 ();
 FILLCELL_X8 FILLER_306_1068 ();
 FILLCELL_X1 FILLER_306_1076 ();
 FILLCELL_X1 FILLER_306_1080 ();
 FILLCELL_X2 FILLER_306_1102 ();
 FILLCELL_X1 FILLER_306_1114 ();
 FILLCELL_X32 FILLER_306_1124 ();
 FILLCELL_X32 FILLER_306_1156 ();
 FILLCELL_X16 FILLER_306_1188 ();
 FILLCELL_X4 FILLER_306_1204 ();
 FILLCELL_X2 FILLER_306_1208 ();
 FILLCELL_X1 FILLER_306_1210 ();
 FILLCELL_X2 FILLER_306_1234 ();
 FILLCELL_X2 FILLER_306_1238 ();
 FILLCELL_X1 FILLER_306_1256 ();
 FILLCELL_X1 FILLER_306_1261 ();
 FILLCELL_X1 FILLER_306_1273 ();
 FILLCELL_X2 FILLER_306_1281 ();
 FILLCELL_X2 FILLER_306_1302 ();
 FILLCELL_X1 FILLER_306_1325 ();
 FILLCELL_X32 FILLER_306_1330 ();
 FILLCELL_X32 FILLER_306_1362 ();
 FILLCELL_X32 FILLER_306_1394 ();
 FILLCELL_X32 FILLER_306_1426 ();
 FILLCELL_X32 FILLER_306_1458 ();
 FILLCELL_X32 FILLER_306_1490 ();
 FILLCELL_X32 FILLER_306_1522 ();
 FILLCELL_X32 FILLER_306_1554 ();
 FILLCELL_X32 FILLER_306_1586 ();
 FILLCELL_X32 FILLER_306_1618 ();
 FILLCELL_X32 FILLER_306_1650 ();
 FILLCELL_X32 FILLER_306_1682 ();
 FILLCELL_X32 FILLER_306_1714 ();
 FILLCELL_X32 FILLER_306_1746 ();
 FILLCELL_X32 FILLER_306_1778 ();
 FILLCELL_X32 FILLER_306_1810 ();
 FILLCELL_X32 FILLER_306_1842 ();
 FILLCELL_X16 FILLER_306_1874 ();
 FILLCELL_X4 FILLER_306_1890 ();
 FILLCELL_X32 FILLER_306_1895 ();
 FILLCELL_X32 FILLER_306_1927 ();
 FILLCELL_X32 FILLER_306_1959 ();
 FILLCELL_X32 FILLER_306_1991 ();
 FILLCELL_X32 FILLER_306_2023 ();
 FILLCELL_X32 FILLER_306_2055 ();
 FILLCELL_X32 FILLER_306_2087 ();
 FILLCELL_X32 FILLER_306_2119 ();
 FILLCELL_X32 FILLER_306_2151 ();
 FILLCELL_X32 FILLER_306_2183 ();
 FILLCELL_X32 FILLER_306_2215 ();
 FILLCELL_X32 FILLER_306_2247 ();
 FILLCELL_X32 FILLER_306_2279 ();
 FILLCELL_X32 FILLER_306_2311 ();
 FILLCELL_X32 FILLER_306_2343 ();
 FILLCELL_X32 FILLER_306_2375 ();
 FILLCELL_X16 FILLER_306_2407 ();
 FILLCELL_X8 FILLER_306_2423 ();
 FILLCELL_X4 FILLER_306_2431 ();
 FILLCELL_X1 FILLER_306_2435 ();
 FILLCELL_X32 FILLER_307_1 ();
 FILLCELL_X32 FILLER_307_33 ();
 FILLCELL_X32 FILLER_307_65 ();
 FILLCELL_X32 FILLER_307_97 ();
 FILLCELL_X32 FILLER_307_129 ();
 FILLCELL_X32 FILLER_307_161 ();
 FILLCELL_X32 FILLER_307_193 ();
 FILLCELL_X32 FILLER_307_225 ();
 FILLCELL_X32 FILLER_307_257 ();
 FILLCELL_X32 FILLER_307_289 ();
 FILLCELL_X32 FILLER_307_321 ();
 FILLCELL_X32 FILLER_307_353 ();
 FILLCELL_X32 FILLER_307_385 ();
 FILLCELL_X32 FILLER_307_417 ();
 FILLCELL_X32 FILLER_307_449 ();
 FILLCELL_X32 FILLER_307_481 ();
 FILLCELL_X32 FILLER_307_513 ();
 FILLCELL_X32 FILLER_307_545 ();
 FILLCELL_X32 FILLER_307_577 ();
 FILLCELL_X32 FILLER_307_609 ();
 FILLCELL_X32 FILLER_307_641 ();
 FILLCELL_X32 FILLER_307_673 ();
 FILLCELL_X32 FILLER_307_705 ();
 FILLCELL_X32 FILLER_307_737 ();
 FILLCELL_X32 FILLER_307_769 ();
 FILLCELL_X32 FILLER_307_801 ();
 FILLCELL_X32 FILLER_307_833 ();
 FILLCELL_X32 FILLER_307_865 ();
 FILLCELL_X16 FILLER_307_897 ();
 FILLCELL_X8 FILLER_307_913 ();
 FILLCELL_X4 FILLER_307_921 ();
 FILLCELL_X2 FILLER_307_925 ();
 FILLCELL_X1 FILLER_307_927 ();
 FILLCELL_X8 FILLER_307_930 ();
 FILLCELL_X4 FILLER_307_938 ();
 FILLCELL_X2 FILLER_307_942 ();
 FILLCELL_X8 FILLER_307_946 ();
 FILLCELL_X8 FILLER_307_958 ();
 FILLCELL_X4 FILLER_307_966 ();
 FILLCELL_X2 FILLER_307_970 ();
 FILLCELL_X2 FILLER_307_976 ();
 FILLCELL_X1 FILLER_307_978 ();
 FILLCELL_X16 FILLER_307_991 ();
 FILLCELL_X2 FILLER_307_1007 ();
 FILLCELL_X1 FILLER_307_1009 ();
 FILLCELL_X4 FILLER_307_1014 ();
 FILLCELL_X2 FILLER_307_1018 ();
 FILLCELL_X1 FILLER_307_1020 ();
 FILLCELL_X2 FILLER_307_1046 ();
 FILLCELL_X1 FILLER_307_1048 ();
 FILLCELL_X4 FILLER_307_1062 ();
 FILLCELL_X32 FILLER_307_1090 ();
 FILLCELL_X8 FILLER_307_1122 ();
 FILLCELL_X1 FILLER_307_1130 ();
 FILLCELL_X32 FILLER_307_1152 ();
 FILLCELL_X16 FILLER_307_1184 ();
 FILLCELL_X8 FILLER_307_1200 ();
 FILLCELL_X4 FILLER_307_1208 ();
 FILLCELL_X2 FILLER_307_1212 ();
 FILLCELL_X1 FILLER_307_1214 ();
 FILLCELL_X1 FILLER_307_1242 ();
 FILLCELL_X1 FILLER_307_1248 ();
 FILLCELL_X2 FILLER_307_1260 ();
 FILLCELL_X1 FILLER_307_1262 ();
 FILLCELL_X1 FILLER_307_1264 ();
 FILLCELL_X1 FILLER_307_1272 ();
 FILLCELL_X4 FILLER_307_1276 ();
 FILLCELL_X4 FILLER_307_1287 ();
 FILLCELL_X2 FILLER_307_1291 ();
 FILLCELL_X4 FILLER_307_1296 ();
 FILLCELL_X2 FILLER_307_1300 ();
 FILLCELL_X2 FILLER_307_1309 ();
 FILLCELL_X1 FILLER_307_1311 ();
 FILLCELL_X2 FILLER_307_1322 ();
 FILLCELL_X32 FILLER_307_1335 ();
 FILLCELL_X32 FILLER_307_1367 ();
 FILLCELL_X32 FILLER_307_1399 ();
 FILLCELL_X32 FILLER_307_1431 ();
 FILLCELL_X32 FILLER_307_1463 ();
 FILLCELL_X32 FILLER_307_1495 ();
 FILLCELL_X32 FILLER_307_1527 ();
 FILLCELL_X32 FILLER_307_1559 ();
 FILLCELL_X32 FILLER_307_1591 ();
 FILLCELL_X32 FILLER_307_1623 ();
 FILLCELL_X32 FILLER_307_1655 ();
 FILLCELL_X32 FILLER_307_1687 ();
 FILLCELL_X32 FILLER_307_1719 ();
 FILLCELL_X32 FILLER_307_1751 ();
 FILLCELL_X32 FILLER_307_1783 ();
 FILLCELL_X32 FILLER_307_1815 ();
 FILLCELL_X32 FILLER_307_1847 ();
 FILLCELL_X32 FILLER_307_1879 ();
 FILLCELL_X32 FILLER_307_1911 ();
 FILLCELL_X32 FILLER_307_1943 ();
 FILLCELL_X32 FILLER_307_1975 ();
 FILLCELL_X32 FILLER_307_2007 ();
 FILLCELL_X32 FILLER_307_2039 ();
 FILLCELL_X32 FILLER_307_2071 ();
 FILLCELL_X32 FILLER_307_2103 ();
 FILLCELL_X32 FILLER_307_2135 ();
 FILLCELL_X32 FILLER_307_2167 ();
 FILLCELL_X32 FILLER_307_2199 ();
 FILLCELL_X32 FILLER_307_2231 ();
 FILLCELL_X32 FILLER_307_2263 ();
 FILLCELL_X32 FILLER_307_2295 ();
 FILLCELL_X32 FILLER_307_2327 ();
 FILLCELL_X32 FILLER_307_2359 ();
 FILLCELL_X32 FILLER_307_2391 ();
 FILLCELL_X8 FILLER_307_2423 ();
 FILLCELL_X4 FILLER_307_2431 ();
 FILLCELL_X1 FILLER_307_2435 ();
 FILLCELL_X32 FILLER_308_1 ();
 FILLCELL_X32 FILLER_308_33 ();
 FILLCELL_X32 FILLER_308_65 ();
 FILLCELL_X32 FILLER_308_97 ();
 FILLCELL_X32 FILLER_308_129 ();
 FILLCELL_X32 FILLER_308_161 ();
 FILLCELL_X32 FILLER_308_193 ();
 FILLCELL_X32 FILLER_308_225 ();
 FILLCELL_X32 FILLER_308_257 ();
 FILLCELL_X32 FILLER_308_289 ();
 FILLCELL_X32 FILLER_308_321 ();
 FILLCELL_X32 FILLER_308_353 ();
 FILLCELL_X32 FILLER_308_385 ();
 FILLCELL_X32 FILLER_308_417 ();
 FILLCELL_X32 FILLER_308_449 ();
 FILLCELL_X32 FILLER_308_481 ();
 FILLCELL_X32 FILLER_308_513 ();
 FILLCELL_X32 FILLER_308_545 ();
 FILLCELL_X32 FILLER_308_577 ();
 FILLCELL_X16 FILLER_308_609 ();
 FILLCELL_X4 FILLER_308_625 ();
 FILLCELL_X2 FILLER_308_629 ();
 FILLCELL_X32 FILLER_308_632 ();
 FILLCELL_X32 FILLER_308_664 ();
 FILLCELL_X32 FILLER_308_696 ();
 FILLCELL_X32 FILLER_308_728 ();
 FILLCELL_X32 FILLER_308_760 ();
 FILLCELL_X32 FILLER_308_792 ();
 FILLCELL_X32 FILLER_308_824 ();
 FILLCELL_X32 FILLER_308_856 ();
 FILLCELL_X32 FILLER_308_888 ();
 FILLCELL_X8 FILLER_308_920 ();
 FILLCELL_X1 FILLER_308_928 ();
 FILLCELL_X16 FILLER_308_945 ();
 FILLCELL_X8 FILLER_308_961 ();
 FILLCELL_X4 FILLER_308_969 ();
 FILLCELL_X1 FILLER_308_973 ();
 FILLCELL_X8 FILLER_308_984 ();
 FILLCELL_X2 FILLER_308_992 ();
 FILLCELL_X1 FILLER_308_994 ();
 FILLCELL_X1 FILLER_308_1002 ();
 FILLCELL_X2 FILLER_308_1008 ();
 FILLCELL_X2 FILLER_308_1014 ();
 FILLCELL_X32 FILLER_308_1034 ();
 FILLCELL_X8 FILLER_308_1066 ();
 FILLCELL_X4 FILLER_308_1074 ();
 FILLCELL_X2 FILLER_308_1078 ();
 FILLCELL_X16 FILLER_308_1087 ();
 FILLCELL_X8 FILLER_308_1103 ();
 FILLCELL_X2 FILLER_308_1111 ();
 FILLCELL_X4 FILLER_308_1118 ();
 FILLCELL_X4 FILLER_308_1129 ();
 FILLCELL_X2 FILLER_308_1133 ();
 FILLCELL_X4 FILLER_308_1151 ();
 FILLCELL_X1 FILLER_308_1155 ();
 FILLCELL_X4 FILLER_308_1163 ();
 FILLCELL_X2 FILLER_308_1167 ();
 FILLCELL_X1 FILLER_308_1169 ();
 FILLCELL_X1 FILLER_308_1180 ();
 FILLCELL_X2 FILLER_308_1191 ();
 FILLCELL_X1 FILLER_308_1193 ();
 FILLCELL_X8 FILLER_308_1199 ();
 FILLCELL_X2 FILLER_308_1215 ();
 FILLCELL_X1 FILLER_308_1247 ();
 FILLCELL_X32 FILLER_308_1268 ();
 FILLCELL_X8 FILLER_308_1300 ();
 FILLCELL_X2 FILLER_308_1317 ();
 FILLCELL_X32 FILLER_308_1336 ();
 FILLCELL_X32 FILLER_308_1368 ();
 FILLCELL_X32 FILLER_308_1400 ();
 FILLCELL_X32 FILLER_308_1432 ();
 FILLCELL_X32 FILLER_308_1464 ();
 FILLCELL_X32 FILLER_308_1496 ();
 FILLCELL_X32 FILLER_308_1528 ();
 FILLCELL_X32 FILLER_308_1560 ();
 FILLCELL_X32 FILLER_308_1592 ();
 FILLCELL_X32 FILLER_308_1624 ();
 FILLCELL_X32 FILLER_308_1656 ();
 FILLCELL_X32 FILLER_308_1688 ();
 FILLCELL_X32 FILLER_308_1720 ();
 FILLCELL_X32 FILLER_308_1752 ();
 FILLCELL_X32 FILLER_308_1784 ();
 FILLCELL_X32 FILLER_308_1816 ();
 FILLCELL_X32 FILLER_308_1848 ();
 FILLCELL_X8 FILLER_308_1880 ();
 FILLCELL_X4 FILLER_308_1888 ();
 FILLCELL_X2 FILLER_308_1892 ();
 FILLCELL_X32 FILLER_308_1895 ();
 FILLCELL_X32 FILLER_308_1927 ();
 FILLCELL_X32 FILLER_308_1959 ();
 FILLCELL_X32 FILLER_308_1991 ();
 FILLCELL_X32 FILLER_308_2023 ();
 FILLCELL_X32 FILLER_308_2055 ();
 FILLCELL_X32 FILLER_308_2087 ();
 FILLCELL_X32 FILLER_308_2119 ();
 FILLCELL_X32 FILLER_308_2151 ();
 FILLCELL_X32 FILLER_308_2183 ();
 FILLCELL_X32 FILLER_308_2215 ();
 FILLCELL_X32 FILLER_308_2247 ();
 FILLCELL_X32 FILLER_308_2279 ();
 FILLCELL_X32 FILLER_308_2311 ();
 FILLCELL_X32 FILLER_308_2343 ();
 FILLCELL_X32 FILLER_308_2375 ();
 FILLCELL_X16 FILLER_308_2407 ();
 FILLCELL_X8 FILLER_308_2423 ();
 FILLCELL_X4 FILLER_308_2431 ();
 FILLCELL_X1 FILLER_308_2435 ();
 FILLCELL_X32 FILLER_309_1 ();
 FILLCELL_X32 FILLER_309_33 ();
 FILLCELL_X32 FILLER_309_65 ();
 FILLCELL_X32 FILLER_309_97 ();
 FILLCELL_X32 FILLER_309_129 ();
 FILLCELL_X32 FILLER_309_161 ();
 FILLCELL_X32 FILLER_309_193 ();
 FILLCELL_X32 FILLER_309_225 ();
 FILLCELL_X32 FILLER_309_257 ();
 FILLCELL_X32 FILLER_309_289 ();
 FILLCELL_X32 FILLER_309_321 ();
 FILLCELL_X32 FILLER_309_353 ();
 FILLCELL_X32 FILLER_309_385 ();
 FILLCELL_X32 FILLER_309_417 ();
 FILLCELL_X32 FILLER_309_449 ();
 FILLCELL_X32 FILLER_309_481 ();
 FILLCELL_X32 FILLER_309_513 ();
 FILLCELL_X32 FILLER_309_545 ();
 FILLCELL_X32 FILLER_309_577 ();
 FILLCELL_X32 FILLER_309_609 ();
 FILLCELL_X32 FILLER_309_641 ();
 FILLCELL_X32 FILLER_309_673 ();
 FILLCELL_X32 FILLER_309_705 ();
 FILLCELL_X32 FILLER_309_737 ();
 FILLCELL_X32 FILLER_309_769 ();
 FILLCELL_X32 FILLER_309_801 ();
 FILLCELL_X32 FILLER_309_833 ();
 FILLCELL_X32 FILLER_309_865 ();
 FILLCELL_X32 FILLER_309_897 ();
 FILLCELL_X4 FILLER_309_929 ();
 FILLCELL_X4 FILLER_309_947 ();
 FILLCELL_X2 FILLER_309_951 ();
 FILLCELL_X16 FILLER_309_961 ();
 FILLCELL_X2 FILLER_309_977 ();
 FILLCELL_X1 FILLER_309_979 ();
 FILLCELL_X16 FILLER_309_990 ();
 FILLCELL_X4 FILLER_309_1006 ();
 FILLCELL_X2 FILLER_309_1010 ();
 FILLCELL_X16 FILLER_309_1019 ();
 FILLCELL_X8 FILLER_309_1035 ();
 FILLCELL_X4 FILLER_309_1043 ();
 FILLCELL_X1 FILLER_309_1047 ();
 FILLCELL_X32 FILLER_309_1055 ();
 FILLCELL_X16 FILLER_309_1087 ();
 FILLCELL_X8 FILLER_309_1103 ();
 FILLCELL_X2 FILLER_309_1111 ();
 FILLCELL_X32 FILLER_309_1123 ();
 FILLCELL_X32 FILLER_309_1155 ();
 FILLCELL_X16 FILLER_309_1187 ();
 FILLCELL_X8 FILLER_309_1203 ();
 FILLCELL_X2 FILLER_309_1211 ();
 FILLCELL_X1 FILLER_309_1213 ();
 FILLCELL_X2 FILLER_309_1223 ();
 FILLCELL_X2 FILLER_309_1234 ();
 FILLCELL_X32 FILLER_309_1264 ();
 FILLCELL_X8 FILLER_309_1296 ();
 FILLCELL_X4 FILLER_309_1304 ();
 FILLCELL_X32 FILLER_309_1310 ();
 FILLCELL_X32 FILLER_309_1342 ();
 FILLCELL_X32 FILLER_309_1374 ();
 FILLCELL_X32 FILLER_309_1406 ();
 FILLCELL_X32 FILLER_309_1438 ();
 FILLCELL_X32 FILLER_309_1470 ();
 FILLCELL_X32 FILLER_309_1502 ();
 FILLCELL_X32 FILLER_309_1534 ();
 FILLCELL_X32 FILLER_309_1566 ();
 FILLCELL_X32 FILLER_309_1598 ();
 FILLCELL_X32 FILLER_309_1630 ();
 FILLCELL_X32 FILLER_309_1662 ();
 FILLCELL_X32 FILLER_309_1694 ();
 FILLCELL_X32 FILLER_309_1726 ();
 FILLCELL_X32 FILLER_309_1758 ();
 FILLCELL_X32 FILLER_309_1790 ();
 FILLCELL_X32 FILLER_309_1822 ();
 FILLCELL_X32 FILLER_309_1854 ();
 FILLCELL_X32 FILLER_309_1886 ();
 FILLCELL_X32 FILLER_309_1918 ();
 FILLCELL_X32 FILLER_309_1950 ();
 FILLCELL_X32 FILLER_309_1982 ();
 FILLCELL_X32 FILLER_309_2014 ();
 FILLCELL_X32 FILLER_309_2046 ();
 FILLCELL_X32 FILLER_309_2078 ();
 FILLCELL_X32 FILLER_309_2110 ();
 FILLCELL_X32 FILLER_309_2142 ();
 FILLCELL_X32 FILLER_309_2174 ();
 FILLCELL_X32 FILLER_309_2206 ();
 FILLCELL_X32 FILLER_309_2238 ();
 FILLCELL_X32 FILLER_309_2270 ();
 FILLCELL_X32 FILLER_309_2302 ();
 FILLCELL_X32 FILLER_309_2334 ();
 FILLCELL_X32 FILLER_309_2366 ();
 FILLCELL_X32 FILLER_309_2398 ();
 FILLCELL_X4 FILLER_309_2430 ();
 FILLCELL_X2 FILLER_309_2434 ();
 FILLCELL_X32 FILLER_310_1 ();
 FILLCELL_X32 FILLER_310_33 ();
 FILLCELL_X32 FILLER_310_65 ();
 FILLCELL_X32 FILLER_310_97 ();
 FILLCELL_X32 FILLER_310_129 ();
 FILLCELL_X32 FILLER_310_161 ();
 FILLCELL_X32 FILLER_310_193 ();
 FILLCELL_X32 FILLER_310_225 ();
 FILLCELL_X32 FILLER_310_257 ();
 FILLCELL_X32 FILLER_310_289 ();
 FILLCELL_X32 FILLER_310_321 ();
 FILLCELL_X32 FILLER_310_353 ();
 FILLCELL_X32 FILLER_310_385 ();
 FILLCELL_X32 FILLER_310_417 ();
 FILLCELL_X32 FILLER_310_449 ();
 FILLCELL_X32 FILLER_310_481 ();
 FILLCELL_X32 FILLER_310_513 ();
 FILLCELL_X32 FILLER_310_545 ();
 FILLCELL_X32 FILLER_310_577 ();
 FILLCELL_X16 FILLER_310_609 ();
 FILLCELL_X4 FILLER_310_625 ();
 FILLCELL_X2 FILLER_310_629 ();
 FILLCELL_X32 FILLER_310_632 ();
 FILLCELL_X32 FILLER_310_664 ();
 FILLCELL_X32 FILLER_310_696 ();
 FILLCELL_X32 FILLER_310_728 ();
 FILLCELL_X32 FILLER_310_760 ();
 FILLCELL_X32 FILLER_310_792 ();
 FILLCELL_X32 FILLER_310_824 ();
 FILLCELL_X32 FILLER_310_856 ();
 FILLCELL_X32 FILLER_310_888 ();
 FILLCELL_X4 FILLER_310_920 ();
 FILLCELL_X2 FILLER_310_924 ();
 FILLCELL_X1 FILLER_310_926 ();
 FILLCELL_X32 FILLER_310_943 ();
 FILLCELL_X16 FILLER_310_975 ();
 FILLCELL_X2 FILLER_310_991 ();
 FILLCELL_X1 FILLER_310_993 ();
 FILLCELL_X8 FILLER_310_1004 ();
 FILLCELL_X4 FILLER_310_1012 ();
 FILLCELL_X2 FILLER_310_1016 ();
 FILLCELL_X1 FILLER_310_1018 ();
 FILLCELL_X16 FILLER_310_1024 ();
 FILLCELL_X4 FILLER_310_1040 ();
 FILLCELL_X2 FILLER_310_1044 ();
 FILLCELL_X16 FILLER_310_1056 ();
 FILLCELL_X4 FILLER_310_1072 ();
 FILLCELL_X2 FILLER_310_1076 ();
 FILLCELL_X1 FILLER_310_1078 ();
 FILLCELL_X16 FILLER_310_1089 ();
 FILLCELL_X32 FILLER_310_1115 ();
 FILLCELL_X8 FILLER_310_1147 ();
 FILLCELL_X4 FILLER_310_1155 ();
 FILLCELL_X32 FILLER_310_1181 ();
 FILLCELL_X16 FILLER_310_1213 ();
 FILLCELL_X4 FILLER_310_1229 ();
 FILLCELL_X2 FILLER_310_1233 ();
 FILLCELL_X1 FILLER_310_1235 ();
 FILLCELL_X2 FILLER_310_1239 ();
 FILLCELL_X1 FILLER_310_1241 ();
 FILLCELL_X32 FILLER_310_1250 ();
 FILLCELL_X4 FILLER_310_1282 ();
 FILLCELL_X2 FILLER_310_1286 ();
 FILLCELL_X32 FILLER_310_1291 ();
 FILLCELL_X32 FILLER_310_1323 ();
 FILLCELL_X32 FILLER_310_1355 ();
 FILLCELL_X32 FILLER_310_1387 ();
 FILLCELL_X32 FILLER_310_1419 ();
 FILLCELL_X32 FILLER_310_1451 ();
 FILLCELL_X32 FILLER_310_1483 ();
 FILLCELL_X32 FILLER_310_1515 ();
 FILLCELL_X32 FILLER_310_1547 ();
 FILLCELL_X32 FILLER_310_1579 ();
 FILLCELL_X32 FILLER_310_1611 ();
 FILLCELL_X32 FILLER_310_1643 ();
 FILLCELL_X32 FILLER_310_1675 ();
 FILLCELL_X32 FILLER_310_1707 ();
 FILLCELL_X32 FILLER_310_1739 ();
 FILLCELL_X32 FILLER_310_1771 ();
 FILLCELL_X32 FILLER_310_1803 ();
 FILLCELL_X32 FILLER_310_1835 ();
 FILLCELL_X16 FILLER_310_1867 ();
 FILLCELL_X8 FILLER_310_1883 ();
 FILLCELL_X2 FILLER_310_1891 ();
 FILLCELL_X1 FILLER_310_1893 ();
 FILLCELL_X32 FILLER_310_1895 ();
 FILLCELL_X32 FILLER_310_1927 ();
 FILLCELL_X32 FILLER_310_1959 ();
 FILLCELL_X32 FILLER_310_1991 ();
 FILLCELL_X32 FILLER_310_2023 ();
 FILLCELL_X32 FILLER_310_2055 ();
 FILLCELL_X32 FILLER_310_2087 ();
 FILLCELL_X32 FILLER_310_2119 ();
 FILLCELL_X32 FILLER_310_2151 ();
 FILLCELL_X32 FILLER_310_2183 ();
 FILLCELL_X32 FILLER_310_2215 ();
 FILLCELL_X32 FILLER_310_2247 ();
 FILLCELL_X32 FILLER_310_2279 ();
 FILLCELL_X32 FILLER_310_2311 ();
 FILLCELL_X32 FILLER_310_2343 ();
 FILLCELL_X32 FILLER_310_2375 ();
 FILLCELL_X16 FILLER_310_2407 ();
 FILLCELL_X8 FILLER_310_2423 ();
 FILLCELL_X4 FILLER_310_2431 ();
 FILLCELL_X1 FILLER_310_2435 ();
 FILLCELL_X32 FILLER_311_1 ();
 FILLCELL_X32 FILLER_311_33 ();
 FILLCELL_X32 FILLER_311_65 ();
 FILLCELL_X32 FILLER_311_97 ();
 FILLCELL_X32 FILLER_311_129 ();
 FILLCELL_X32 FILLER_311_161 ();
 FILLCELL_X32 FILLER_311_193 ();
 FILLCELL_X32 FILLER_311_225 ();
 FILLCELL_X32 FILLER_311_257 ();
 FILLCELL_X32 FILLER_311_289 ();
 FILLCELL_X32 FILLER_311_321 ();
 FILLCELL_X32 FILLER_311_353 ();
 FILLCELL_X32 FILLER_311_385 ();
 FILLCELL_X32 FILLER_311_417 ();
 FILLCELL_X32 FILLER_311_449 ();
 FILLCELL_X32 FILLER_311_481 ();
 FILLCELL_X32 FILLER_311_513 ();
 FILLCELL_X32 FILLER_311_545 ();
 FILLCELL_X32 FILLER_311_577 ();
 FILLCELL_X32 FILLER_311_609 ();
 FILLCELL_X32 FILLER_311_641 ();
 FILLCELL_X32 FILLER_311_673 ();
 FILLCELL_X32 FILLER_311_705 ();
 FILLCELL_X32 FILLER_311_737 ();
 FILLCELL_X32 FILLER_311_769 ();
 FILLCELL_X32 FILLER_311_801 ();
 FILLCELL_X32 FILLER_311_833 ();
 FILLCELL_X32 FILLER_311_865 ();
 FILLCELL_X32 FILLER_311_897 ();
 FILLCELL_X32 FILLER_311_929 ();
 FILLCELL_X2 FILLER_311_961 ();
 FILLCELL_X1 FILLER_311_963 ();
 FILLCELL_X16 FILLER_311_966 ();
 FILLCELL_X8 FILLER_311_984 ();
 FILLCELL_X4 FILLER_311_992 ();
 FILLCELL_X1 FILLER_311_996 ();
 FILLCELL_X8 FILLER_311_999 ();
 FILLCELL_X4 FILLER_311_1007 ();
 FILLCELL_X32 FILLER_311_1021 ();
 FILLCELL_X32 FILLER_311_1053 ();
 FILLCELL_X16 FILLER_311_1085 ();
 FILLCELL_X2 FILLER_311_1101 ();
 FILLCELL_X16 FILLER_311_1105 ();
 FILLCELL_X4 FILLER_311_1121 ();
 FILLCELL_X1 FILLER_311_1125 ();
 FILLCELL_X32 FILLER_311_1136 ();
 FILLCELL_X32 FILLER_311_1168 ();
 FILLCELL_X32 FILLER_311_1200 ();
 FILLCELL_X16 FILLER_311_1232 ();
 FILLCELL_X8 FILLER_311_1248 ();
 FILLCELL_X4 FILLER_311_1256 ();
 FILLCELL_X2 FILLER_311_1260 ();
 FILLCELL_X1 FILLER_311_1262 ();
 FILLCELL_X8 FILLER_311_1264 ();
 FILLCELL_X4 FILLER_311_1272 ();
 FILLCELL_X2 FILLER_311_1276 ();
 FILLCELL_X8 FILLER_311_1302 ();
 FILLCELL_X2 FILLER_311_1310 ();
 FILLCELL_X8 FILLER_311_1316 ();
 FILLCELL_X2 FILLER_311_1324 ();
 FILLCELL_X32 FILLER_311_1329 ();
 FILLCELL_X32 FILLER_311_1361 ();
 FILLCELL_X32 FILLER_311_1393 ();
 FILLCELL_X32 FILLER_311_1425 ();
 FILLCELL_X32 FILLER_311_1457 ();
 FILLCELL_X32 FILLER_311_1489 ();
 FILLCELL_X32 FILLER_311_1521 ();
 FILLCELL_X32 FILLER_311_1553 ();
 FILLCELL_X32 FILLER_311_1585 ();
 FILLCELL_X32 FILLER_311_1617 ();
 FILLCELL_X32 FILLER_311_1649 ();
 FILLCELL_X32 FILLER_311_1681 ();
 FILLCELL_X32 FILLER_311_1713 ();
 FILLCELL_X32 FILLER_311_1745 ();
 FILLCELL_X32 FILLER_311_1777 ();
 FILLCELL_X32 FILLER_311_1809 ();
 FILLCELL_X32 FILLER_311_1841 ();
 FILLCELL_X32 FILLER_311_1873 ();
 FILLCELL_X32 FILLER_311_1905 ();
 FILLCELL_X32 FILLER_311_1937 ();
 FILLCELL_X32 FILLER_311_1969 ();
 FILLCELL_X32 FILLER_311_2001 ();
 FILLCELL_X32 FILLER_311_2033 ();
 FILLCELL_X32 FILLER_311_2065 ();
 FILLCELL_X32 FILLER_311_2097 ();
 FILLCELL_X32 FILLER_311_2129 ();
 FILLCELL_X32 FILLER_311_2161 ();
 FILLCELL_X32 FILLER_311_2193 ();
 FILLCELL_X32 FILLER_311_2225 ();
 FILLCELL_X32 FILLER_311_2257 ();
 FILLCELL_X32 FILLER_311_2289 ();
 FILLCELL_X32 FILLER_311_2321 ();
 FILLCELL_X32 FILLER_311_2353 ();
 FILLCELL_X32 FILLER_311_2385 ();
 FILLCELL_X16 FILLER_311_2417 ();
 FILLCELL_X2 FILLER_311_2433 ();
 FILLCELL_X1 FILLER_311_2435 ();
 FILLCELL_X32 FILLER_312_1 ();
 FILLCELL_X32 FILLER_312_33 ();
 FILLCELL_X32 FILLER_312_65 ();
 FILLCELL_X32 FILLER_312_97 ();
 FILLCELL_X32 FILLER_312_129 ();
 FILLCELL_X32 FILLER_312_161 ();
 FILLCELL_X32 FILLER_312_193 ();
 FILLCELL_X32 FILLER_312_225 ();
 FILLCELL_X32 FILLER_312_257 ();
 FILLCELL_X32 FILLER_312_289 ();
 FILLCELL_X32 FILLER_312_321 ();
 FILLCELL_X32 FILLER_312_353 ();
 FILLCELL_X32 FILLER_312_385 ();
 FILLCELL_X32 FILLER_312_417 ();
 FILLCELL_X32 FILLER_312_449 ();
 FILLCELL_X32 FILLER_312_481 ();
 FILLCELL_X32 FILLER_312_513 ();
 FILLCELL_X32 FILLER_312_545 ();
 FILLCELL_X32 FILLER_312_577 ();
 FILLCELL_X16 FILLER_312_609 ();
 FILLCELL_X4 FILLER_312_625 ();
 FILLCELL_X2 FILLER_312_629 ();
 FILLCELL_X32 FILLER_312_632 ();
 FILLCELL_X32 FILLER_312_664 ();
 FILLCELL_X32 FILLER_312_696 ();
 FILLCELL_X32 FILLER_312_728 ();
 FILLCELL_X32 FILLER_312_760 ();
 FILLCELL_X32 FILLER_312_792 ();
 FILLCELL_X32 FILLER_312_824 ();
 FILLCELL_X32 FILLER_312_856 ();
 FILLCELL_X32 FILLER_312_888 ();
 FILLCELL_X8 FILLER_312_920 ();
 FILLCELL_X4 FILLER_312_928 ();
 FILLCELL_X2 FILLER_312_932 ();
 FILLCELL_X16 FILLER_312_938 ();
 FILLCELL_X4 FILLER_312_954 ();
 FILLCELL_X2 FILLER_312_958 ();
 FILLCELL_X1 FILLER_312_960 ();
 FILLCELL_X2 FILLER_312_977 ();
 FILLCELL_X1 FILLER_312_979 ();
 FILLCELL_X1 FILLER_312_982 ();
 FILLCELL_X16 FILLER_312_999 ();
 FILLCELL_X1 FILLER_312_1015 ();
 FILLCELL_X8 FILLER_312_1018 ();
 FILLCELL_X1 FILLER_312_1026 ();
 FILLCELL_X32 FILLER_312_1029 ();
 FILLCELL_X1 FILLER_312_1061 ();
 FILLCELL_X16 FILLER_312_1081 ();
 FILLCELL_X8 FILLER_312_1097 ();
 FILLCELL_X2 FILLER_312_1105 ();
 FILLCELL_X1 FILLER_312_1125 ();
 FILLCELL_X8 FILLER_312_1128 ();
 FILLCELL_X2 FILLER_312_1136 ();
 FILLCELL_X1 FILLER_312_1138 ();
 FILLCELL_X16 FILLER_312_1149 ();
 FILLCELL_X8 FILLER_312_1167 ();
 FILLCELL_X2 FILLER_312_1175 ();
 FILLCELL_X1 FILLER_312_1177 ();
 FILLCELL_X8 FILLER_312_1182 ();
 FILLCELL_X1 FILLER_312_1190 ();
 FILLCELL_X2 FILLER_312_1201 ();
 FILLCELL_X32 FILLER_312_1217 ();
 FILLCELL_X16 FILLER_312_1249 ();
 FILLCELL_X8 FILLER_312_1265 ();
 FILLCELL_X2 FILLER_312_1273 ();
 FILLCELL_X1 FILLER_312_1275 ();
 FILLCELL_X4 FILLER_312_1290 ();
 FILLCELL_X2 FILLER_312_1294 ();
 FILLCELL_X2 FILLER_312_1308 ();
 FILLCELL_X1 FILLER_312_1316 ();
 FILLCELL_X32 FILLER_312_1350 ();
 FILLCELL_X32 FILLER_312_1382 ();
 FILLCELL_X32 FILLER_312_1414 ();
 FILLCELL_X32 FILLER_312_1446 ();
 FILLCELL_X32 FILLER_312_1478 ();
 FILLCELL_X32 FILLER_312_1510 ();
 FILLCELL_X32 FILLER_312_1542 ();
 FILLCELL_X32 FILLER_312_1574 ();
 FILLCELL_X32 FILLER_312_1606 ();
 FILLCELL_X32 FILLER_312_1638 ();
 FILLCELL_X32 FILLER_312_1670 ();
 FILLCELL_X32 FILLER_312_1702 ();
 FILLCELL_X32 FILLER_312_1734 ();
 FILLCELL_X32 FILLER_312_1766 ();
 FILLCELL_X32 FILLER_312_1798 ();
 FILLCELL_X32 FILLER_312_1830 ();
 FILLCELL_X32 FILLER_312_1862 ();
 FILLCELL_X32 FILLER_312_1895 ();
 FILLCELL_X32 FILLER_312_1927 ();
 FILLCELL_X32 FILLER_312_1959 ();
 FILLCELL_X32 FILLER_312_1991 ();
 FILLCELL_X32 FILLER_312_2023 ();
 FILLCELL_X32 FILLER_312_2055 ();
 FILLCELL_X32 FILLER_312_2087 ();
 FILLCELL_X32 FILLER_312_2119 ();
 FILLCELL_X32 FILLER_312_2151 ();
 FILLCELL_X32 FILLER_312_2183 ();
 FILLCELL_X32 FILLER_312_2215 ();
 FILLCELL_X32 FILLER_312_2247 ();
 FILLCELL_X32 FILLER_312_2279 ();
 FILLCELL_X32 FILLER_312_2311 ();
 FILLCELL_X32 FILLER_312_2343 ();
 FILLCELL_X32 FILLER_312_2375 ();
 FILLCELL_X16 FILLER_312_2407 ();
 FILLCELL_X8 FILLER_312_2423 ();
 FILLCELL_X4 FILLER_312_2431 ();
 FILLCELL_X1 FILLER_312_2435 ();
 FILLCELL_X32 FILLER_313_1 ();
 FILLCELL_X32 FILLER_313_33 ();
 FILLCELL_X32 FILLER_313_65 ();
 FILLCELL_X32 FILLER_313_97 ();
 FILLCELL_X32 FILLER_313_129 ();
 FILLCELL_X32 FILLER_313_161 ();
 FILLCELL_X32 FILLER_313_193 ();
 FILLCELL_X32 FILLER_313_225 ();
 FILLCELL_X32 FILLER_313_257 ();
 FILLCELL_X32 FILLER_313_289 ();
 FILLCELL_X32 FILLER_313_321 ();
 FILLCELL_X32 FILLER_313_353 ();
 FILLCELL_X32 FILLER_313_385 ();
 FILLCELL_X32 FILLER_313_417 ();
 FILLCELL_X32 FILLER_313_449 ();
 FILLCELL_X32 FILLER_313_481 ();
 FILLCELL_X32 FILLER_313_513 ();
 FILLCELL_X32 FILLER_313_545 ();
 FILLCELL_X32 FILLER_313_577 ();
 FILLCELL_X32 FILLER_313_609 ();
 FILLCELL_X32 FILLER_313_641 ();
 FILLCELL_X32 FILLER_313_673 ();
 FILLCELL_X32 FILLER_313_705 ();
 FILLCELL_X32 FILLER_313_737 ();
 FILLCELL_X32 FILLER_313_769 ();
 FILLCELL_X32 FILLER_313_801 ();
 FILLCELL_X32 FILLER_313_833 ();
 FILLCELL_X32 FILLER_313_865 ();
 FILLCELL_X32 FILLER_313_897 ();
 FILLCELL_X4 FILLER_313_929 ();
 FILLCELL_X2 FILLER_313_933 ();
 FILLCELL_X1 FILLER_313_935 ();
 FILLCELL_X16 FILLER_313_946 ();
 FILLCELL_X4 FILLER_313_962 ();
 FILLCELL_X2 FILLER_313_966 ();
 FILLCELL_X8 FILLER_313_970 ();
 FILLCELL_X2 FILLER_313_978 ();
 FILLCELL_X16 FILLER_313_982 ();
 FILLCELL_X32 FILLER_313_1000 ();
 FILLCELL_X8 FILLER_313_1032 ();
 FILLCELL_X4 FILLER_313_1040 ();
 FILLCELL_X2 FILLER_313_1044 ();
 FILLCELL_X16 FILLER_313_1049 ();
 FILLCELL_X16 FILLER_313_1095 ();
 FILLCELL_X8 FILLER_313_1111 ();
 FILLCELL_X2 FILLER_313_1119 ();
 FILLCELL_X8 FILLER_313_1123 ();
 FILLCELL_X4 FILLER_313_1131 ();
 FILLCELL_X2 FILLER_313_1135 ();
 FILLCELL_X1 FILLER_313_1137 ();
 FILLCELL_X4 FILLER_313_1140 ();
 FILLCELL_X1 FILLER_313_1144 ();
 FILLCELL_X2 FILLER_313_1163 ();
 FILLCELL_X1 FILLER_313_1165 ();
 FILLCELL_X8 FILLER_313_1186 ();
 FILLCELL_X4 FILLER_313_1194 ();
 FILLCELL_X1 FILLER_313_1198 ();
 FILLCELL_X2 FILLER_313_1209 ();
 FILLCELL_X32 FILLER_313_1231 ();
 FILLCELL_X4 FILLER_313_1264 ();
 FILLCELL_X2 FILLER_313_1268 ();
 FILLCELL_X1 FILLER_313_1281 ();
 FILLCELL_X1 FILLER_313_1285 ();
 FILLCELL_X4 FILLER_313_1299 ();
 FILLCELL_X32 FILLER_313_1346 ();
 FILLCELL_X32 FILLER_313_1378 ();
 FILLCELL_X32 FILLER_313_1410 ();
 FILLCELL_X32 FILLER_313_1442 ();
 FILLCELL_X32 FILLER_313_1474 ();
 FILLCELL_X32 FILLER_313_1506 ();
 FILLCELL_X32 FILLER_313_1538 ();
 FILLCELL_X32 FILLER_313_1570 ();
 FILLCELL_X32 FILLER_313_1602 ();
 FILLCELL_X32 FILLER_313_1634 ();
 FILLCELL_X32 FILLER_313_1666 ();
 FILLCELL_X32 FILLER_313_1698 ();
 FILLCELL_X32 FILLER_313_1730 ();
 FILLCELL_X32 FILLER_313_1762 ();
 FILLCELL_X32 FILLER_313_1794 ();
 FILLCELL_X32 FILLER_313_1826 ();
 FILLCELL_X32 FILLER_313_1858 ();
 FILLCELL_X32 FILLER_313_1890 ();
 FILLCELL_X32 FILLER_313_1922 ();
 FILLCELL_X32 FILLER_313_1954 ();
 FILLCELL_X32 FILLER_313_1986 ();
 FILLCELL_X32 FILLER_313_2018 ();
 FILLCELL_X32 FILLER_313_2050 ();
 FILLCELL_X32 FILLER_313_2082 ();
 FILLCELL_X32 FILLER_313_2114 ();
 FILLCELL_X32 FILLER_313_2146 ();
 FILLCELL_X32 FILLER_313_2178 ();
 FILLCELL_X32 FILLER_313_2210 ();
 FILLCELL_X32 FILLER_313_2242 ();
 FILLCELL_X32 FILLER_313_2274 ();
 FILLCELL_X32 FILLER_313_2306 ();
 FILLCELL_X32 FILLER_313_2338 ();
 FILLCELL_X32 FILLER_313_2370 ();
 FILLCELL_X32 FILLER_313_2402 ();
 FILLCELL_X2 FILLER_313_2434 ();
 FILLCELL_X32 FILLER_314_1 ();
 FILLCELL_X32 FILLER_314_33 ();
 FILLCELL_X32 FILLER_314_65 ();
 FILLCELL_X32 FILLER_314_97 ();
 FILLCELL_X32 FILLER_314_129 ();
 FILLCELL_X32 FILLER_314_161 ();
 FILLCELL_X32 FILLER_314_193 ();
 FILLCELL_X32 FILLER_314_225 ();
 FILLCELL_X32 FILLER_314_257 ();
 FILLCELL_X32 FILLER_314_289 ();
 FILLCELL_X32 FILLER_314_321 ();
 FILLCELL_X32 FILLER_314_353 ();
 FILLCELL_X32 FILLER_314_385 ();
 FILLCELL_X32 FILLER_314_417 ();
 FILLCELL_X32 FILLER_314_449 ();
 FILLCELL_X32 FILLER_314_481 ();
 FILLCELL_X32 FILLER_314_513 ();
 FILLCELL_X32 FILLER_314_545 ();
 FILLCELL_X32 FILLER_314_577 ();
 FILLCELL_X16 FILLER_314_609 ();
 FILLCELL_X4 FILLER_314_625 ();
 FILLCELL_X2 FILLER_314_629 ();
 FILLCELL_X32 FILLER_314_632 ();
 FILLCELL_X32 FILLER_314_664 ();
 FILLCELL_X32 FILLER_314_696 ();
 FILLCELL_X32 FILLER_314_728 ();
 FILLCELL_X32 FILLER_314_760 ();
 FILLCELL_X32 FILLER_314_792 ();
 FILLCELL_X32 FILLER_314_824 ();
 FILLCELL_X32 FILLER_314_856 ();
 FILLCELL_X32 FILLER_314_888 ();
 FILLCELL_X8 FILLER_314_920 ();
 FILLCELL_X4 FILLER_314_928 ();
 FILLCELL_X2 FILLER_314_932 ();
 FILLCELL_X2 FILLER_314_958 ();
 FILLCELL_X1 FILLER_314_960 ();
 FILLCELL_X2 FILLER_314_977 ();
 FILLCELL_X1 FILLER_314_979 ();
 FILLCELL_X8 FILLER_314_982 ();
 FILLCELL_X2 FILLER_314_990 ();
 FILLCELL_X1 FILLER_314_992 ();
 FILLCELL_X8 FILLER_314_995 ();
 FILLCELL_X4 FILLER_314_1003 ();
 FILLCELL_X4 FILLER_314_1025 ();
 FILLCELL_X2 FILLER_314_1047 ();
 FILLCELL_X1 FILLER_314_1049 ();
 FILLCELL_X16 FILLER_314_1052 ();
 FILLCELL_X1 FILLER_314_1068 ();
 FILLCELL_X32 FILLER_314_1072 ();
 FILLCELL_X32 FILLER_314_1104 ();
 FILLCELL_X16 FILLER_314_1136 ();
 FILLCELL_X8 FILLER_314_1152 ();
 FILLCELL_X4 FILLER_314_1160 ();
 FILLCELL_X1 FILLER_314_1167 ();
 FILLCELL_X16 FILLER_314_1170 ();
 FILLCELL_X8 FILLER_314_1186 ();
 FILLCELL_X4 FILLER_314_1194 ();
 FILLCELL_X1 FILLER_314_1198 ();
 FILLCELL_X8 FILLER_314_1228 ();
 FILLCELL_X1 FILLER_314_1236 ();
 FILLCELL_X32 FILLER_314_1247 ();
 FILLCELL_X4 FILLER_314_1279 ();
 FILLCELL_X1 FILLER_314_1294 ();
 FILLCELL_X4 FILLER_314_1318 ();
 FILLCELL_X2 FILLER_314_1322 ();
 FILLCELL_X1 FILLER_314_1324 ();
 FILLCELL_X32 FILLER_314_1327 ();
 FILLCELL_X32 FILLER_314_1359 ();
 FILLCELL_X32 FILLER_314_1391 ();
 FILLCELL_X32 FILLER_314_1423 ();
 FILLCELL_X32 FILLER_314_1455 ();
 FILLCELL_X32 FILLER_314_1487 ();
 FILLCELL_X32 FILLER_314_1519 ();
 FILLCELL_X32 FILLER_314_1551 ();
 FILLCELL_X32 FILLER_314_1583 ();
 FILLCELL_X32 FILLER_314_1615 ();
 FILLCELL_X32 FILLER_314_1647 ();
 FILLCELL_X32 FILLER_314_1679 ();
 FILLCELL_X32 FILLER_314_1711 ();
 FILLCELL_X32 FILLER_314_1743 ();
 FILLCELL_X32 FILLER_314_1775 ();
 FILLCELL_X32 FILLER_314_1807 ();
 FILLCELL_X32 FILLER_314_1839 ();
 FILLCELL_X16 FILLER_314_1871 ();
 FILLCELL_X4 FILLER_314_1887 ();
 FILLCELL_X2 FILLER_314_1891 ();
 FILLCELL_X1 FILLER_314_1893 ();
 FILLCELL_X32 FILLER_314_1895 ();
 FILLCELL_X32 FILLER_314_1927 ();
 FILLCELL_X32 FILLER_314_1959 ();
 FILLCELL_X32 FILLER_314_1991 ();
 FILLCELL_X32 FILLER_314_2023 ();
 FILLCELL_X32 FILLER_314_2055 ();
 FILLCELL_X32 FILLER_314_2087 ();
 FILLCELL_X32 FILLER_314_2119 ();
 FILLCELL_X32 FILLER_314_2151 ();
 FILLCELL_X32 FILLER_314_2183 ();
 FILLCELL_X32 FILLER_314_2215 ();
 FILLCELL_X32 FILLER_314_2247 ();
 FILLCELL_X32 FILLER_314_2279 ();
 FILLCELL_X32 FILLER_314_2311 ();
 FILLCELL_X32 FILLER_314_2343 ();
 FILLCELL_X32 FILLER_314_2375 ();
 FILLCELL_X16 FILLER_314_2407 ();
 FILLCELL_X8 FILLER_314_2423 ();
 FILLCELL_X4 FILLER_314_2431 ();
 FILLCELL_X1 FILLER_314_2435 ();
 FILLCELL_X32 FILLER_315_1 ();
 FILLCELL_X32 FILLER_315_33 ();
 FILLCELL_X32 FILLER_315_65 ();
 FILLCELL_X32 FILLER_315_97 ();
 FILLCELL_X32 FILLER_315_129 ();
 FILLCELL_X32 FILLER_315_161 ();
 FILLCELL_X32 FILLER_315_193 ();
 FILLCELL_X32 FILLER_315_225 ();
 FILLCELL_X32 FILLER_315_257 ();
 FILLCELL_X32 FILLER_315_289 ();
 FILLCELL_X32 FILLER_315_321 ();
 FILLCELL_X32 FILLER_315_353 ();
 FILLCELL_X32 FILLER_315_385 ();
 FILLCELL_X32 FILLER_315_417 ();
 FILLCELL_X32 FILLER_315_449 ();
 FILLCELL_X32 FILLER_315_481 ();
 FILLCELL_X32 FILLER_315_513 ();
 FILLCELL_X32 FILLER_315_545 ();
 FILLCELL_X32 FILLER_315_577 ();
 FILLCELL_X32 FILLER_315_609 ();
 FILLCELL_X32 FILLER_315_641 ();
 FILLCELL_X32 FILLER_315_673 ();
 FILLCELL_X32 FILLER_315_705 ();
 FILLCELL_X32 FILLER_315_737 ();
 FILLCELL_X32 FILLER_315_769 ();
 FILLCELL_X32 FILLER_315_801 ();
 FILLCELL_X32 FILLER_315_833 ();
 FILLCELL_X32 FILLER_315_865 ();
 FILLCELL_X32 FILLER_315_897 ();
 FILLCELL_X32 FILLER_315_929 ();
 FILLCELL_X4 FILLER_315_961 ();
 FILLCELL_X2 FILLER_315_965 ();
 FILLCELL_X1 FILLER_315_967 ();
 FILLCELL_X2 FILLER_315_984 ();
 FILLCELL_X2 FILLER_315_990 ();
 FILLCELL_X1 FILLER_315_992 ();
 FILLCELL_X8 FILLER_315_1012 ();
 FILLCELL_X4 FILLER_315_1020 ();
 FILLCELL_X16 FILLER_315_1026 ();
 FILLCELL_X8 FILLER_315_1042 ();
 FILLCELL_X4 FILLER_315_1050 ();
 FILLCELL_X16 FILLER_315_1058 ();
 FILLCELL_X8 FILLER_315_1074 ();
 FILLCELL_X2 FILLER_315_1082 ();
 FILLCELL_X1 FILLER_315_1084 ();
 FILLCELL_X8 FILLER_315_1089 ();
 FILLCELL_X4 FILLER_315_1097 ();
 FILLCELL_X2 FILLER_315_1101 ();
 FILLCELL_X1 FILLER_315_1103 ();
 FILLCELL_X16 FILLER_315_1136 ();
 FILLCELL_X1 FILLER_315_1155 ();
 FILLCELL_X1 FILLER_315_1164 ();
 FILLCELL_X32 FILLER_315_1179 ();
 FILLCELL_X16 FILLER_315_1211 ();
 FILLCELL_X8 FILLER_315_1227 ();
 FILLCELL_X4 FILLER_315_1235 ();
 FILLCELL_X2 FILLER_315_1239 ();
 FILLCELL_X1 FILLER_315_1243 ();
 FILLCELL_X4 FILLER_315_1246 ();
 FILLCELL_X1 FILLER_315_1250 ();
 FILLCELL_X2 FILLER_315_1260 ();
 FILLCELL_X1 FILLER_315_1262 ();
 FILLCELL_X2 FILLER_315_1264 ();
 FILLCELL_X16 FILLER_315_1280 ();
 FILLCELL_X2 FILLER_315_1296 ();
 FILLCELL_X4 FILLER_315_1319 ();
 FILLCELL_X32 FILLER_315_1328 ();
 FILLCELL_X32 FILLER_315_1360 ();
 FILLCELL_X32 FILLER_315_1392 ();
 FILLCELL_X32 FILLER_315_1424 ();
 FILLCELL_X32 FILLER_315_1456 ();
 FILLCELL_X32 FILLER_315_1488 ();
 FILLCELL_X32 FILLER_315_1520 ();
 FILLCELL_X32 FILLER_315_1552 ();
 FILLCELL_X32 FILLER_315_1584 ();
 FILLCELL_X32 FILLER_315_1616 ();
 FILLCELL_X32 FILLER_315_1648 ();
 FILLCELL_X32 FILLER_315_1680 ();
 FILLCELL_X32 FILLER_315_1712 ();
 FILLCELL_X32 FILLER_315_1744 ();
 FILLCELL_X32 FILLER_315_1776 ();
 FILLCELL_X32 FILLER_315_1808 ();
 FILLCELL_X32 FILLER_315_1840 ();
 FILLCELL_X32 FILLER_315_1872 ();
 FILLCELL_X32 FILLER_315_1904 ();
 FILLCELL_X32 FILLER_315_1936 ();
 FILLCELL_X32 FILLER_315_1968 ();
 FILLCELL_X32 FILLER_315_2000 ();
 FILLCELL_X32 FILLER_315_2032 ();
 FILLCELL_X32 FILLER_315_2064 ();
 FILLCELL_X32 FILLER_315_2096 ();
 FILLCELL_X32 FILLER_315_2128 ();
 FILLCELL_X32 FILLER_315_2160 ();
 FILLCELL_X32 FILLER_315_2192 ();
 FILLCELL_X32 FILLER_315_2224 ();
 FILLCELL_X32 FILLER_315_2256 ();
 FILLCELL_X32 FILLER_315_2288 ();
 FILLCELL_X32 FILLER_315_2320 ();
 FILLCELL_X32 FILLER_315_2352 ();
 FILLCELL_X32 FILLER_315_2384 ();
 FILLCELL_X16 FILLER_315_2416 ();
 FILLCELL_X4 FILLER_315_2432 ();
 FILLCELL_X32 FILLER_316_1 ();
 FILLCELL_X32 FILLER_316_33 ();
 FILLCELL_X32 FILLER_316_65 ();
 FILLCELL_X32 FILLER_316_97 ();
 FILLCELL_X32 FILLER_316_129 ();
 FILLCELL_X32 FILLER_316_161 ();
 FILLCELL_X32 FILLER_316_193 ();
 FILLCELL_X32 FILLER_316_225 ();
 FILLCELL_X32 FILLER_316_257 ();
 FILLCELL_X32 FILLER_316_289 ();
 FILLCELL_X32 FILLER_316_321 ();
 FILLCELL_X32 FILLER_316_353 ();
 FILLCELL_X32 FILLER_316_385 ();
 FILLCELL_X32 FILLER_316_417 ();
 FILLCELL_X32 FILLER_316_449 ();
 FILLCELL_X32 FILLER_316_481 ();
 FILLCELL_X32 FILLER_316_513 ();
 FILLCELL_X32 FILLER_316_545 ();
 FILLCELL_X32 FILLER_316_577 ();
 FILLCELL_X16 FILLER_316_609 ();
 FILLCELL_X4 FILLER_316_625 ();
 FILLCELL_X2 FILLER_316_629 ();
 FILLCELL_X32 FILLER_316_632 ();
 FILLCELL_X32 FILLER_316_664 ();
 FILLCELL_X32 FILLER_316_696 ();
 FILLCELL_X32 FILLER_316_728 ();
 FILLCELL_X32 FILLER_316_760 ();
 FILLCELL_X32 FILLER_316_792 ();
 FILLCELL_X32 FILLER_316_824 ();
 FILLCELL_X32 FILLER_316_856 ();
 FILLCELL_X32 FILLER_316_888 ();
 FILLCELL_X16 FILLER_316_920 ();
 FILLCELL_X1 FILLER_316_936 ();
 FILLCELL_X32 FILLER_316_941 ();
 FILLCELL_X2 FILLER_316_973 ();
 FILLCELL_X1 FILLER_316_975 ();
 FILLCELL_X8 FILLER_316_980 ();
 FILLCELL_X2 FILLER_316_988 ();
 FILLCELL_X1 FILLER_316_990 ();
 FILLCELL_X16 FILLER_316_1007 ();
 FILLCELL_X4 FILLER_316_1023 ();
 FILLCELL_X1 FILLER_316_1030 ();
 FILLCELL_X8 FILLER_316_1035 ();
 FILLCELL_X4 FILLER_316_1043 ();
 FILLCELL_X1 FILLER_316_1047 ();
 FILLCELL_X8 FILLER_316_1068 ();
 FILLCELL_X2 FILLER_316_1076 ();
 FILLCELL_X32 FILLER_316_1082 ();
 FILLCELL_X32 FILLER_316_1114 ();
 FILLCELL_X8 FILLER_316_1146 ();
 FILLCELL_X2 FILLER_316_1154 ();
 FILLCELL_X32 FILLER_316_1170 ();
 FILLCELL_X16 FILLER_316_1202 ();
 FILLCELL_X8 FILLER_316_1218 ();
 FILLCELL_X4 FILLER_316_1226 ();
 FILLCELL_X32 FILLER_316_1269 ();
 FILLCELL_X2 FILLER_316_1305 ();
 FILLCELL_X32 FILLER_316_1310 ();
 FILLCELL_X32 FILLER_316_1342 ();
 FILLCELL_X32 FILLER_316_1374 ();
 FILLCELL_X32 FILLER_316_1406 ();
 FILLCELL_X32 FILLER_316_1438 ();
 FILLCELL_X32 FILLER_316_1470 ();
 FILLCELL_X32 FILLER_316_1502 ();
 FILLCELL_X32 FILLER_316_1534 ();
 FILLCELL_X32 FILLER_316_1566 ();
 FILLCELL_X32 FILLER_316_1598 ();
 FILLCELL_X32 FILLER_316_1630 ();
 FILLCELL_X32 FILLER_316_1662 ();
 FILLCELL_X32 FILLER_316_1694 ();
 FILLCELL_X32 FILLER_316_1726 ();
 FILLCELL_X32 FILLER_316_1758 ();
 FILLCELL_X32 FILLER_316_1790 ();
 FILLCELL_X32 FILLER_316_1822 ();
 FILLCELL_X32 FILLER_316_1854 ();
 FILLCELL_X8 FILLER_316_1886 ();
 FILLCELL_X32 FILLER_316_1895 ();
 FILLCELL_X32 FILLER_316_1927 ();
 FILLCELL_X32 FILLER_316_1959 ();
 FILLCELL_X32 FILLER_316_1991 ();
 FILLCELL_X32 FILLER_316_2023 ();
 FILLCELL_X32 FILLER_316_2055 ();
 FILLCELL_X32 FILLER_316_2087 ();
 FILLCELL_X32 FILLER_316_2119 ();
 FILLCELL_X32 FILLER_316_2151 ();
 FILLCELL_X32 FILLER_316_2183 ();
 FILLCELL_X32 FILLER_316_2215 ();
 FILLCELL_X32 FILLER_316_2247 ();
 FILLCELL_X32 FILLER_316_2279 ();
 FILLCELL_X32 FILLER_316_2311 ();
 FILLCELL_X32 FILLER_316_2343 ();
 FILLCELL_X32 FILLER_316_2375 ();
 FILLCELL_X16 FILLER_316_2407 ();
 FILLCELL_X8 FILLER_316_2423 ();
 FILLCELL_X4 FILLER_316_2431 ();
 FILLCELL_X1 FILLER_316_2435 ();
 FILLCELL_X32 FILLER_317_1 ();
 FILLCELL_X32 FILLER_317_33 ();
 FILLCELL_X32 FILLER_317_65 ();
 FILLCELL_X32 FILLER_317_97 ();
 FILLCELL_X32 FILLER_317_129 ();
 FILLCELL_X32 FILLER_317_161 ();
 FILLCELL_X32 FILLER_317_193 ();
 FILLCELL_X32 FILLER_317_225 ();
 FILLCELL_X32 FILLER_317_257 ();
 FILLCELL_X32 FILLER_317_289 ();
 FILLCELL_X32 FILLER_317_321 ();
 FILLCELL_X32 FILLER_317_353 ();
 FILLCELL_X32 FILLER_317_385 ();
 FILLCELL_X32 FILLER_317_417 ();
 FILLCELL_X32 FILLER_317_449 ();
 FILLCELL_X32 FILLER_317_481 ();
 FILLCELL_X32 FILLER_317_513 ();
 FILLCELL_X32 FILLER_317_545 ();
 FILLCELL_X32 FILLER_317_577 ();
 FILLCELL_X32 FILLER_317_609 ();
 FILLCELL_X32 FILLER_317_641 ();
 FILLCELL_X32 FILLER_317_673 ();
 FILLCELL_X32 FILLER_317_705 ();
 FILLCELL_X32 FILLER_317_737 ();
 FILLCELL_X32 FILLER_317_769 ();
 FILLCELL_X32 FILLER_317_801 ();
 FILLCELL_X32 FILLER_317_833 ();
 FILLCELL_X32 FILLER_317_865 ();
 FILLCELL_X32 FILLER_317_897 ();
 FILLCELL_X2 FILLER_317_929 ();
 FILLCELL_X1 FILLER_317_931 ();
 FILLCELL_X8 FILLER_317_948 ();
 FILLCELL_X4 FILLER_317_956 ();
 FILLCELL_X1 FILLER_317_960 ();
 FILLCELL_X4 FILLER_317_965 ();
 FILLCELL_X1 FILLER_317_969 ();
 FILLCELL_X16 FILLER_317_972 ();
 FILLCELL_X8 FILLER_317_988 ();
 FILLCELL_X2 FILLER_317_996 ();
 FILLCELL_X16 FILLER_317_1000 ();
 FILLCELL_X8 FILLER_317_1016 ();
 FILLCELL_X2 FILLER_317_1040 ();
 FILLCELL_X8 FILLER_317_1046 ();
 FILLCELL_X2 FILLER_317_1070 ();
 FILLCELL_X16 FILLER_317_1104 ();
 FILLCELL_X8 FILLER_317_1120 ();
 FILLCELL_X2 FILLER_317_1128 ();
 FILLCELL_X32 FILLER_317_1149 ();
 FILLCELL_X2 FILLER_317_1181 ();
 FILLCELL_X32 FILLER_317_1203 ();
 FILLCELL_X16 FILLER_317_1235 ();
 FILLCELL_X8 FILLER_317_1251 ();
 FILLCELL_X4 FILLER_317_1259 ();
 FILLCELL_X4 FILLER_317_1264 ();
 FILLCELL_X1 FILLER_317_1290 ();
 FILLCELL_X32 FILLER_317_1296 ();
 FILLCELL_X32 FILLER_317_1328 ();
 FILLCELL_X32 FILLER_317_1360 ();
 FILLCELL_X32 FILLER_317_1392 ();
 FILLCELL_X32 FILLER_317_1424 ();
 FILLCELL_X32 FILLER_317_1456 ();
 FILLCELL_X32 FILLER_317_1488 ();
 FILLCELL_X32 FILLER_317_1520 ();
 FILLCELL_X32 FILLER_317_1552 ();
 FILLCELL_X32 FILLER_317_1584 ();
 FILLCELL_X32 FILLER_317_1616 ();
 FILLCELL_X32 FILLER_317_1648 ();
 FILLCELL_X32 FILLER_317_1680 ();
 FILLCELL_X32 FILLER_317_1712 ();
 FILLCELL_X32 FILLER_317_1744 ();
 FILLCELL_X32 FILLER_317_1776 ();
 FILLCELL_X32 FILLER_317_1808 ();
 FILLCELL_X32 FILLER_317_1840 ();
 FILLCELL_X32 FILLER_317_1872 ();
 FILLCELL_X32 FILLER_317_1904 ();
 FILLCELL_X32 FILLER_317_1936 ();
 FILLCELL_X32 FILLER_317_1968 ();
 FILLCELL_X32 FILLER_317_2000 ();
 FILLCELL_X32 FILLER_317_2032 ();
 FILLCELL_X32 FILLER_317_2064 ();
 FILLCELL_X32 FILLER_317_2096 ();
 FILLCELL_X32 FILLER_317_2128 ();
 FILLCELL_X32 FILLER_317_2160 ();
 FILLCELL_X32 FILLER_317_2192 ();
 FILLCELL_X32 FILLER_317_2224 ();
 FILLCELL_X32 FILLER_317_2256 ();
 FILLCELL_X32 FILLER_317_2288 ();
 FILLCELL_X32 FILLER_317_2320 ();
 FILLCELL_X32 FILLER_317_2352 ();
 FILLCELL_X32 FILLER_317_2384 ();
 FILLCELL_X16 FILLER_317_2416 ();
 FILLCELL_X4 FILLER_317_2432 ();
 FILLCELL_X32 FILLER_318_1 ();
 FILLCELL_X32 FILLER_318_33 ();
 FILLCELL_X32 FILLER_318_65 ();
 FILLCELL_X32 FILLER_318_97 ();
 FILLCELL_X32 FILLER_318_129 ();
 FILLCELL_X32 FILLER_318_161 ();
 FILLCELL_X32 FILLER_318_193 ();
 FILLCELL_X32 FILLER_318_225 ();
 FILLCELL_X32 FILLER_318_257 ();
 FILLCELL_X32 FILLER_318_289 ();
 FILLCELL_X32 FILLER_318_321 ();
 FILLCELL_X32 FILLER_318_353 ();
 FILLCELL_X32 FILLER_318_385 ();
 FILLCELL_X32 FILLER_318_417 ();
 FILLCELL_X32 FILLER_318_449 ();
 FILLCELL_X32 FILLER_318_481 ();
 FILLCELL_X32 FILLER_318_513 ();
 FILLCELL_X32 FILLER_318_545 ();
 FILLCELL_X32 FILLER_318_577 ();
 FILLCELL_X16 FILLER_318_609 ();
 FILLCELL_X4 FILLER_318_625 ();
 FILLCELL_X2 FILLER_318_629 ();
 FILLCELL_X32 FILLER_318_632 ();
 FILLCELL_X32 FILLER_318_664 ();
 FILLCELL_X32 FILLER_318_696 ();
 FILLCELL_X32 FILLER_318_728 ();
 FILLCELL_X32 FILLER_318_760 ();
 FILLCELL_X32 FILLER_318_792 ();
 FILLCELL_X32 FILLER_318_824 ();
 FILLCELL_X32 FILLER_318_856 ();
 FILLCELL_X32 FILLER_318_888 ();
 FILLCELL_X32 FILLER_318_920 ();
 FILLCELL_X8 FILLER_318_952 ();
 FILLCELL_X2 FILLER_318_960 ();
 FILLCELL_X32 FILLER_318_966 ();
 FILLCELL_X2 FILLER_318_998 ();
 FILLCELL_X16 FILLER_318_1002 ();
 FILLCELL_X8 FILLER_318_1018 ();
 FILLCELL_X16 FILLER_318_1042 ();
 FILLCELL_X8 FILLER_318_1058 ();
 FILLCELL_X2 FILLER_318_1066 ();
 FILLCELL_X1 FILLER_318_1068 ();
 FILLCELL_X2 FILLER_318_1073 ();
 FILLCELL_X32 FILLER_318_1079 ();
 FILLCELL_X4 FILLER_318_1111 ();
 FILLCELL_X1 FILLER_318_1115 ();
 FILLCELL_X16 FILLER_318_1120 ();
 FILLCELL_X2 FILLER_318_1136 ();
 FILLCELL_X1 FILLER_318_1138 ();
 FILLCELL_X8 FILLER_318_1142 ();
 FILLCELL_X4 FILLER_318_1150 ();
 FILLCELL_X2 FILLER_318_1154 ();
 FILLCELL_X32 FILLER_318_1160 ();
 FILLCELL_X4 FILLER_318_1195 ();
 FILLCELL_X2 FILLER_318_1199 ();
 FILLCELL_X1 FILLER_318_1201 ();
 FILLCELL_X32 FILLER_318_1227 ();
 FILLCELL_X8 FILLER_318_1259 ();
 FILLCELL_X32 FILLER_318_1295 ();
 FILLCELL_X32 FILLER_318_1327 ();
 FILLCELL_X32 FILLER_318_1359 ();
 FILLCELL_X32 FILLER_318_1391 ();
 FILLCELL_X32 FILLER_318_1423 ();
 FILLCELL_X32 FILLER_318_1455 ();
 FILLCELL_X32 FILLER_318_1487 ();
 FILLCELL_X32 FILLER_318_1519 ();
 FILLCELL_X32 FILLER_318_1551 ();
 FILLCELL_X32 FILLER_318_1583 ();
 FILLCELL_X32 FILLER_318_1615 ();
 FILLCELL_X32 FILLER_318_1647 ();
 FILLCELL_X32 FILLER_318_1679 ();
 FILLCELL_X32 FILLER_318_1711 ();
 FILLCELL_X32 FILLER_318_1743 ();
 FILLCELL_X32 FILLER_318_1775 ();
 FILLCELL_X32 FILLER_318_1807 ();
 FILLCELL_X32 FILLER_318_1839 ();
 FILLCELL_X16 FILLER_318_1871 ();
 FILLCELL_X4 FILLER_318_1887 ();
 FILLCELL_X2 FILLER_318_1891 ();
 FILLCELL_X1 FILLER_318_1893 ();
 FILLCELL_X32 FILLER_318_1895 ();
 FILLCELL_X32 FILLER_318_1927 ();
 FILLCELL_X32 FILLER_318_1959 ();
 FILLCELL_X32 FILLER_318_1991 ();
 FILLCELL_X32 FILLER_318_2023 ();
 FILLCELL_X32 FILLER_318_2055 ();
 FILLCELL_X32 FILLER_318_2087 ();
 FILLCELL_X32 FILLER_318_2119 ();
 FILLCELL_X32 FILLER_318_2151 ();
 FILLCELL_X32 FILLER_318_2183 ();
 FILLCELL_X32 FILLER_318_2215 ();
 FILLCELL_X32 FILLER_318_2247 ();
 FILLCELL_X32 FILLER_318_2279 ();
 FILLCELL_X32 FILLER_318_2311 ();
 FILLCELL_X32 FILLER_318_2343 ();
 FILLCELL_X32 FILLER_318_2375 ();
 FILLCELL_X16 FILLER_318_2407 ();
 FILLCELL_X8 FILLER_318_2423 ();
 FILLCELL_X4 FILLER_318_2431 ();
 FILLCELL_X1 FILLER_318_2435 ();
 FILLCELL_X32 FILLER_319_1 ();
 FILLCELL_X32 FILLER_319_33 ();
 FILLCELL_X32 FILLER_319_65 ();
 FILLCELL_X32 FILLER_319_97 ();
 FILLCELL_X32 FILLER_319_129 ();
 FILLCELL_X32 FILLER_319_161 ();
 FILLCELL_X32 FILLER_319_193 ();
 FILLCELL_X32 FILLER_319_225 ();
 FILLCELL_X32 FILLER_319_257 ();
 FILLCELL_X32 FILLER_319_289 ();
 FILLCELL_X32 FILLER_319_321 ();
 FILLCELL_X32 FILLER_319_353 ();
 FILLCELL_X32 FILLER_319_385 ();
 FILLCELL_X32 FILLER_319_417 ();
 FILLCELL_X32 FILLER_319_449 ();
 FILLCELL_X32 FILLER_319_481 ();
 FILLCELL_X32 FILLER_319_513 ();
 FILLCELL_X32 FILLER_319_545 ();
 FILLCELL_X32 FILLER_319_577 ();
 FILLCELL_X32 FILLER_319_609 ();
 FILLCELL_X32 FILLER_319_641 ();
 FILLCELL_X32 FILLER_319_673 ();
 FILLCELL_X32 FILLER_319_705 ();
 FILLCELL_X32 FILLER_319_737 ();
 FILLCELL_X32 FILLER_319_769 ();
 FILLCELL_X32 FILLER_319_801 ();
 FILLCELL_X32 FILLER_319_833 ();
 FILLCELL_X32 FILLER_319_865 ();
 FILLCELL_X32 FILLER_319_897 ();
 FILLCELL_X16 FILLER_319_929 ();
 FILLCELL_X8 FILLER_319_945 ();
 FILLCELL_X4 FILLER_319_953 ();
 FILLCELL_X2 FILLER_319_957 ();
 FILLCELL_X16 FILLER_319_973 ();
 FILLCELL_X8 FILLER_319_989 ();
 FILLCELL_X16 FILLER_319_1011 ();
 FILLCELL_X2 FILLER_319_1027 ();
 FILLCELL_X32 FILLER_319_1031 ();
 FILLCELL_X32 FILLER_319_1063 ();
 FILLCELL_X8 FILLER_319_1095 ();
 FILLCELL_X2 FILLER_319_1103 ();
 FILLCELL_X1 FILLER_319_1105 ();
 FILLCELL_X32 FILLER_319_1129 ();
 FILLCELL_X16 FILLER_319_1161 ();
 FILLCELL_X8 FILLER_319_1177 ();
 FILLCELL_X4 FILLER_319_1185 ();
 FILLCELL_X2 FILLER_319_1189 ();
 FILLCELL_X1 FILLER_319_1191 ();
 FILLCELL_X16 FILLER_319_1194 ();
 FILLCELL_X4 FILLER_319_1210 ();
 FILLCELL_X2 FILLER_319_1214 ();
 FILLCELL_X32 FILLER_319_1222 ();
 FILLCELL_X8 FILLER_319_1254 ();
 FILLCELL_X1 FILLER_319_1262 ();
 FILLCELL_X2 FILLER_319_1264 ();
 FILLCELL_X1 FILLER_319_1266 ();
 FILLCELL_X4 FILLER_319_1277 ();
 FILLCELL_X32 FILLER_319_1291 ();
 FILLCELL_X32 FILLER_319_1323 ();
 FILLCELL_X32 FILLER_319_1355 ();
 FILLCELL_X32 FILLER_319_1387 ();
 FILLCELL_X32 FILLER_319_1419 ();
 FILLCELL_X32 FILLER_319_1451 ();
 FILLCELL_X32 FILLER_319_1483 ();
 FILLCELL_X32 FILLER_319_1515 ();
 FILLCELL_X32 FILLER_319_1547 ();
 FILLCELL_X32 FILLER_319_1579 ();
 FILLCELL_X32 FILLER_319_1611 ();
 FILLCELL_X32 FILLER_319_1643 ();
 FILLCELL_X32 FILLER_319_1675 ();
 FILLCELL_X32 FILLER_319_1707 ();
 FILLCELL_X32 FILLER_319_1739 ();
 FILLCELL_X32 FILLER_319_1771 ();
 FILLCELL_X32 FILLER_319_1803 ();
 FILLCELL_X32 FILLER_319_1835 ();
 FILLCELL_X32 FILLER_319_1867 ();
 FILLCELL_X32 FILLER_319_1899 ();
 FILLCELL_X32 FILLER_319_1931 ();
 FILLCELL_X32 FILLER_319_1963 ();
 FILLCELL_X32 FILLER_319_1995 ();
 FILLCELL_X32 FILLER_319_2027 ();
 FILLCELL_X32 FILLER_319_2059 ();
 FILLCELL_X32 FILLER_319_2091 ();
 FILLCELL_X32 FILLER_319_2123 ();
 FILLCELL_X32 FILLER_319_2155 ();
 FILLCELL_X32 FILLER_319_2187 ();
 FILLCELL_X32 FILLER_319_2219 ();
 FILLCELL_X32 FILLER_319_2251 ();
 FILLCELL_X32 FILLER_319_2283 ();
 FILLCELL_X32 FILLER_319_2315 ();
 FILLCELL_X32 FILLER_319_2347 ();
 FILLCELL_X32 FILLER_319_2379 ();
 FILLCELL_X16 FILLER_319_2411 ();
 FILLCELL_X8 FILLER_319_2427 ();
 FILLCELL_X1 FILLER_319_2435 ();
 FILLCELL_X32 FILLER_320_1 ();
 FILLCELL_X32 FILLER_320_33 ();
 FILLCELL_X32 FILLER_320_65 ();
 FILLCELL_X32 FILLER_320_97 ();
 FILLCELL_X32 FILLER_320_129 ();
 FILLCELL_X32 FILLER_320_161 ();
 FILLCELL_X32 FILLER_320_193 ();
 FILLCELL_X32 FILLER_320_225 ();
 FILLCELL_X32 FILLER_320_257 ();
 FILLCELL_X32 FILLER_320_289 ();
 FILLCELL_X32 FILLER_320_321 ();
 FILLCELL_X32 FILLER_320_353 ();
 FILLCELL_X32 FILLER_320_385 ();
 FILLCELL_X32 FILLER_320_417 ();
 FILLCELL_X32 FILLER_320_449 ();
 FILLCELL_X32 FILLER_320_481 ();
 FILLCELL_X32 FILLER_320_513 ();
 FILLCELL_X32 FILLER_320_545 ();
 FILLCELL_X32 FILLER_320_577 ();
 FILLCELL_X16 FILLER_320_609 ();
 FILLCELL_X4 FILLER_320_625 ();
 FILLCELL_X2 FILLER_320_629 ();
 FILLCELL_X32 FILLER_320_632 ();
 FILLCELL_X32 FILLER_320_664 ();
 FILLCELL_X32 FILLER_320_696 ();
 FILLCELL_X32 FILLER_320_728 ();
 FILLCELL_X32 FILLER_320_760 ();
 FILLCELL_X32 FILLER_320_792 ();
 FILLCELL_X32 FILLER_320_824 ();
 FILLCELL_X32 FILLER_320_856 ();
 FILLCELL_X32 FILLER_320_888 ();
 FILLCELL_X32 FILLER_320_920 ();
 FILLCELL_X16 FILLER_320_952 ();
 FILLCELL_X1 FILLER_320_968 ();
 FILLCELL_X8 FILLER_320_985 ();
 FILLCELL_X4 FILLER_320_993 ();
 FILLCELL_X1 FILLER_320_997 ();
 FILLCELL_X16 FILLER_320_1018 ();
 FILLCELL_X4 FILLER_320_1034 ();
 FILLCELL_X2 FILLER_320_1038 ();
 FILLCELL_X32 FILLER_320_1059 ();
 FILLCELL_X4 FILLER_320_1091 ();
 FILLCELL_X2 FILLER_320_1095 ();
 FILLCELL_X16 FILLER_320_1099 ();
 FILLCELL_X32 FILLER_320_1119 ();
 FILLCELL_X2 FILLER_320_1151 ();
 FILLCELL_X8 FILLER_320_1162 ();
 FILLCELL_X1 FILLER_320_1170 ();
 FILLCELL_X8 FILLER_320_1181 ();
 FILLCELL_X1 FILLER_320_1189 ();
 FILLCELL_X8 FILLER_320_1196 ();
 FILLCELL_X2 FILLER_320_1204 ();
 FILLCELL_X1 FILLER_320_1206 ();
 FILLCELL_X4 FILLER_320_1212 ();
 FILLCELL_X2 FILLER_320_1216 ();
 FILLCELL_X1 FILLER_320_1218 ();
 FILLCELL_X32 FILLER_320_1224 ();
 FILLCELL_X16 FILLER_320_1256 ();
 FILLCELL_X4 FILLER_320_1272 ();
 FILLCELL_X1 FILLER_320_1276 ();
 FILLCELL_X32 FILLER_320_1284 ();
 FILLCELL_X32 FILLER_320_1316 ();
 FILLCELL_X32 FILLER_320_1348 ();
 FILLCELL_X32 FILLER_320_1380 ();
 FILLCELL_X32 FILLER_320_1412 ();
 FILLCELL_X32 FILLER_320_1444 ();
 FILLCELL_X32 FILLER_320_1476 ();
 FILLCELL_X32 FILLER_320_1508 ();
 FILLCELL_X32 FILLER_320_1540 ();
 FILLCELL_X32 FILLER_320_1572 ();
 FILLCELL_X32 FILLER_320_1604 ();
 FILLCELL_X32 FILLER_320_1636 ();
 FILLCELL_X32 FILLER_320_1668 ();
 FILLCELL_X32 FILLER_320_1700 ();
 FILLCELL_X32 FILLER_320_1732 ();
 FILLCELL_X32 FILLER_320_1764 ();
 FILLCELL_X32 FILLER_320_1796 ();
 FILLCELL_X32 FILLER_320_1828 ();
 FILLCELL_X32 FILLER_320_1860 ();
 FILLCELL_X2 FILLER_320_1892 ();
 FILLCELL_X32 FILLER_320_1895 ();
 FILLCELL_X32 FILLER_320_1927 ();
 FILLCELL_X32 FILLER_320_1959 ();
 FILLCELL_X32 FILLER_320_1991 ();
 FILLCELL_X32 FILLER_320_2023 ();
 FILLCELL_X32 FILLER_320_2055 ();
 FILLCELL_X32 FILLER_320_2087 ();
 FILLCELL_X32 FILLER_320_2119 ();
 FILLCELL_X32 FILLER_320_2151 ();
 FILLCELL_X32 FILLER_320_2183 ();
 FILLCELL_X32 FILLER_320_2215 ();
 FILLCELL_X32 FILLER_320_2247 ();
 FILLCELL_X32 FILLER_320_2279 ();
 FILLCELL_X32 FILLER_320_2311 ();
 FILLCELL_X32 FILLER_320_2343 ();
 FILLCELL_X32 FILLER_320_2375 ();
 FILLCELL_X16 FILLER_320_2407 ();
 FILLCELL_X8 FILLER_320_2423 ();
 FILLCELL_X4 FILLER_320_2431 ();
 FILLCELL_X1 FILLER_320_2435 ();
 FILLCELL_X32 FILLER_321_1 ();
 FILLCELL_X32 FILLER_321_33 ();
 FILLCELL_X32 FILLER_321_65 ();
 FILLCELL_X32 FILLER_321_97 ();
 FILLCELL_X32 FILLER_321_129 ();
 FILLCELL_X32 FILLER_321_161 ();
 FILLCELL_X32 FILLER_321_193 ();
 FILLCELL_X32 FILLER_321_225 ();
 FILLCELL_X32 FILLER_321_257 ();
 FILLCELL_X32 FILLER_321_289 ();
 FILLCELL_X32 FILLER_321_321 ();
 FILLCELL_X32 FILLER_321_353 ();
 FILLCELL_X32 FILLER_321_385 ();
 FILLCELL_X32 FILLER_321_417 ();
 FILLCELL_X32 FILLER_321_449 ();
 FILLCELL_X32 FILLER_321_481 ();
 FILLCELL_X32 FILLER_321_513 ();
 FILLCELL_X32 FILLER_321_545 ();
 FILLCELL_X32 FILLER_321_577 ();
 FILLCELL_X32 FILLER_321_609 ();
 FILLCELL_X32 FILLER_321_641 ();
 FILLCELL_X32 FILLER_321_673 ();
 FILLCELL_X32 FILLER_321_705 ();
 FILLCELL_X32 FILLER_321_737 ();
 FILLCELL_X32 FILLER_321_769 ();
 FILLCELL_X32 FILLER_321_801 ();
 FILLCELL_X32 FILLER_321_833 ();
 FILLCELL_X32 FILLER_321_865 ();
 FILLCELL_X32 FILLER_321_897 ();
 FILLCELL_X4 FILLER_321_929 ();
 FILLCELL_X1 FILLER_321_933 ();
 FILLCELL_X4 FILLER_321_968 ();
 FILLCELL_X4 FILLER_321_982 ();
 FILLCELL_X32 FILLER_321_990 ();
 FILLCELL_X16 FILLER_321_1022 ();
 FILLCELL_X1 FILLER_321_1038 ();
 FILLCELL_X8 FILLER_321_1043 ();
 FILLCELL_X4 FILLER_321_1051 ();
 FILLCELL_X2 FILLER_321_1055 ();
 FILLCELL_X1 FILLER_321_1057 ();
 FILLCELL_X1 FILLER_321_1062 ();
 FILLCELL_X4 FILLER_321_1079 ();
 FILLCELL_X32 FILLER_321_1097 ();
 FILLCELL_X8 FILLER_321_1129 ();
 FILLCELL_X4 FILLER_321_1137 ();
 FILLCELL_X2 FILLER_321_1141 ();
 FILLCELL_X1 FILLER_321_1143 ();
 FILLCELL_X4 FILLER_321_1173 ();
 FILLCELL_X2 FILLER_321_1177 ();
 FILLCELL_X8 FILLER_321_1181 ();
 FILLCELL_X4 FILLER_321_1189 ();
 FILLCELL_X1 FILLER_321_1193 ();
 FILLCELL_X2 FILLER_321_1197 ();
 FILLCELL_X1 FILLER_321_1199 ();
 FILLCELL_X2 FILLER_321_1205 ();
 FILLCELL_X1 FILLER_321_1213 ();
 FILLCELL_X16 FILLER_321_1217 ();
 FILLCELL_X2 FILLER_321_1233 ();
 FILLCELL_X1 FILLER_321_1235 ();
 FILLCELL_X16 FILLER_321_1243 ();
 FILLCELL_X4 FILLER_321_1259 ();
 FILLCELL_X8 FILLER_321_1264 ();
 FILLCELL_X2 FILLER_321_1272 ();
 FILLCELL_X32 FILLER_321_1277 ();
 FILLCELL_X32 FILLER_321_1309 ();
 FILLCELL_X32 FILLER_321_1341 ();
 FILLCELL_X32 FILLER_321_1373 ();
 FILLCELL_X32 FILLER_321_1405 ();
 FILLCELL_X32 FILLER_321_1437 ();
 FILLCELL_X32 FILLER_321_1469 ();
 FILLCELL_X32 FILLER_321_1501 ();
 FILLCELL_X32 FILLER_321_1533 ();
 FILLCELL_X32 FILLER_321_1565 ();
 FILLCELL_X32 FILLER_321_1597 ();
 FILLCELL_X32 FILLER_321_1629 ();
 FILLCELL_X32 FILLER_321_1661 ();
 FILLCELL_X32 FILLER_321_1693 ();
 FILLCELL_X32 FILLER_321_1725 ();
 FILLCELL_X32 FILLER_321_1757 ();
 FILLCELL_X32 FILLER_321_1789 ();
 FILLCELL_X32 FILLER_321_1821 ();
 FILLCELL_X32 FILLER_321_1853 ();
 FILLCELL_X32 FILLER_321_1885 ();
 FILLCELL_X32 FILLER_321_1917 ();
 FILLCELL_X32 FILLER_321_1949 ();
 FILLCELL_X32 FILLER_321_1981 ();
 FILLCELL_X32 FILLER_321_2013 ();
 FILLCELL_X32 FILLER_321_2045 ();
 FILLCELL_X32 FILLER_321_2077 ();
 FILLCELL_X32 FILLER_321_2109 ();
 FILLCELL_X32 FILLER_321_2141 ();
 FILLCELL_X32 FILLER_321_2173 ();
 FILLCELL_X32 FILLER_321_2205 ();
 FILLCELL_X32 FILLER_321_2237 ();
 FILLCELL_X32 FILLER_321_2269 ();
 FILLCELL_X32 FILLER_321_2301 ();
 FILLCELL_X32 FILLER_321_2333 ();
 FILLCELL_X32 FILLER_321_2365 ();
 FILLCELL_X32 FILLER_321_2397 ();
 FILLCELL_X4 FILLER_321_2429 ();
 FILLCELL_X2 FILLER_321_2433 ();
 FILLCELL_X1 FILLER_321_2435 ();
 FILLCELL_X32 FILLER_322_1 ();
 FILLCELL_X32 FILLER_322_33 ();
 FILLCELL_X32 FILLER_322_65 ();
 FILLCELL_X32 FILLER_322_97 ();
 FILLCELL_X32 FILLER_322_129 ();
 FILLCELL_X32 FILLER_322_161 ();
 FILLCELL_X32 FILLER_322_193 ();
 FILLCELL_X32 FILLER_322_225 ();
 FILLCELL_X32 FILLER_322_257 ();
 FILLCELL_X32 FILLER_322_289 ();
 FILLCELL_X32 FILLER_322_321 ();
 FILLCELL_X32 FILLER_322_353 ();
 FILLCELL_X32 FILLER_322_385 ();
 FILLCELL_X32 FILLER_322_417 ();
 FILLCELL_X32 FILLER_322_449 ();
 FILLCELL_X32 FILLER_322_481 ();
 FILLCELL_X32 FILLER_322_513 ();
 FILLCELL_X32 FILLER_322_545 ();
 FILLCELL_X32 FILLER_322_577 ();
 FILLCELL_X16 FILLER_322_609 ();
 FILLCELL_X4 FILLER_322_625 ();
 FILLCELL_X2 FILLER_322_629 ();
 FILLCELL_X32 FILLER_322_632 ();
 FILLCELL_X32 FILLER_322_664 ();
 FILLCELL_X32 FILLER_322_696 ();
 FILLCELL_X32 FILLER_322_728 ();
 FILLCELL_X32 FILLER_322_760 ();
 FILLCELL_X32 FILLER_322_792 ();
 FILLCELL_X32 FILLER_322_824 ();
 FILLCELL_X32 FILLER_322_856 ();
 FILLCELL_X32 FILLER_322_888 ();
 FILLCELL_X32 FILLER_322_920 ();
 FILLCELL_X8 FILLER_322_952 ();
 FILLCELL_X4 FILLER_322_960 ();
 FILLCELL_X4 FILLER_322_968 ();
 FILLCELL_X16 FILLER_322_976 ();
 FILLCELL_X8 FILLER_322_992 ();
 FILLCELL_X4 FILLER_322_1000 ();
 FILLCELL_X8 FILLER_322_1008 ();
 FILLCELL_X2 FILLER_322_1016 ();
 FILLCELL_X8 FILLER_322_1020 ();
 FILLCELL_X4 FILLER_322_1028 ();
 FILLCELL_X1 FILLER_322_1032 ();
 FILLCELL_X8 FILLER_322_1049 ();
 FILLCELL_X4 FILLER_322_1081 ();
 FILLCELL_X16 FILLER_322_1101 ();
 FILLCELL_X4 FILLER_322_1117 ();
 FILLCELL_X8 FILLER_322_1134 ();
 FILLCELL_X2 FILLER_322_1142 ();
 FILLCELL_X16 FILLER_322_1148 ();
 FILLCELL_X4 FILLER_322_1168 ();
 FILLCELL_X1 FILLER_322_1172 ();
 FILLCELL_X8 FILLER_322_1177 ();
 FILLCELL_X4 FILLER_322_1185 ();
 FILLCELL_X1 FILLER_322_1189 ();
 FILLCELL_X1 FILLER_322_1212 ();
 FILLCELL_X4 FILLER_322_1219 ();
 FILLCELL_X1 FILLER_322_1236 ();
 FILLCELL_X1 FILLER_322_1240 ();
 FILLCELL_X2 FILLER_322_1243 ();
 FILLCELL_X32 FILLER_322_1254 ();
 FILLCELL_X32 FILLER_322_1286 ();
 FILLCELL_X32 FILLER_322_1318 ();
 FILLCELL_X32 FILLER_322_1350 ();
 FILLCELL_X32 FILLER_322_1382 ();
 FILLCELL_X32 FILLER_322_1414 ();
 FILLCELL_X32 FILLER_322_1446 ();
 FILLCELL_X32 FILLER_322_1478 ();
 FILLCELL_X32 FILLER_322_1510 ();
 FILLCELL_X32 FILLER_322_1542 ();
 FILLCELL_X32 FILLER_322_1574 ();
 FILLCELL_X32 FILLER_322_1606 ();
 FILLCELL_X32 FILLER_322_1638 ();
 FILLCELL_X32 FILLER_322_1670 ();
 FILLCELL_X32 FILLER_322_1702 ();
 FILLCELL_X32 FILLER_322_1734 ();
 FILLCELL_X32 FILLER_322_1766 ();
 FILLCELL_X32 FILLER_322_1798 ();
 FILLCELL_X32 FILLER_322_1830 ();
 FILLCELL_X32 FILLER_322_1862 ();
 FILLCELL_X32 FILLER_322_1895 ();
 FILLCELL_X32 FILLER_322_1927 ();
 FILLCELL_X32 FILLER_322_1959 ();
 FILLCELL_X32 FILLER_322_1991 ();
 FILLCELL_X32 FILLER_322_2023 ();
 FILLCELL_X32 FILLER_322_2055 ();
 FILLCELL_X32 FILLER_322_2087 ();
 FILLCELL_X32 FILLER_322_2119 ();
 FILLCELL_X32 FILLER_322_2151 ();
 FILLCELL_X32 FILLER_322_2183 ();
 FILLCELL_X32 FILLER_322_2215 ();
 FILLCELL_X32 FILLER_322_2247 ();
 FILLCELL_X32 FILLER_322_2279 ();
 FILLCELL_X32 FILLER_322_2311 ();
 FILLCELL_X32 FILLER_322_2343 ();
 FILLCELL_X32 FILLER_322_2375 ();
 FILLCELL_X16 FILLER_322_2407 ();
 FILLCELL_X8 FILLER_322_2423 ();
 FILLCELL_X4 FILLER_322_2431 ();
 FILLCELL_X1 FILLER_322_2435 ();
 FILLCELL_X32 FILLER_323_1 ();
 FILLCELL_X32 FILLER_323_33 ();
 FILLCELL_X32 FILLER_323_65 ();
 FILLCELL_X32 FILLER_323_97 ();
 FILLCELL_X32 FILLER_323_129 ();
 FILLCELL_X32 FILLER_323_161 ();
 FILLCELL_X32 FILLER_323_193 ();
 FILLCELL_X32 FILLER_323_225 ();
 FILLCELL_X32 FILLER_323_257 ();
 FILLCELL_X32 FILLER_323_289 ();
 FILLCELL_X32 FILLER_323_321 ();
 FILLCELL_X32 FILLER_323_353 ();
 FILLCELL_X32 FILLER_323_385 ();
 FILLCELL_X32 FILLER_323_417 ();
 FILLCELL_X32 FILLER_323_449 ();
 FILLCELL_X32 FILLER_323_481 ();
 FILLCELL_X32 FILLER_323_513 ();
 FILLCELL_X32 FILLER_323_545 ();
 FILLCELL_X32 FILLER_323_577 ();
 FILLCELL_X32 FILLER_323_609 ();
 FILLCELL_X32 FILLER_323_641 ();
 FILLCELL_X32 FILLER_323_673 ();
 FILLCELL_X32 FILLER_323_705 ();
 FILLCELL_X32 FILLER_323_737 ();
 FILLCELL_X32 FILLER_323_769 ();
 FILLCELL_X32 FILLER_323_801 ();
 FILLCELL_X32 FILLER_323_833 ();
 FILLCELL_X32 FILLER_323_865 ();
 FILLCELL_X32 FILLER_323_897 ();
 FILLCELL_X32 FILLER_323_929 ();
 FILLCELL_X16 FILLER_323_961 ();
 FILLCELL_X1 FILLER_323_977 ();
 FILLCELL_X4 FILLER_323_998 ();
 FILLCELL_X1 FILLER_323_1002 ();
 FILLCELL_X16 FILLER_323_1013 ();
 FILLCELL_X8 FILLER_323_1029 ();
 FILLCELL_X2 FILLER_323_1037 ();
 FILLCELL_X1 FILLER_323_1039 ();
 FILLCELL_X16 FILLER_323_1044 ();
 FILLCELL_X8 FILLER_323_1060 ();
 FILLCELL_X32 FILLER_323_1072 ();
 FILLCELL_X32 FILLER_323_1104 ();
 FILLCELL_X8 FILLER_323_1136 ();
 FILLCELL_X1 FILLER_323_1144 ();
 FILLCELL_X16 FILLER_323_1151 ();
 FILLCELL_X4 FILLER_323_1167 ();
 FILLCELL_X1 FILLER_323_1171 ();
 FILLCELL_X32 FILLER_323_1182 ();
 FILLCELL_X4 FILLER_323_1214 ();
 FILLCELL_X1 FILLER_323_1218 ();
 FILLCELL_X32 FILLER_323_1264 ();
 FILLCELL_X32 FILLER_323_1296 ();
 FILLCELL_X32 FILLER_323_1328 ();
 FILLCELL_X32 FILLER_323_1360 ();
 FILLCELL_X32 FILLER_323_1392 ();
 FILLCELL_X32 FILLER_323_1424 ();
 FILLCELL_X32 FILLER_323_1456 ();
 FILLCELL_X32 FILLER_323_1488 ();
 FILLCELL_X32 FILLER_323_1520 ();
 FILLCELL_X32 FILLER_323_1552 ();
 FILLCELL_X32 FILLER_323_1584 ();
 FILLCELL_X32 FILLER_323_1616 ();
 FILLCELL_X32 FILLER_323_1648 ();
 FILLCELL_X32 FILLER_323_1680 ();
 FILLCELL_X32 FILLER_323_1712 ();
 FILLCELL_X32 FILLER_323_1744 ();
 FILLCELL_X32 FILLER_323_1776 ();
 FILLCELL_X32 FILLER_323_1808 ();
 FILLCELL_X32 FILLER_323_1840 ();
 FILLCELL_X32 FILLER_323_1872 ();
 FILLCELL_X32 FILLER_323_1904 ();
 FILLCELL_X32 FILLER_323_1936 ();
 FILLCELL_X32 FILLER_323_1968 ();
 FILLCELL_X32 FILLER_323_2000 ();
 FILLCELL_X32 FILLER_323_2032 ();
 FILLCELL_X32 FILLER_323_2064 ();
 FILLCELL_X32 FILLER_323_2096 ();
 FILLCELL_X32 FILLER_323_2128 ();
 FILLCELL_X32 FILLER_323_2160 ();
 FILLCELL_X32 FILLER_323_2192 ();
 FILLCELL_X32 FILLER_323_2224 ();
 FILLCELL_X32 FILLER_323_2256 ();
 FILLCELL_X32 FILLER_323_2288 ();
 FILLCELL_X32 FILLER_323_2320 ();
 FILLCELL_X32 FILLER_323_2352 ();
 FILLCELL_X32 FILLER_323_2384 ();
 FILLCELL_X16 FILLER_323_2416 ();
 FILLCELL_X4 FILLER_323_2432 ();
 FILLCELL_X32 FILLER_324_1 ();
 FILLCELL_X32 FILLER_324_33 ();
 FILLCELL_X32 FILLER_324_65 ();
 FILLCELL_X32 FILLER_324_97 ();
 FILLCELL_X32 FILLER_324_129 ();
 FILLCELL_X32 FILLER_324_161 ();
 FILLCELL_X32 FILLER_324_193 ();
 FILLCELL_X32 FILLER_324_225 ();
 FILLCELL_X32 FILLER_324_257 ();
 FILLCELL_X32 FILLER_324_289 ();
 FILLCELL_X32 FILLER_324_321 ();
 FILLCELL_X32 FILLER_324_353 ();
 FILLCELL_X32 FILLER_324_385 ();
 FILLCELL_X32 FILLER_324_417 ();
 FILLCELL_X32 FILLER_324_449 ();
 FILLCELL_X32 FILLER_324_481 ();
 FILLCELL_X32 FILLER_324_513 ();
 FILLCELL_X32 FILLER_324_545 ();
 FILLCELL_X32 FILLER_324_577 ();
 FILLCELL_X16 FILLER_324_609 ();
 FILLCELL_X4 FILLER_324_625 ();
 FILLCELL_X2 FILLER_324_629 ();
 FILLCELL_X32 FILLER_324_632 ();
 FILLCELL_X32 FILLER_324_664 ();
 FILLCELL_X32 FILLER_324_696 ();
 FILLCELL_X32 FILLER_324_728 ();
 FILLCELL_X32 FILLER_324_760 ();
 FILLCELL_X32 FILLER_324_792 ();
 FILLCELL_X32 FILLER_324_824 ();
 FILLCELL_X32 FILLER_324_856 ();
 FILLCELL_X32 FILLER_324_888 ();
 FILLCELL_X32 FILLER_324_920 ();
 FILLCELL_X32 FILLER_324_952 ();
 FILLCELL_X4 FILLER_324_984 ();
 FILLCELL_X1 FILLER_324_988 ();
 FILLCELL_X8 FILLER_324_993 ();
 FILLCELL_X2 FILLER_324_1001 ();
 FILLCELL_X32 FILLER_324_1019 ();
 FILLCELL_X32 FILLER_324_1051 ();
 FILLCELL_X32 FILLER_324_1083 ();
 FILLCELL_X16 FILLER_324_1115 ();
 FILLCELL_X8 FILLER_324_1131 ();
 FILLCELL_X4 FILLER_324_1139 ();
 FILLCELL_X2 FILLER_324_1143 ();
 FILLCELL_X16 FILLER_324_1147 ();
 FILLCELL_X8 FILLER_324_1163 ();
 FILLCELL_X2 FILLER_324_1171 ();
 FILLCELL_X1 FILLER_324_1173 ();
 FILLCELL_X32 FILLER_324_1176 ();
 FILLCELL_X16 FILLER_324_1208 ();
 FILLCELL_X2 FILLER_324_1224 ();
 FILLCELL_X1 FILLER_324_1226 ();
 FILLCELL_X16 FILLER_324_1232 ();
 FILLCELL_X4 FILLER_324_1248 ();
 FILLCELL_X2 FILLER_324_1252 ();
 FILLCELL_X32 FILLER_324_1262 ();
 FILLCELL_X32 FILLER_324_1294 ();
 FILLCELL_X32 FILLER_324_1326 ();
 FILLCELL_X32 FILLER_324_1358 ();
 FILLCELL_X32 FILLER_324_1390 ();
 FILLCELL_X32 FILLER_324_1422 ();
 FILLCELL_X32 FILLER_324_1454 ();
 FILLCELL_X32 FILLER_324_1486 ();
 FILLCELL_X32 FILLER_324_1518 ();
 FILLCELL_X32 FILLER_324_1550 ();
 FILLCELL_X32 FILLER_324_1582 ();
 FILLCELL_X32 FILLER_324_1614 ();
 FILLCELL_X32 FILLER_324_1646 ();
 FILLCELL_X32 FILLER_324_1678 ();
 FILLCELL_X32 FILLER_324_1710 ();
 FILLCELL_X32 FILLER_324_1742 ();
 FILLCELL_X32 FILLER_324_1774 ();
 FILLCELL_X32 FILLER_324_1806 ();
 FILLCELL_X32 FILLER_324_1838 ();
 FILLCELL_X16 FILLER_324_1870 ();
 FILLCELL_X8 FILLER_324_1886 ();
 FILLCELL_X32 FILLER_324_1895 ();
 FILLCELL_X32 FILLER_324_1927 ();
 FILLCELL_X32 FILLER_324_1959 ();
 FILLCELL_X32 FILLER_324_1991 ();
 FILLCELL_X32 FILLER_324_2023 ();
 FILLCELL_X32 FILLER_324_2055 ();
 FILLCELL_X32 FILLER_324_2087 ();
 FILLCELL_X32 FILLER_324_2119 ();
 FILLCELL_X32 FILLER_324_2151 ();
 FILLCELL_X32 FILLER_324_2183 ();
 FILLCELL_X32 FILLER_324_2215 ();
 FILLCELL_X32 FILLER_324_2247 ();
 FILLCELL_X32 FILLER_324_2279 ();
 FILLCELL_X32 FILLER_324_2311 ();
 FILLCELL_X32 FILLER_324_2343 ();
 FILLCELL_X32 FILLER_324_2375 ();
 FILLCELL_X16 FILLER_324_2407 ();
 FILLCELL_X8 FILLER_324_2423 ();
 FILLCELL_X4 FILLER_324_2431 ();
 FILLCELL_X1 FILLER_324_2435 ();
 FILLCELL_X32 FILLER_325_1 ();
 FILLCELL_X32 FILLER_325_33 ();
 FILLCELL_X32 FILLER_325_65 ();
 FILLCELL_X32 FILLER_325_97 ();
 FILLCELL_X32 FILLER_325_129 ();
 FILLCELL_X32 FILLER_325_161 ();
 FILLCELL_X32 FILLER_325_193 ();
 FILLCELL_X32 FILLER_325_225 ();
 FILLCELL_X32 FILLER_325_257 ();
 FILLCELL_X32 FILLER_325_289 ();
 FILLCELL_X32 FILLER_325_321 ();
 FILLCELL_X32 FILLER_325_353 ();
 FILLCELL_X32 FILLER_325_385 ();
 FILLCELL_X32 FILLER_325_417 ();
 FILLCELL_X32 FILLER_325_449 ();
 FILLCELL_X32 FILLER_325_481 ();
 FILLCELL_X32 FILLER_325_513 ();
 FILLCELL_X32 FILLER_325_545 ();
 FILLCELL_X32 FILLER_325_577 ();
 FILLCELL_X32 FILLER_325_609 ();
 FILLCELL_X32 FILLER_325_641 ();
 FILLCELL_X32 FILLER_325_673 ();
 FILLCELL_X32 FILLER_325_705 ();
 FILLCELL_X32 FILLER_325_737 ();
 FILLCELL_X32 FILLER_325_769 ();
 FILLCELL_X32 FILLER_325_801 ();
 FILLCELL_X32 FILLER_325_833 ();
 FILLCELL_X32 FILLER_325_865 ();
 FILLCELL_X32 FILLER_325_897 ();
 FILLCELL_X32 FILLER_325_929 ();
 FILLCELL_X32 FILLER_325_961 ();
 FILLCELL_X8 FILLER_325_993 ();
 FILLCELL_X4 FILLER_325_1001 ();
 FILLCELL_X2 FILLER_325_1005 ();
 FILLCELL_X1 FILLER_325_1007 ();
 FILLCELL_X32 FILLER_325_1012 ();
 FILLCELL_X16 FILLER_325_1044 ();
 FILLCELL_X8 FILLER_325_1060 ();
 FILLCELL_X2 FILLER_325_1068 ();
 FILLCELL_X1 FILLER_325_1070 ();
 FILLCELL_X32 FILLER_325_1073 ();
 FILLCELL_X32 FILLER_325_1105 ();
 FILLCELL_X4 FILLER_325_1137 ();
 FILLCELL_X2 FILLER_325_1141 ();
 FILLCELL_X1 FILLER_325_1143 ();
 FILLCELL_X16 FILLER_325_1151 ();
 FILLCELL_X8 FILLER_325_1167 ();
 FILLCELL_X8 FILLER_325_1179 ();
 FILLCELL_X4 FILLER_325_1187 ();
 FILLCELL_X2 FILLER_325_1191 ();
 FILLCELL_X1 FILLER_325_1193 ();
 FILLCELL_X1 FILLER_325_1196 ();
 FILLCELL_X32 FILLER_325_1207 ();
 FILLCELL_X8 FILLER_325_1239 ();
 FILLCELL_X2 FILLER_325_1247 ();
 FILLCELL_X1 FILLER_325_1249 ();
 FILLCELL_X8 FILLER_325_1254 ();
 FILLCELL_X1 FILLER_325_1262 ();
 FILLCELL_X1 FILLER_325_1264 ();
 FILLCELL_X32 FILLER_325_1287 ();
 FILLCELL_X32 FILLER_325_1319 ();
 FILLCELL_X32 FILLER_325_1351 ();
 FILLCELL_X32 FILLER_325_1383 ();
 FILLCELL_X32 FILLER_325_1415 ();
 FILLCELL_X32 FILLER_325_1447 ();
 FILLCELL_X32 FILLER_325_1479 ();
 FILLCELL_X32 FILLER_325_1511 ();
 FILLCELL_X32 FILLER_325_1543 ();
 FILLCELL_X32 FILLER_325_1575 ();
 FILLCELL_X32 FILLER_325_1607 ();
 FILLCELL_X32 FILLER_325_1639 ();
 FILLCELL_X32 FILLER_325_1671 ();
 FILLCELL_X32 FILLER_325_1703 ();
 FILLCELL_X32 FILLER_325_1735 ();
 FILLCELL_X32 FILLER_325_1767 ();
 FILLCELL_X32 FILLER_325_1799 ();
 FILLCELL_X32 FILLER_325_1831 ();
 FILLCELL_X32 FILLER_325_1863 ();
 FILLCELL_X32 FILLER_325_1895 ();
 FILLCELL_X32 FILLER_325_1927 ();
 FILLCELL_X32 FILLER_325_1959 ();
 FILLCELL_X32 FILLER_325_1991 ();
 FILLCELL_X32 FILLER_325_2023 ();
 FILLCELL_X32 FILLER_325_2055 ();
 FILLCELL_X32 FILLER_325_2087 ();
 FILLCELL_X32 FILLER_325_2119 ();
 FILLCELL_X32 FILLER_325_2151 ();
 FILLCELL_X32 FILLER_325_2183 ();
 FILLCELL_X32 FILLER_325_2215 ();
 FILLCELL_X32 FILLER_325_2247 ();
 FILLCELL_X32 FILLER_325_2279 ();
 FILLCELL_X32 FILLER_325_2311 ();
 FILLCELL_X32 FILLER_325_2343 ();
 FILLCELL_X32 FILLER_325_2375 ();
 FILLCELL_X16 FILLER_325_2407 ();
 FILLCELL_X8 FILLER_325_2423 ();
 FILLCELL_X4 FILLER_325_2431 ();
 FILLCELL_X1 FILLER_325_2435 ();
 FILLCELL_X32 FILLER_326_1 ();
 FILLCELL_X32 FILLER_326_33 ();
 FILLCELL_X32 FILLER_326_65 ();
 FILLCELL_X32 FILLER_326_97 ();
 FILLCELL_X32 FILLER_326_129 ();
 FILLCELL_X32 FILLER_326_161 ();
 FILLCELL_X32 FILLER_326_193 ();
 FILLCELL_X32 FILLER_326_225 ();
 FILLCELL_X32 FILLER_326_257 ();
 FILLCELL_X32 FILLER_326_289 ();
 FILLCELL_X32 FILLER_326_321 ();
 FILLCELL_X32 FILLER_326_353 ();
 FILLCELL_X32 FILLER_326_385 ();
 FILLCELL_X32 FILLER_326_417 ();
 FILLCELL_X32 FILLER_326_449 ();
 FILLCELL_X32 FILLER_326_481 ();
 FILLCELL_X32 FILLER_326_513 ();
 FILLCELL_X32 FILLER_326_545 ();
 FILLCELL_X32 FILLER_326_577 ();
 FILLCELL_X16 FILLER_326_609 ();
 FILLCELL_X4 FILLER_326_625 ();
 FILLCELL_X2 FILLER_326_629 ();
 FILLCELL_X32 FILLER_326_632 ();
 FILLCELL_X32 FILLER_326_664 ();
 FILLCELL_X32 FILLER_326_696 ();
 FILLCELL_X32 FILLER_326_728 ();
 FILLCELL_X32 FILLER_326_760 ();
 FILLCELL_X32 FILLER_326_792 ();
 FILLCELL_X32 FILLER_326_824 ();
 FILLCELL_X32 FILLER_326_856 ();
 FILLCELL_X32 FILLER_326_888 ();
 FILLCELL_X32 FILLER_326_920 ();
 FILLCELL_X32 FILLER_326_952 ();
 FILLCELL_X32 FILLER_326_984 ();
 FILLCELL_X32 FILLER_326_1016 ();
 FILLCELL_X4 FILLER_326_1048 ();
 FILLCELL_X2 FILLER_326_1052 ();
 FILLCELL_X16 FILLER_326_1078 ();
 FILLCELL_X16 FILLER_326_1107 ();
 FILLCELL_X2 FILLER_326_1123 ();
 FILLCELL_X4 FILLER_326_1129 ();
 FILLCELL_X2 FILLER_326_1133 ();
 FILLCELL_X2 FILLER_326_1142 ();
 FILLCELL_X1 FILLER_326_1144 ();
 FILLCELL_X4 FILLER_326_1151 ();
 FILLCELL_X1 FILLER_326_1155 ();
 FILLCELL_X4 FILLER_326_1178 ();
 FILLCELL_X2 FILLER_326_1188 ();
 FILLCELL_X1 FILLER_326_1190 ();
 FILLCELL_X1 FILLER_326_1197 ();
 FILLCELL_X8 FILLER_326_1208 ();
 FILLCELL_X4 FILLER_326_1216 ();
 FILLCELL_X2 FILLER_326_1220 ();
 FILLCELL_X1 FILLER_326_1222 ();
 FILLCELL_X8 FILLER_326_1235 ();
 FILLCELL_X2 FILLER_326_1243 ();
 FILLCELL_X1 FILLER_326_1249 ();
 FILLCELL_X32 FILLER_326_1260 ();
 FILLCELL_X32 FILLER_326_1292 ();
 FILLCELL_X32 FILLER_326_1324 ();
 FILLCELL_X32 FILLER_326_1356 ();
 FILLCELL_X32 FILLER_326_1388 ();
 FILLCELL_X32 FILLER_326_1420 ();
 FILLCELL_X32 FILLER_326_1452 ();
 FILLCELL_X32 FILLER_326_1484 ();
 FILLCELL_X32 FILLER_326_1516 ();
 FILLCELL_X32 FILLER_326_1548 ();
 FILLCELL_X32 FILLER_326_1580 ();
 FILLCELL_X32 FILLER_326_1612 ();
 FILLCELL_X32 FILLER_326_1644 ();
 FILLCELL_X32 FILLER_326_1676 ();
 FILLCELL_X32 FILLER_326_1708 ();
 FILLCELL_X32 FILLER_326_1740 ();
 FILLCELL_X32 FILLER_326_1772 ();
 FILLCELL_X32 FILLER_326_1804 ();
 FILLCELL_X32 FILLER_326_1836 ();
 FILLCELL_X16 FILLER_326_1868 ();
 FILLCELL_X8 FILLER_326_1884 ();
 FILLCELL_X2 FILLER_326_1892 ();
 FILLCELL_X32 FILLER_326_1895 ();
 FILLCELL_X32 FILLER_326_1927 ();
 FILLCELL_X32 FILLER_326_1959 ();
 FILLCELL_X32 FILLER_326_1991 ();
 FILLCELL_X32 FILLER_326_2023 ();
 FILLCELL_X32 FILLER_326_2055 ();
 FILLCELL_X32 FILLER_326_2087 ();
 FILLCELL_X32 FILLER_326_2119 ();
 FILLCELL_X32 FILLER_326_2151 ();
 FILLCELL_X32 FILLER_326_2183 ();
 FILLCELL_X32 FILLER_326_2215 ();
 FILLCELL_X32 FILLER_326_2247 ();
 FILLCELL_X32 FILLER_326_2279 ();
 FILLCELL_X32 FILLER_326_2311 ();
 FILLCELL_X32 FILLER_326_2343 ();
 FILLCELL_X32 FILLER_326_2375 ();
 FILLCELL_X16 FILLER_326_2407 ();
 FILLCELL_X8 FILLER_326_2423 ();
 FILLCELL_X4 FILLER_326_2431 ();
 FILLCELL_X1 FILLER_326_2435 ();
 FILLCELL_X32 FILLER_327_1 ();
 FILLCELL_X32 FILLER_327_33 ();
 FILLCELL_X32 FILLER_327_65 ();
 FILLCELL_X32 FILLER_327_97 ();
 FILLCELL_X32 FILLER_327_129 ();
 FILLCELL_X32 FILLER_327_161 ();
 FILLCELL_X32 FILLER_327_193 ();
 FILLCELL_X32 FILLER_327_225 ();
 FILLCELL_X32 FILLER_327_257 ();
 FILLCELL_X32 FILLER_327_289 ();
 FILLCELL_X32 FILLER_327_321 ();
 FILLCELL_X32 FILLER_327_353 ();
 FILLCELL_X32 FILLER_327_385 ();
 FILLCELL_X32 FILLER_327_417 ();
 FILLCELL_X32 FILLER_327_449 ();
 FILLCELL_X32 FILLER_327_481 ();
 FILLCELL_X32 FILLER_327_513 ();
 FILLCELL_X32 FILLER_327_545 ();
 FILLCELL_X32 FILLER_327_577 ();
 FILLCELL_X32 FILLER_327_609 ();
 FILLCELL_X32 FILLER_327_641 ();
 FILLCELL_X32 FILLER_327_673 ();
 FILLCELL_X32 FILLER_327_705 ();
 FILLCELL_X32 FILLER_327_737 ();
 FILLCELL_X32 FILLER_327_769 ();
 FILLCELL_X32 FILLER_327_801 ();
 FILLCELL_X32 FILLER_327_833 ();
 FILLCELL_X32 FILLER_327_865 ();
 FILLCELL_X32 FILLER_327_897 ();
 FILLCELL_X32 FILLER_327_929 ();
 FILLCELL_X32 FILLER_327_961 ();
 FILLCELL_X32 FILLER_327_993 ();
 FILLCELL_X4 FILLER_327_1025 ();
 FILLCELL_X1 FILLER_327_1029 ();
 FILLCELL_X16 FILLER_327_1044 ();
 FILLCELL_X4 FILLER_327_1060 ();
 FILLCELL_X32 FILLER_327_1068 ();
 FILLCELL_X16 FILLER_327_1100 ();
 FILLCELL_X8 FILLER_327_1116 ();
 FILLCELL_X1 FILLER_327_1138 ();
 FILLCELL_X1 FILLER_327_1145 ();
 FILLCELL_X4 FILLER_327_1160 ();
 FILLCELL_X2 FILLER_327_1166 ();
 FILLCELL_X1 FILLER_327_1168 ();
 FILLCELL_X2 FILLER_327_1173 ();
 FILLCELL_X16 FILLER_327_1187 ();
 FILLCELL_X8 FILLER_327_1203 ();
 FILLCELL_X2 FILLER_327_1233 ();
 FILLCELL_X1 FILLER_327_1235 ();
 FILLCELL_X8 FILLER_327_1239 ();
 FILLCELL_X4 FILLER_327_1247 ();
 FILLCELL_X2 FILLER_327_1251 ();
 FILLCELL_X1 FILLER_327_1253 ();
 FILLCELL_X32 FILLER_327_1286 ();
 FILLCELL_X32 FILLER_327_1318 ();
 FILLCELL_X32 FILLER_327_1350 ();
 FILLCELL_X32 FILLER_327_1382 ();
 FILLCELL_X32 FILLER_327_1414 ();
 FILLCELL_X32 FILLER_327_1446 ();
 FILLCELL_X32 FILLER_327_1478 ();
 FILLCELL_X32 FILLER_327_1510 ();
 FILLCELL_X32 FILLER_327_1542 ();
 FILLCELL_X32 FILLER_327_1574 ();
 FILLCELL_X32 FILLER_327_1606 ();
 FILLCELL_X32 FILLER_327_1638 ();
 FILLCELL_X32 FILLER_327_1670 ();
 FILLCELL_X32 FILLER_327_1702 ();
 FILLCELL_X32 FILLER_327_1734 ();
 FILLCELL_X32 FILLER_327_1766 ();
 FILLCELL_X32 FILLER_327_1798 ();
 FILLCELL_X32 FILLER_327_1830 ();
 FILLCELL_X32 FILLER_327_1862 ();
 FILLCELL_X32 FILLER_327_1894 ();
 FILLCELL_X32 FILLER_327_1926 ();
 FILLCELL_X32 FILLER_327_1958 ();
 FILLCELL_X32 FILLER_327_1990 ();
 FILLCELL_X32 FILLER_327_2022 ();
 FILLCELL_X32 FILLER_327_2054 ();
 FILLCELL_X32 FILLER_327_2086 ();
 FILLCELL_X32 FILLER_327_2118 ();
 FILLCELL_X32 FILLER_327_2150 ();
 FILLCELL_X32 FILLER_327_2182 ();
 FILLCELL_X32 FILLER_327_2214 ();
 FILLCELL_X32 FILLER_327_2246 ();
 FILLCELL_X32 FILLER_327_2278 ();
 FILLCELL_X32 FILLER_327_2310 ();
 FILLCELL_X32 FILLER_327_2342 ();
 FILLCELL_X32 FILLER_327_2374 ();
 FILLCELL_X16 FILLER_327_2406 ();
 FILLCELL_X8 FILLER_327_2422 ();
 FILLCELL_X4 FILLER_327_2430 ();
 FILLCELL_X2 FILLER_327_2434 ();
 FILLCELL_X32 FILLER_328_1 ();
 FILLCELL_X32 FILLER_328_33 ();
 FILLCELL_X32 FILLER_328_65 ();
 FILLCELL_X32 FILLER_328_97 ();
 FILLCELL_X32 FILLER_328_129 ();
 FILLCELL_X32 FILLER_328_161 ();
 FILLCELL_X32 FILLER_328_193 ();
 FILLCELL_X32 FILLER_328_225 ();
 FILLCELL_X32 FILLER_328_257 ();
 FILLCELL_X32 FILLER_328_289 ();
 FILLCELL_X32 FILLER_328_321 ();
 FILLCELL_X32 FILLER_328_353 ();
 FILLCELL_X32 FILLER_328_385 ();
 FILLCELL_X32 FILLER_328_417 ();
 FILLCELL_X32 FILLER_328_449 ();
 FILLCELL_X32 FILLER_328_481 ();
 FILLCELL_X32 FILLER_328_513 ();
 FILLCELL_X32 FILLER_328_545 ();
 FILLCELL_X32 FILLER_328_577 ();
 FILLCELL_X16 FILLER_328_609 ();
 FILLCELL_X4 FILLER_328_625 ();
 FILLCELL_X2 FILLER_328_629 ();
 FILLCELL_X32 FILLER_328_632 ();
 FILLCELL_X32 FILLER_328_664 ();
 FILLCELL_X32 FILLER_328_696 ();
 FILLCELL_X32 FILLER_328_728 ();
 FILLCELL_X32 FILLER_328_760 ();
 FILLCELL_X32 FILLER_328_792 ();
 FILLCELL_X32 FILLER_328_824 ();
 FILLCELL_X32 FILLER_328_856 ();
 FILLCELL_X32 FILLER_328_888 ();
 FILLCELL_X32 FILLER_328_920 ();
 FILLCELL_X32 FILLER_328_952 ();
 FILLCELL_X32 FILLER_328_984 ();
 FILLCELL_X8 FILLER_328_1016 ();
 FILLCELL_X4 FILLER_328_1024 ();
 FILLCELL_X2 FILLER_328_1028 ();
 FILLCELL_X1 FILLER_328_1030 ();
 FILLCELL_X32 FILLER_328_1035 ();
 FILLCELL_X32 FILLER_328_1067 ();
 FILLCELL_X32 FILLER_328_1099 ();
 FILLCELL_X4 FILLER_328_1131 ();
 FILLCELL_X2 FILLER_328_1135 ();
 FILLCELL_X1 FILLER_328_1137 ();
 FILLCELL_X8 FILLER_328_1146 ();
 FILLCELL_X1 FILLER_328_1154 ();
 FILLCELL_X8 FILLER_328_1159 ();
 FILLCELL_X4 FILLER_328_1167 ();
 FILLCELL_X32 FILLER_328_1181 ();
 FILLCELL_X16 FILLER_328_1213 ();
 FILLCELL_X2 FILLER_328_1229 ();
 FILLCELL_X32 FILLER_328_1253 ();
 FILLCELL_X32 FILLER_328_1285 ();
 FILLCELL_X32 FILLER_328_1317 ();
 FILLCELL_X32 FILLER_328_1349 ();
 FILLCELL_X32 FILLER_328_1381 ();
 FILLCELL_X32 FILLER_328_1413 ();
 FILLCELL_X32 FILLER_328_1445 ();
 FILLCELL_X32 FILLER_328_1477 ();
 FILLCELL_X32 FILLER_328_1509 ();
 FILLCELL_X32 FILLER_328_1541 ();
 FILLCELL_X32 FILLER_328_1573 ();
 FILLCELL_X32 FILLER_328_1605 ();
 FILLCELL_X32 FILLER_328_1637 ();
 FILLCELL_X32 FILLER_328_1669 ();
 FILLCELL_X32 FILLER_328_1701 ();
 FILLCELL_X32 FILLER_328_1733 ();
 FILLCELL_X32 FILLER_328_1765 ();
 FILLCELL_X32 FILLER_328_1797 ();
 FILLCELL_X32 FILLER_328_1829 ();
 FILLCELL_X32 FILLER_328_1861 ();
 FILLCELL_X1 FILLER_328_1893 ();
 FILLCELL_X32 FILLER_328_1895 ();
 FILLCELL_X32 FILLER_328_1927 ();
 FILLCELL_X32 FILLER_328_1959 ();
 FILLCELL_X32 FILLER_328_1991 ();
 FILLCELL_X32 FILLER_328_2023 ();
 FILLCELL_X32 FILLER_328_2055 ();
 FILLCELL_X32 FILLER_328_2087 ();
 FILLCELL_X32 FILLER_328_2119 ();
 FILLCELL_X32 FILLER_328_2151 ();
 FILLCELL_X32 FILLER_328_2183 ();
 FILLCELL_X32 FILLER_328_2215 ();
 FILLCELL_X32 FILLER_328_2247 ();
 FILLCELL_X32 FILLER_328_2279 ();
 FILLCELL_X32 FILLER_328_2311 ();
 FILLCELL_X32 FILLER_328_2343 ();
 FILLCELL_X32 FILLER_328_2375 ();
 FILLCELL_X16 FILLER_328_2407 ();
 FILLCELL_X8 FILLER_328_2423 ();
 FILLCELL_X4 FILLER_328_2431 ();
 FILLCELL_X1 FILLER_328_2435 ();
 FILLCELL_X32 FILLER_329_1 ();
 FILLCELL_X32 FILLER_329_33 ();
 FILLCELL_X32 FILLER_329_65 ();
 FILLCELL_X32 FILLER_329_97 ();
 FILLCELL_X32 FILLER_329_129 ();
 FILLCELL_X32 FILLER_329_161 ();
 FILLCELL_X32 FILLER_329_193 ();
 FILLCELL_X32 FILLER_329_225 ();
 FILLCELL_X32 FILLER_329_257 ();
 FILLCELL_X32 FILLER_329_289 ();
 FILLCELL_X32 FILLER_329_321 ();
 FILLCELL_X32 FILLER_329_353 ();
 FILLCELL_X32 FILLER_329_385 ();
 FILLCELL_X32 FILLER_329_417 ();
 FILLCELL_X32 FILLER_329_449 ();
 FILLCELL_X32 FILLER_329_481 ();
 FILLCELL_X32 FILLER_329_513 ();
 FILLCELL_X32 FILLER_329_545 ();
 FILLCELL_X32 FILLER_329_577 ();
 FILLCELL_X16 FILLER_329_609 ();
 FILLCELL_X4 FILLER_329_625 ();
 FILLCELL_X2 FILLER_329_629 ();
 FILLCELL_X32 FILLER_329_632 ();
 FILLCELL_X32 FILLER_329_664 ();
 FILLCELL_X32 FILLER_329_696 ();
 FILLCELL_X32 FILLER_329_728 ();
 FILLCELL_X32 FILLER_329_760 ();
 FILLCELL_X32 FILLER_329_792 ();
 FILLCELL_X32 FILLER_329_824 ();
 FILLCELL_X32 FILLER_329_856 ();
 FILLCELL_X32 FILLER_329_888 ();
 FILLCELL_X32 FILLER_329_920 ();
 FILLCELL_X32 FILLER_329_952 ();
 FILLCELL_X16 FILLER_329_984 ();
 FILLCELL_X8 FILLER_329_1000 ();
 FILLCELL_X4 FILLER_329_1008 ();
 FILLCELL_X1 FILLER_329_1012 ();
 FILLCELL_X16 FILLER_329_1033 ();
 FILLCELL_X1 FILLER_329_1049 ();
 FILLCELL_X32 FILLER_329_1063 ();
 FILLCELL_X1 FILLER_329_1095 ();
 FILLCELL_X2 FILLER_329_1100 ();
 FILLCELL_X16 FILLER_329_1106 ();
 FILLCELL_X4 FILLER_329_1122 ();
 FILLCELL_X2 FILLER_329_1126 ();
 FILLCELL_X1 FILLER_329_1128 ();
 FILLCELL_X8 FILLER_329_1132 ();
 FILLCELL_X1 FILLER_329_1140 ();
 FILLCELL_X8 FILLER_329_1144 ();
 FILLCELL_X1 FILLER_329_1152 ();
 FILLCELL_X32 FILLER_329_1164 ();
 FILLCELL_X32 FILLER_329_1196 ();
 FILLCELL_X16 FILLER_329_1228 ();
 FILLCELL_X2 FILLER_329_1244 ();
 FILLCELL_X1 FILLER_329_1246 ();
 FILLCELL_X4 FILLER_329_1257 ();
 FILLCELL_X1 FILLER_329_1261 ();
 FILLCELL_X32 FILLER_329_1263 ();
 FILLCELL_X32 FILLER_329_1295 ();
 FILLCELL_X32 FILLER_329_1327 ();
 FILLCELL_X32 FILLER_329_1359 ();
 FILLCELL_X32 FILLER_329_1391 ();
 FILLCELL_X32 FILLER_329_1423 ();
 FILLCELL_X32 FILLER_329_1455 ();
 FILLCELL_X32 FILLER_329_1487 ();
 FILLCELL_X32 FILLER_329_1519 ();
 FILLCELL_X32 FILLER_329_1551 ();
 FILLCELL_X32 FILLER_329_1583 ();
 FILLCELL_X32 FILLER_329_1615 ();
 FILLCELL_X32 FILLER_329_1647 ();
 FILLCELL_X32 FILLER_329_1679 ();
 FILLCELL_X32 FILLER_329_1711 ();
 FILLCELL_X32 FILLER_329_1743 ();
 FILLCELL_X32 FILLER_329_1775 ();
 FILLCELL_X32 FILLER_329_1807 ();
 FILLCELL_X32 FILLER_329_1839 ();
 FILLCELL_X16 FILLER_329_1871 ();
 FILLCELL_X4 FILLER_329_1887 ();
 FILLCELL_X2 FILLER_329_1891 ();
 FILLCELL_X32 FILLER_329_1894 ();
 FILLCELL_X32 FILLER_329_1926 ();
 FILLCELL_X32 FILLER_329_1958 ();
 FILLCELL_X32 FILLER_329_1990 ();
 FILLCELL_X32 FILLER_329_2022 ();
 FILLCELL_X32 FILLER_329_2054 ();
 FILLCELL_X32 FILLER_329_2086 ();
 FILLCELL_X32 FILLER_329_2118 ();
 FILLCELL_X32 FILLER_329_2150 ();
 FILLCELL_X32 FILLER_329_2182 ();
 FILLCELL_X32 FILLER_329_2214 ();
 FILLCELL_X32 FILLER_329_2246 ();
 FILLCELL_X32 FILLER_329_2278 ();
 FILLCELL_X32 FILLER_329_2310 ();
 FILLCELL_X32 FILLER_329_2342 ();
 FILLCELL_X32 FILLER_329_2374 ();
 FILLCELL_X16 FILLER_329_2406 ();
 FILLCELL_X8 FILLER_329_2422 ();
 FILLCELL_X4 FILLER_329_2430 ();
 FILLCELL_X2 FILLER_329_2434 ();
endmodule
