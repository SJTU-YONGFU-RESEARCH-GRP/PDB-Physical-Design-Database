module hamming_code (single_bit_error,
    corrected_code,
    data_in,
    data_out,
    encoded_out,
    received_in);
 output single_bit_error;
 output [6:0] corrected_code;
 input [3:0] data_in;
 output [3:0] data_out;
 output [6:0] encoded_out;
 input [6:0] received_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire p1;
 wire p2;
 wire p3;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;

 sky130_fd_sc_hd__buf_4 _080_ (.A(received_in[2]),
    .X(_009_));
 sky130_fd_sc_hd__xnor2_2 _081_ (.A(_009_),
    .B(net5),
    .Y(_010_));
 sky130_fd_sc_hd__buf_6 _082_ (.A(_010_),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_2 _083_ (.A(received_in[5]),
    .X(_012_));
 sky130_fd_sc_hd__xor2_1 _084_ (.A(_012_),
    .B(net7),
    .X(_013_));
 sky130_fd_sc_hd__xor2_1 _085_ (.A(net8),
    .B(net9),
    .X(_014_));
 sky130_fd_sc_hd__or2_0 _086_ (.A(_013_),
    .B(_014_),
    .X(_015_));
 sky130_fd_sc_hd__nand3_1 _087_ (.A(_013_),
    .B(_014_),
    .C(_011_),
    .Y(_016_));
 sky130_fd_sc_hd__o21ai_1 _088_ (.A1(_011_),
    .A2(_015_),
    .B1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__xnor2_1 _089_ (.A(_009_),
    .B(net6),
    .Y(_018_));
 sky130_fd_sc_hd__buf_2 _090_ (.A(_018_),
    .X(_019_));
 sky130_fd_sc_hd__xnor2_2 _091_ (.A(net9),
    .B(_012_),
    .Y(_020_));
 sky130_fd_sc_hd__xnor2_1 _092_ (.A(_019_),
    .B(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _093_ (.A(_017_),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__xnor2_1 _094_ (.A(net5),
    .B(_022_),
    .Y(net10));
 sky130_fd_sc_hd__xnor2_1 _095_ (.A(_009_),
    .B(_020_),
    .Y(_023_));
 sky130_fd_sc_hd__xor2_1 _096_ (.A(_009_),
    .B(net5),
    .X(_024_));
 sky130_fd_sc_hd__buf_4 _097_ (.A(_024_),
    .X(_025_));
 sky130_fd_sc_hd__nand3_1 _098_ (.A(_013_),
    .B(_014_),
    .C(_024_),
    .Y(_026_));
 sky130_fd_sc_hd__o21ai_1 _099_ (.A1(_025_),
    .A2(_015_),
    .B1(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__mux2_1 _100_ (.A0(net6),
    .A1(_023_),
    .S(_027_),
    .X(net11));
 sky130_fd_sc_hd__xnor2_1 _101_ (.A(net6),
    .B(_020_),
    .Y(_028_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(_009_),
    .A1(_028_),
    .S(_017_),
    .X(net12));
 sky130_fd_sc_hd__buf_2 _103_ (.A(net7),
    .X(_029_));
 sky130_fd_sc_hd__nor2_1 _104_ (.A(_029_),
    .B(_010_),
    .Y(_030_));
 sky130_fd_sc_hd__buf_2 _105_ (.A(net7),
    .X(_031_));
 sky130_fd_sc_hd__xor2_4 _106_ (.A(_009_),
    .B(net6),
    .X(_032_));
 sky130_fd_sc_hd__nand2_1 _107_ (.A(_010_),
    .B(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__buf_2 _108_ (.A(_012_),
    .X(_034_));
 sky130_fd_sc_hd__a21oi_1 _109_ (.A1(_031_),
    .A2(_033_),
    .B1(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__buf_2 _110_ (.A(net9),
    .X(_036_));
 sky130_fd_sc_hd__o21a_1 _111_ (.A1(_030_),
    .A2(_035_),
    .B1(_036_),
    .X(_037_));
 sky130_fd_sc_hd__inv_1 _112_ (.A(_012_),
    .Y(_038_));
 sky130_fd_sc_hd__nand2_1 _113_ (.A(_038_),
    .B(_025_),
    .Y(_039_));
 sky130_fd_sc_hd__o21ai_0 _114_ (.A1(_011_),
    .A2(_019_),
    .B1(_029_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _115_ (.A(_039_),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__buf_2 _116_ (.A(net8),
    .X(_042_));
 sky130_fd_sc_hd__o221ai_1 _117_ (.A1(_031_),
    .A2(_019_),
    .B1(_041_),
    .B2(_036_),
    .C1(_042_),
    .Y(_043_));
 sky130_fd_sc_hd__o21ai_0 _118_ (.A1(_025_),
    .A2(_032_),
    .B1(_031_),
    .Y(_044_));
 sky130_fd_sc_hd__a21oi_1 _119_ (.A1(_038_),
    .A2(_044_),
    .B1(_030_),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_0 _120_ (.A1(_011_),
    .A2(_032_),
    .B1(_031_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_1 _121_ (.A(_042_),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_0 _122_ (.A1(_031_),
    .A2(_032_),
    .B1(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__a31oi_1 _123_ (.A1(_036_),
    .A2(_046_),
    .A3(_039_),
    .B1(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__o21ai_0 _124_ (.A1(_036_),
    .A2(_045_),
    .B1(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__o21ai_0 _125_ (.A1(_037_),
    .A2(_043_),
    .B1(_050_),
    .Y(net13));
 sky130_fd_sc_hd__a21oi_1 _126_ (.A1(_029_),
    .A2(_019_),
    .B1(_042_),
    .Y(_051_));
 sky130_fd_sc_hd__nor3_1 _127_ (.A(_029_),
    .B(_024_),
    .C(_032_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _128_ (.A(_051_),
    .B(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__o22ai_1 _129_ (.A1(_042_),
    .A2(_025_),
    .B1(_053_),
    .B2(_034_),
    .Y(_054_));
 sky130_fd_sc_hd__o21ai_0 _130_ (.A1(_029_),
    .A2(_019_),
    .B1(_047_),
    .Y(_055_));
 sky130_fd_sc_hd__nand3_1 _131_ (.A(_031_),
    .B(_011_),
    .C(_032_),
    .Y(_056_));
 sky130_fd_sc_hd__a21oi_1 _132_ (.A1(_055_),
    .A2(_056_),
    .B1(_038_),
    .Y(_057_));
 sky130_fd_sc_hd__nor3_1 _133_ (.A(_031_),
    .B(_011_),
    .C(_032_),
    .Y(_058_));
 sky130_fd_sc_hd__o21ai_0 _134_ (.A1(_051_),
    .A2(_058_),
    .B1(_034_),
    .Y(_059_));
 sky130_fd_sc_hd__nand3_1 _135_ (.A(_029_),
    .B(_025_),
    .C(_032_),
    .Y(_060_));
 sky130_fd_sc_hd__a21o_1 _136_ (.A1(_055_),
    .A2(_060_),
    .B1(_034_),
    .X(_061_));
 sky130_fd_sc_hd__o2111ai_1 _137_ (.A1(_042_),
    .A2(_011_),
    .B1(_059_),
    .C1(_061_),
    .D1(_036_),
    .Y(_062_));
 sky130_fd_sc_hd__o31ai_2 _138_ (.A1(_036_),
    .A2(_054_),
    .A3(_057_),
    .B1(_062_),
    .Y(net14));
 sky130_fd_sc_hd__a21oi_1 _139_ (.A1(_029_),
    .A2(_011_),
    .B1(_012_),
    .Y(_063_));
 sky130_fd_sc_hd__o21ai_0 _140_ (.A1(_052_),
    .A2(_063_),
    .B1(_047_),
    .Y(_064_));
 sky130_fd_sc_hd__o21ai_0 _141_ (.A1(_034_),
    .A2(_032_),
    .B1(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__nand4_1 _142_ (.A(_042_),
    .B(_031_),
    .C(_025_),
    .D(_019_),
    .Y(_066_));
 sky130_fd_sc_hd__inv_1 _143_ (.A(_036_),
    .Y(_067_));
 sky130_fd_sc_hd__o311ai_1 _144_ (.A1(_047_),
    .A2(_034_),
    .A3(_030_),
    .B1(_066_),
    .C1(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__o21a_1 _145_ (.A1(_034_),
    .A2(_030_),
    .B1(_060_),
    .X(_069_));
 sky130_fd_sc_hd__nor3_1 _146_ (.A(_029_),
    .B(_025_),
    .C(_019_),
    .Y(_070_));
 sky130_fd_sc_hd__o21ai_0 _147_ (.A1(_063_),
    .A2(_070_),
    .B1(_042_),
    .Y(_071_));
 sky130_fd_sc_hd__o221ai_1 _148_ (.A1(_034_),
    .A2(_019_),
    .B1(_069_),
    .B2(_042_),
    .C1(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__o22ai_2 _149_ (.A1(_065_),
    .A2(_068_),
    .B1(_072_),
    .B2(_067_),
    .Y(net15));
 sky130_fd_sc_hd__xnor2_1 _150_ (.A(_034_),
    .B(_019_),
    .Y(_073_));
 sky130_fd_sc_hd__nand2_1 _151_ (.A(net9),
    .B(_033_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_1 _152_ (.A(_012_),
    .B(net7),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _153_ (.A(_011_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__nor2_1 _154_ (.A(net9),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__and3_1 _155_ (.A(_011_),
    .B(_018_),
    .C(_075_),
    .X(_078_));
 sky130_fd_sc_hd__a311oi_1 _156_ (.A1(_034_),
    .A2(_031_),
    .A3(_074_),
    .B1(_077_),
    .C1(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _157_ (.A(_038_),
    .B(_029_),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _158_ (.A(_025_),
    .B(_019_),
    .Y(_001_));
 sky130_fd_sc_hd__a21oi_1 _159_ (.A1(_038_),
    .A2(_029_),
    .B1(_025_),
    .Y(_002_));
 sky130_fd_sc_hd__o22ai_1 _160_ (.A1(_000_),
    .A2(_001_),
    .B1(_002_),
    .B2(_036_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _161_ (.A(_025_),
    .B(_032_),
    .Y(_004_));
 sky130_fd_sc_hd__a211oi_1 _162_ (.A1(_036_),
    .A2(_004_),
    .B1(_031_),
    .C1(_038_),
    .Y(_005_));
 sky130_fd_sc_hd__o21ai_0 _163_ (.A1(_003_),
    .A2(_005_),
    .B1(_042_),
    .Y(_006_));
 sky130_fd_sc_hd__o221a_1 _164_ (.A1(_036_),
    .A2(_073_),
    .B1(_079_),
    .B2(_042_),
    .C1(_006_),
    .X(net16));
 sky130_fd_sc_hd__xnor2_1 _165_ (.A(net4),
    .B(net2),
    .Y(_007_));
 sky130_fd_sc_hd__xnor2_1 _166_ (.A(net1),
    .B(_007_),
    .Y(p1));
 sky130_fd_sc_hd__xnor2_1 _167_ (.A(net1),
    .B(net3),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_1 _168_ (.A(net4),
    .B(_008_),
    .Y(p2));
 sky130_fd_sc_hd__xnor2_1 _169_ (.A(net3),
    .B(_007_),
    .Y(p3));
 sky130_fd_sc_hd__nand2_1 _170_ (.A(_021_),
    .B(_027_),
    .Y(net28));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(net12),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(net14),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(net15),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 _174_ (.A(net16),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 _175_ (.A(p1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 _176_ (.A(p2),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 _177_ (.A(net1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _178_ (.A(p3),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _179_ (.A(net2),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _180_ (.A(net3),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 _181_ (.A(net4),
    .X(net27));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_51 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(data_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(received_in[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(received_in[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(received_in[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(received_in[4]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(received_in[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(corrected_code[0]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(corrected_code[1]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(corrected_code[2]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(corrected_code[3]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(corrected_code[4]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(corrected_code[5]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(corrected_code[6]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(encoded_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(encoded_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(encoded_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(encoded_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(encoded_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(encoded_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(encoded_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(single_bit_error));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_13 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_145 ();
endmodule
