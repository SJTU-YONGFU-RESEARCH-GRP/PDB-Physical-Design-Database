module non_restoring_divider (busy,
    clk,
    error,
    rst_n,
    start,
    valid,
    dividend,
    divisor,
    quotient,
    remainder);
 output busy;
 input clk;
 output error;
 input rst_n;
 input start;
 output valid;
 input [7:0] dividend;
 input [7:0] divisor;
 output [7:0] quotient;
 output [7:0] remainder;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire \div_reg[0] ;
 wire \div_reg[1] ;
 wire \div_reg[2] ;
 wire \div_reg[3] ;
 wire \div_reg[4] ;
 wire \div_reg[5] ;
 wire \div_reg[6] ;
 wire \div_reg[7] ;
 wire \iter[0] ;
 wire \iter[1] ;
 wire \iter[2] ;
 wire \iter[3] ;
 wire \quot[0] ;
 wire \quot[1] ;
 wire \quot[2] ;
 wire \quot[3] ;
 wire \quot[4] ;
 wire \quot[5] ;
 wire \quot[6] ;
 wire \quot[7] ;
 wire \rem[0] ;
 wire \rem[1] ;
 wire \rem[2] ;
 wire \rem[3] ;
 wire \rem[4] ;
 wire \rem[5] ;
 wire \rem[6] ;
 wire \rem[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net38;

 gf180mcu_fd_sc_mcu9t5v0__inv_2 _220_ (.I(\iter[3] ),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _221_ (.I(\iter[2] ),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _222_ (.I(_174_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _223_ (.I0(net5),
    .I1(net4),
    .I2(net3),
    .I3(net2),
    .S0(\iter[0] ),
    .S1(_173_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _224_ (.A1(\iter[0] ),
    .A2(\iter[1] ),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _225_ (.A1(_050_),
    .A2(_051_),
    .A3(_052_),
    .A4(_053_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _226_ (.A1(\iter[2] ),
    .A2(_174_),
    .A3(_052_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _227_ (.I0(net9),
    .I1(net8),
    .I2(net7),
    .I3(net6),
    .S0(\iter[0] ),
    .S1(_173_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _228_ (.A1(\iter[2] ),
    .A2(_051_),
    .A3(_056_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _229_ (.A1(_054_),
    .A2(_055_),
    .A3(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _230_ (.I(\iter[0] ),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _231_ (.I(\iter[1] ),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _232_ (.A1(_170_),
    .A2(_171_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _233_ (.I0(_052_),
    .I1(_056_),
    .S(_174_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _234_ (.A1(_050_),
    .A2(\iter[3] ),
    .A3(_059_),
    .A4(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _235_ (.A1(_049_),
    .A2(_058_),
    .B(_061_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _236_ (.I(_180_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _237_ (.I(\div_reg[0] ),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _238_ (.I(\div_reg[1] ),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _239_ (.I(\div_reg[3] ),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _240_ (.I(\div_reg[2] ),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _241_ (.I(\div_reg[6] ),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _242_ (.I(\div_reg[5] ),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _243_ (.I(\div_reg[4] ),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _244_ (.I(\rem[0] ),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _245_ (.I(\rem[2] ),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _246_ (.I(\rem[1] ),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _247_ (.I(\rem[6] ),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _248_ (.I(\rem[5] ),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _249_ (.I(\rem[4] ),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _250_ (.I(\rem[3] ),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _251_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _252_ (.A1(net18),
    .A2(_062_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _253_ (.A1(net15),
    .A2(net14),
    .A3(net17),
    .A4(net16),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _254_ (.A1(net11),
    .A2(net10),
    .A3(net13),
    .A4(net12),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _255_ (.A1(_064_),
    .A2(_065_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _256_ (.A1(_063_),
    .A2(_066_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _257_ (.I(\state[1] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _258_ (.A1(_068_),
    .A2(\state[0] ),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _259_ (.A1(_050_),
    .A2(_049_),
    .A3(_172_),
    .A4(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _260_ (.I(_070_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _261_ (.A1(\state[1] ),
    .A2(\state[0] ),
    .B(net19),
    .C(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _262_ (.A1(_067_),
    .A2(_072_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _263_ (.I0(net10),
    .I1(\div_reg[0] ),
    .S(_067_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _264_ (.I0(net11),
    .I1(\div_reg[1] ),
    .S(_067_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _265_ (.I0(net12),
    .I1(\div_reg[2] ),
    .S(_067_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _266_ (.I0(net13),
    .I1(\div_reg[3] ),
    .S(_067_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _267_ (.I0(net14),
    .I1(\div_reg[4] ),
    .S(_067_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _268_ (.I0(net15),
    .I1(\div_reg[5] ),
    .S(_067_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _269_ (.I0(net16),
    .I1(\div_reg[6] ),
    .S(_067_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _270_ (.I0(net17),
    .I1(\div_reg[7] ),
    .S(_067_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _271_ (.I(net20),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _272_ (.A1(net18),
    .A2(_062_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _273_ (.A1(_073_),
    .A2(_062_),
    .B1(_074_),
    .B2(_066_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _274_ (.I(_172_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _275_ (.A1(\iter[2] ),
    .A2(\iter[3] ),
    .A3(_075_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _276_ (.A1(_069_),
    .A2(_076_),
    .Z(_077_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _277_ (.I(_077_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _278_ (.A1(_063_),
    .A2(_066_),
    .B1(_069_),
    .B2(_076_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _279_ (.I(_079_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _280_ (.I0(_078_),
    .I1(_080_),
    .S(\iter[0] ),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _281_ (.A1(_069_),
    .A2(_076_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _282_ (.I(_081_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _283_ (.I(_079_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _284_ (.I(_083_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _285_ (.A1(_173_),
    .A2(_082_),
    .B1(_046_),
    .B2(_171_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _286_ (.A1(_174_),
    .A2(_082_),
    .B(_083_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _287_ (.A1(_174_),
    .A2(_078_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _288_ (.I0(_084_),
    .I1(_085_),
    .S(_050_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _289_ (.I(\state[0] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _290_ (.A1(_075_),
    .A2(_053_),
    .B(\iter[2] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _291_ (.A1(\state[1] ),
    .A2(_086_),
    .A3(_087_),
    .B(_046_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _292_ (.A1(_050_),
    .A2(\iter[3] ),
    .A3(_059_),
    .A4(_069_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _293_ (.A1(_049_),
    .A2(_088_),
    .B(_089_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _294_ (.A1(_201_),
    .A2(_204_),
    .A3(_210_),
    .A4(_216_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _295_ (.A1(_189_),
    .A2(_195_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _296_ (.A1(_184_),
    .A2(_179_),
    .A3(_090_),
    .A4(_091_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _297_ (.A1(_201_),
    .A2(_204_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _298_ (.A1(_218_),
    .A2(_210_),
    .B(_212_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _299_ (.A1(_206_),
    .A2(_201_),
    .B(_200_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _300_ (.A1(_093_),
    .A2(_094_),
    .B(_095_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _301_ (.A1(_189_),
    .A2(_195_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _302_ (.I(_178_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _303_ (.A1(_184_),
    .A2(_098_),
    .B(_185_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _304_ (.A1(_197_),
    .A2(_189_),
    .B(_191_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _305_ (.A1(_097_),
    .A2(_099_),
    .B(_100_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _306_ (.A1(_090_),
    .A2(_092_),
    .Z(_102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_4 _307_ (.A1(_092_),
    .A2(_096_),
    .B1(_101_),
    .B2(_102_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _308_ (.A1(_078_),
    .A2(_103_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _309_ (.A1(\quot[0] ),
    .A2(_080_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _310_ (.A1(_104_),
    .A2(_105_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _311_ (.A1(\quot[0] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[1] ),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _312_ (.I(_106_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _313_ (.A1(\quot[1] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[2] ),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _314_ (.I(_107_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _315_ (.A1(\quot[2] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[3] ),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _316_ (.I(_108_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _317_ (.A1(\quot[3] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[4] ),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _318_ (.I(_109_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _319_ (.A1(\quot[4] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[5] ),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _320_ (.I(_110_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _321_ (.A1(\quot[5] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[6] ),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _322_ (.I(_111_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _323_ (.A1(\quot[6] ),
    .A2(_078_),
    .B1(_080_),
    .B2(\quot[7] ),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _324_ (.I(_112_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _325_ (.I0(\quot[0] ),
    .I1(net21),
    .S(_071_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _326_ (.I0(\quot[1] ),
    .I1(net22),
    .S(_071_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _327_ (.I0(\quot[2] ),
    .I1(net23),
    .S(_071_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _328_ (.I0(\quot[3] ),
    .I1(net24),
    .S(_071_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _329_ (.I0(\quot[4] ),
    .I1(net25),
    .S(_071_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _330_ (.I0(\quot[5] ),
    .I1(net26),
    .S(_071_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _331_ (.I0(\quot[6] ),
    .I1(net27),
    .S(_071_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _332_ (.I0(\quot[7] ),
    .I1(net28),
    .S(_070_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _333_ (.I(_184_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _334_ (.I(_185_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _335_ (.A1(_113_),
    .A2(_178_),
    .B(_114_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _336_ (.A1(_197_),
    .A2(_189_),
    .B1(_091_),
    .B2(_115_),
    .C(_191_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _337_ (.A1(_090_),
    .A2(_092_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _338_ (.A1(_092_),
    .A2(_096_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _339_ (.A1(_116_),
    .A2(_117_),
    .B(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _340_ (.I0(_179_),
    .I1(_180_),
    .S(_119_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _341_ (.A1(_166_),
    .A2(_046_),
    .B1(_120_),
    .B2(_082_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _342_ (.I(_169_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _343_ (.I0(_121_),
    .I1(_166_),
    .S(_119_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _344_ (.A1(_196_),
    .A2(_046_),
    .B1(_122_),
    .B2(_082_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _345_ (.A1(_168_),
    .A2(_195_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _346_ (.I0(_196_),
    .I1(_123_),
    .S(_103_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _347_ (.A1(_190_),
    .A2(_046_),
    .B1(_124_),
    .B2(_082_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _348_ (.I(_189_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _349_ (.I(_183_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _350_ (.A1(_113_),
    .A2(_167_),
    .B(_126_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _351_ (.A1(_195_),
    .A2(_127_),
    .B(_194_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _352_ (.A1(_125_),
    .A2(_128_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _353_ (.I0(_190_),
    .I1(_129_),
    .S(_103_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _354_ (.A1(_217_),
    .A2(_046_),
    .B1(_130_),
    .B2(_082_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _355_ (.I(_168_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _356_ (.A1(_131_),
    .A2(_195_),
    .B(_194_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _357_ (.I(_188_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _358_ (.A1(_125_),
    .A2(_132_),
    .B(_133_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _359_ (.A1(_216_),
    .A2(_134_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _360_ (.I0(_217_),
    .I1(_135_),
    .S(_103_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _361_ (.A1(_211_),
    .A2(_046_),
    .B1(_136_),
    .B2(_082_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _362_ (.I(_210_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _363_ (.I(_167_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _364_ (.A1(_184_),
    .A2(_138_),
    .B(_183_),
    .C(_194_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _365_ (.A1(_195_),
    .A2(_194_),
    .B(_189_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _366_ (.A1(_139_),
    .A2(_140_),
    .B(_133_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _367_ (.A1(_216_),
    .A2(_141_),
    .B(_215_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _368_ (.A1(_137_),
    .A2(_142_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _369_ (.A1(_211_),
    .A2(_082_),
    .A3(_103_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _370_ (.A1(_205_),
    .A2(_046_),
    .B1(_104_),
    .B2(_143_),
    .C(_144_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _371_ (.A1(_131_),
    .A2(_195_),
    .B(_188_),
    .C(_194_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _372_ (.A1(_189_),
    .A2(_188_),
    .B(_216_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _373_ (.I(_215_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _374_ (.A1(_145_),
    .A2(_146_),
    .B(_147_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _375_ (.A1(_210_),
    .A2(_148_),
    .B(_209_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _376_ (.A1(_204_),
    .A2(_149_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _377_ (.A1(_205_),
    .A2(_082_),
    .A3(_103_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _378_ (.A1(_199_),
    .A2(_046_),
    .B1(_104_),
    .B2(_150_),
    .C(_151_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _379_ (.I(_203_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _380_ (.A1(_216_),
    .A2(_188_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _381_ (.A1(_147_),
    .A2(_153_),
    .B(_137_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _382_ (.A1(_210_),
    .A2(_216_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _383_ (.A1(_155_),
    .A2(_139_),
    .A3(_140_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _384_ (.A1(_209_),
    .A2(_154_),
    .A3(_156_),
    .B(_204_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _385_ (.A1(_201_),
    .A2(_081_),
    .Z(_158_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _386_ (.A1(_152_),
    .A2(_157_),
    .B(_158_),
    .C(_119_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _387_ (.A1(_201_),
    .A2(_077_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _388_ (.A1(_152_),
    .A2(_103_),
    .A3(_157_),
    .A4(_160_),
    .Z(_161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _389_ (.A1(\rem[7] ),
    .A2(_080_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _390_ (.A1(_199_),
    .A2(_082_),
    .A3(_103_),
    .B(_162_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _391_ (.A1(_159_),
    .A2(_161_),
    .A3(_163_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _392_ (.I0(\rem[0] ),
    .I1(net29),
    .S(_070_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _393_ (.I0(\rem[1] ),
    .I1(net30),
    .S(_070_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _394_ (.I0(\rem[2] ),
    .I1(net31),
    .S(_070_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _395_ (.I0(\rem[3] ),
    .I1(net32),
    .S(_070_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _396_ (.I0(\rem[4] ),
    .I1(net33),
    .S(_070_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _397_ (.I0(\rem[5] ),
    .I1(net34),
    .S(_070_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _398_ (.I0(\rem[6] ),
    .I1(net35),
    .S(_070_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _399_ (.I0(\rem[7] ),
    .I1(net36),
    .S(_070_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _400_ (.A1(net18),
    .A2(_068_),
    .A3(\state[0] ),
    .B(_071_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _401_ (.A1(net18),
    .A2(_068_),
    .B(_086_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _402_ (.A1(net37),
    .A2(_164_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _403_ (.A1(_071_),
    .A2(_165_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _404_ (.A(\div_reg[1] ),
    .B(_166_),
    .CI(_167_),
    .CO(_168_),
    .S(_169_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _405_ (.A(_170_),
    .B(_171_),
    .CO(_172_),
    .S(_173_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _406_ (.A(_170_),
    .B(_171_),
    .CO(_174_),
    .S(_175_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _407_ (.A(_176_),
    .B(_177_),
    .CO(_178_),
    .S(_179_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _408_ (.A(\div_reg[0] ),
    .B(_180_),
    .CO(_167_),
    .S(_181_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _409_ (.A(_182_),
    .B(\rem[0] ),
    .CO(_183_),
    .S(_184_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _410_ (.A(\div_reg[1] ),
    .B(_166_),
    .CO(_185_),
    .S(_186_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _411_ (.A(_187_),
    .B(\rem[2] ),
    .CO(_188_),
    .S(_189_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _412_ (.A(\div_reg[3] ),
    .B(_190_),
    .CO(_191_),
    .S(_192_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _413_ (.A(_193_),
    .B(\rem[1] ),
    .CO(_194_),
    .S(_195_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _414_ (.A(\div_reg[2] ),
    .B(_196_),
    .CO(_197_),
    .S(_198_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _415_ (.A(\div_reg[7] ),
    .B(_199_),
    .CO(_200_),
    .S(_201_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _416_ (.A(_202_),
    .B(\rem[5] ),
    .CO(_203_),
    .S(_204_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _417_ (.A(\div_reg[6] ),
    .B(_205_),
    .CO(_206_),
    .S(_207_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _418_ (.A(_208_),
    .B(\rem[4] ),
    .CO(_209_),
    .S(_210_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _419_ (.A(\div_reg[5] ),
    .B(_211_),
    .CO(_212_),
    .S(_213_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _420_ (.A(_214_),
    .B(\rem[3] ),
    .CO(_215_),
    .S(_216_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _421_ (.A(\div_reg[4] ),
    .B(_217_),
    .CO(_218_),
    .S(_219_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \busy$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\div_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\div_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\div_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[3]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\div_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[4]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\div_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[5]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\div_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[6]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\div_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \div_reg[7]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\div_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \error$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \iter[0]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\iter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \iter[1]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\iter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \iter[2]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\iter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \iter[3]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\iter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[0]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\quot[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[1]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\quot[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[2]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\quot[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[3]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\quot[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[4]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\quot[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[5]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\quot[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[6]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\quot[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quot[7]$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\quot[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[0]$_DFFE_PN0P_  (.D(_022_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[1]$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[2]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[3]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[4]$_DFFE_PN0P_  (.D(_026_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[5]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[6]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \quotient[7]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[0]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rem[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[1]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rem[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[2]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rem[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[3]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rem[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[4]$_DFFE_PN0P_  (.D(_034_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rem[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[5]$_DFFE_PN0P_  (.D(_035_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rem[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[6]$_DFFE_PN0P_  (.D(_036_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rem[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rem[7]$_DFFE_PN0P_  (.D(_037_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rem[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[0]$_DFFE_PN0P_  (.D(_038_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[1]$_DFFE_PN0P_  (.D(_039_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[2]$_DFFE_PN0P_  (.D(_040_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[3]$_DFFE_PN0P_  (.D(_041_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[4]$_DFFE_PN0P_  (.D(_042_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[5]$_DFFE_PN0P_  (.D(_043_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net34));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[6]$_DFFE_PN0P_  (.D(_044_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net35));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \remainder[7]$_DFFE_PN0P_  (.D(_045_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net36));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[0]$_DFFE_PN0P_  (.D(_046_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFFE_PN0P_  (.D(_047_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \valid$_DFFE_PN0P_  (.D(_048_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu9t5v0__buf_16 hold1 (.I(net38),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_72 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_73 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_74 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_75 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_76 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_77 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_78 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_79 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_80 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_81 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_82 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(dividend[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(dividend[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(dividend[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(dividend[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(dividend[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(dividend[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(dividend[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(dividend[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(divisor[0]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(divisor[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(divisor[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(divisor[3]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(divisor[4]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(divisor[5]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(divisor[6]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(divisor[7]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input17 (.I(start),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(busy));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(error));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(quotient[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(quotient[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(quotient[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(quotient[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(quotient[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output25 (.I(net26),
    .Z(quotient[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output26 (.I(net27),
    .Z(quotient[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output27 (.I(net28),
    .Z(quotient[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output28 (.I(net29),
    .Z(remainder[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output29 (.I(net30),
    .Z(remainder[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output30 (.I(net31),
    .Z(remainder[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output31 (.I(net32),
    .Z(remainder[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output32 (.I(net33),
    .Z(remainder[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output33 (.I(net34),
    .Z(remainder[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output34 (.I(net35),
    .Z(remainder[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output35 (.I(net36),
    .Z(remainder[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output36 (.I(net37),
    .Z(valid));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_27 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_307 ();
endmodule
