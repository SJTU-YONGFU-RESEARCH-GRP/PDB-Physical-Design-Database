module fixed_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire \bit_counter[0] ;
 wire \bit_counter[1] ;
 wire \bit_counter[2] ;
 wire \bit_counter[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__inv_3 _119_ (.I(\bit_counter[3] ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _120_ (.A1(\bit_counter[2] ),
    .A2(_101_),
    .A3(_099_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _121_ (.I(_105_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _122_ (.I(\state[0] ),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _123_ (.A1(_098_),
    .A2(\state[1] ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _124_ (.I(_034_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _125_ (.A1(\bit_counter[2] ),
    .A2(\bit_counter[0] ),
    .A3(\bit_counter[1] ),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _126_ (.A1(\bit_counter[3] ),
    .A2(_102_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _127_ (.A1(\bit_counter[2] ),
    .A2(_101_),
    .A3(_099_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _128_ (.I(\state[1] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _129_ (.I(\bit_counter[0] ),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _130_ (.A1(_035_),
    .A2(_036_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _131_ (.I(_108_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _132_ (.A1(net22),
    .A2(_038_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _133_ (.I0(\bit_counter[0] ),
    .I1(_037_),
    .S(_039_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _134_ (.A1(\state[1] ),
    .A2(\bit_counter[0] ),
    .B1(_040_),
    .B2(\state[0] ),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _135_ (.I(_041_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _136_ (.A1(_035_),
    .A2(_100_),
    .Z(_042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _137_ (.I0(\bit_counter[1] ),
    .I1(_042_),
    .S(_039_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _138_ (.A1(\state[1] ),
    .A2(\bit_counter[1] ),
    .B1(_043_),
    .B2(\state[0] ),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _139_ (.I(_044_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _140_ (.A1(_099_),
    .A2(_039_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _141_ (.A1(\state[0] ),
    .A2(_035_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _142_ (.A1(_045_),
    .A2(_046_),
    .Z(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _143_ (.A1(_098_),
    .A2(_045_),
    .B(_035_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _144_ (.I0(_047_),
    .I1(_048_),
    .S(\bit_counter[2] ),
    .Z(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _145_ (.I(_104_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _146_ (.A1(net22),
    .A2(_038_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _147_ (.A1(\state[0] ),
    .A2(_035_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _148_ (.A1(\state[0] ),
    .A2(_050_),
    .B(\state[1] ),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _149_ (.A1(_049_),
    .A2(_050_),
    .A3(_051_),
    .B1(_052_),
    .B2(_101_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _150_ (.I0(\rx_shift_reg[0] ),
    .I1(net13),
    .S(_034_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(\rx_shift_reg[1] ),
    .I1(net14),
    .S(_034_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(\rx_shift_reg[2] ),
    .I1(net15),
    .S(_034_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(\rx_shift_reg[3] ),
    .I1(net16),
    .S(_034_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _154_ (.I0(\rx_shift_reg[4] ),
    .I1(net17),
    .S(_034_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _155_ (.I0(\rx_shift_reg[5] ),
    .I1(net18),
    .S(_034_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _156_ (.I0(\rx_shift_reg[6] ),
    .I1(net19),
    .S(_034_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _157_ (.I0(\rx_shift_reg[7] ),
    .I1(net20),
    .S(_034_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _158_ (.A1(_107_),
    .A2(_115_),
    .A3(_118_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _159_ (.A1(net22),
    .A2(_108_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _160_ (.A1(\bit_counter[2] ),
    .A2(_099_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _161_ (.A1(_100_),
    .A2(_051_),
    .A3(_054_),
    .A4(_055_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _162_ (.I(_111_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _163_ (.A1(\bit_counter[0] ),
    .A2(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _164_ (.A1(_049_),
    .A2(_103_),
    .A3(_114_),
    .A4(_117_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _165_ (.A1(_053_),
    .A2(_056_),
    .A3(_058_),
    .A4(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _166_ (.I0(net3),
    .I1(\rx_shift_reg[0] ),
    .S(_060_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _167_ (.A1(_098_),
    .A2(\state[1] ),
    .A3(_104_),
    .A4(_054_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _168_ (.A1(_100_),
    .A2(_055_),
    .A3(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _169_ (.I(net3),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _170_ (.A1(_057_),
    .A2(_103_),
    .A3(_114_),
    .A4(_117_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _171_ (.A1(_108_),
    .A2(_107_),
    .A3(_115_),
    .A4(_118_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _172_ (.A1(\bit_counter[0] ),
    .A2(_063_),
    .A3(_064_),
    .A4(_065_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _173_ (.A1(_101_),
    .A2(_036_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _174_ (.A1(_067_),
    .A2(_062_),
    .B(\rx_shift_reg[1] ),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _175_ (.A1(_062_),
    .A2(_066_),
    .B(_068_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _176_ (.A1(_036_),
    .A2(_064_),
    .A3(_065_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _177_ (.A1(_100_),
    .A2(_055_),
    .A3(_061_),
    .A4(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _178_ (.I0(\rx_shift_reg[2] ),
    .I1(net3),
    .S(_070_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _179_ (.A1(\bit_counter[2] ),
    .A2(_099_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _180_ (.A1(_100_),
    .A2(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _181_ (.A1(_061_),
    .A2(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _182_ (.A1(_067_),
    .A2(_073_),
    .B(\rx_shift_reg[3] ),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _183_ (.A1(_066_),
    .A2(_073_),
    .B(_074_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _184_ (.A1(_061_),
    .A2(_069_),
    .A3(_072_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _185_ (.I0(net3),
    .I1(\rx_shift_reg[4] ),
    .S(_075_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _186_ (.A1(_100_),
    .A2(_071_),
    .A3(_061_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _187_ (.A1(_067_),
    .A2(_076_),
    .B(\rx_shift_reg[5] ),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _188_ (.A1(_066_),
    .A2(_076_),
    .B(_077_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _189_ (.A1(_100_),
    .A2(_071_),
    .A3(_061_),
    .A4(_069_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _190_ (.I0(\rx_shift_reg[6] ),
    .I1(net3),
    .S(_078_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _191_ (.A1(_104_),
    .A2(_056_),
    .A3(_067_),
    .B(\rx_shift_reg[7] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _192_ (.A1(_104_),
    .A2(_056_),
    .A3(_066_),
    .B(_079_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _193_ (.A1(net22),
    .A2(\state[1] ),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _194_ (.A1(\state[0] ),
    .A2(_080_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _195_ (.A1(_035_),
    .A2(net12),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _196_ (.I0(net23),
    .I1(_081_),
    .S(_098_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _197_ (.I0(net11),
    .I1(\tx_shift_reg[6] ),
    .S(_046_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _198_ (.A1(net22),
    .A2(_106_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _199_ (.I0(net12),
    .I1(_083_),
    .S(\state[0] ),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _200_ (.A1(_035_),
    .A2(_084_),
    .Z(_085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _201_ (.I0(net24),
    .I1(_082_),
    .S(_085_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _202_ (.I(net12),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _203_ (.I(_106_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _204_ (.A1(net22),
    .A2(_087_),
    .A3(_105_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _205_ (.I0(_086_),
    .I1(_088_),
    .S(\state[0] ),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _206_ (.A1(\state[1] ),
    .A2(_089_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _207_ (.A1(_046_),
    .A2(_088_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _208_ (.A1(_098_),
    .A2(_035_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(_086_),
    .I1(net25),
    .S(_090_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _210_ (.A1(net4),
    .A2(_051_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(\tx_shift_reg[0] ),
    .I1(_091_),
    .S(_085_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(net5),
    .I1(\tx_shift_reg[0] ),
    .S(_046_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _213_ (.I0(\tx_shift_reg[1] ),
    .I1(_092_),
    .S(_085_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(net6),
    .I1(\tx_shift_reg[1] ),
    .S(_046_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(\tx_shift_reg[2] ),
    .I1(_093_),
    .S(_085_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(net7),
    .I1(\tx_shift_reg[2] ),
    .S(_046_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _217_ (.I0(\tx_shift_reg[3] ),
    .I1(_094_),
    .S(_085_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _218_ (.I0(net8),
    .I1(\tx_shift_reg[3] ),
    .S(_046_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _219_ (.I0(\tx_shift_reg[4] ),
    .I1(_095_),
    .S(_085_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _220_ (.I0(net9),
    .I1(\tx_shift_reg[4] ),
    .S(_046_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(\tx_shift_reg[5] ),
    .I1(_096_),
    .S(_085_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _222_ (.I0(net10),
    .I1(\tx_shift_reg[5] ),
    .S(_046_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(\tx_shift_reg[6] ),
    .I1(_097_),
    .S(_085_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _224_ (.A(\bit_counter[0] ),
    .B(\bit_counter[1] ),
    .CO(_099_),
    .S(_100_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _225_ (.A(_101_),
    .B(_102_),
    .CO(_103_),
    .S(_104_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _226_ (.A(_101_),
    .B(_105_),
    .CO(_106_),
    .S(_107_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _227_ (.A(\bit_counter[3] ),
    .B(_105_),
    .CO(_108_),
    .S(_109_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _228_ (.A(\bit_counter[3] ),
    .B(_110_),
    .CO(_111_),
    .S(_112_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _229_ (.A(_101_),
    .B(_113_),
    .CO(_114_),
    .S(_115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _230_ (.A(_101_),
    .B(_116_),
    .CO(_117_),
    .S(_118_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[0]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_counter[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[1]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\bit_counter[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[2]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\bit_counter[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_counter[3]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_counter[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[0]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[1]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[2]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[3]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[4]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[5]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[6]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[7]$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFF_PN0_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_022_),
    .SETN(net2),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[1]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_026_),
    .SETN(net2),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[2]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[3]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[4]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[5]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[6]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_65 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_55 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_240 ();
endmodule
