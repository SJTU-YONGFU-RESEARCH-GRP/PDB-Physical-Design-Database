module clock_domain_crossing (dst_clk,
    dst_ready,
    dst_rst_n,
    dst_valid,
    src_clk,
    src_ready,
    src_rst_n,
    src_valid,
    dst_data,
    src_data);
 input dst_clk;
 input dst_ready;
 input dst_rst_n;
 output dst_valid;
 input src_clk;
 output src_ready;
 input src_rst_n;
 input src_valid;
 output [31:0] dst_data;
 input [31:0] src_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire dst_ack;
 wire dst_req_prev;
 wire \dst_req_sync[0] ;
 wire \dst_req_sync[1] ;
 wire src_ack;
 wire \src_ack_sync[0] ;
 wire \src_data_reg[0] ;
 wire \src_data_reg[10] ;
 wire \src_data_reg[11] ;
 wire \src_data_reg[12] ;
 wire \src_data_reg[13] ;
 wire \src_data_reg[14] ;
 wire \src_data_reg[15] ;
 wire \src_data_reg[16] ;
 wire \src_data_reg[17] ;
 wire \src_data_reg[18] ;
 wire \src_data_reg[19] ;
 wire \src_data_reg[1] ;
 wire \src_data_reg[20] ;
 wire \src_data_reg[21] ;
 wire \src_data_reg[22] ;
 wire \src_data_reg[23] ;
 wire \src_data_reg[24] ;
 wire \src_data_reg[25] ;
 wire \src_data_reg[26] ;
 wire \src_data_reg[27] ;
 wire \src_data_reg[28] ;
 wire \src_data_reg[29] ;
 wire \src_data_reg[2] ;
 wire \src_data_reg[30] ;
 wire \src_data_reg[31] ;
 wire \src_data_reg[3] ;
 wire \src_data_reg[4] ;
 wire \src_data_reg[5] ;
 wire \src_data_reg[6] ;
 wire \src_data_reg[7] ;
 wire \src_data_reg[8] ;
 wire \src_data_reg[9] ;
 wire src_req;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire clknet_0_src_clk;
 wire clknet_2_0__leaf_src_clk;
 wire clknet_2_1__leaf_src_clk;
 wire clknet_2_2__leaf_src_clk;
 wire clknet_2_3__leaf_src_clk;
 wire net72;

 sky130_fd_sc_hd__xor2_4 _077_ (.A(dst_req_prev),
    .B(\dst_req_sync[1] ),
    .X(_067_));
 sky130_fd_sc_hd__buf_6 _078_ (.A(_067_),
    .X(_068_));
 sky130_fd_sc_hd__and2_0 _079_ (.A(net4),
    .B(_068_),
    .X(_000_));
 sky130_fd_sc_hd__xnor2_1 _080_ (.A(src_req),
    .B(src_ack),
    .Y(net71));
 sky130_fd_sc_hd__mux2_1 _081_ (.A0(net38),
    .A1(\src_data_reg[0] ),
    .S(_068_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _082_ (.A0(net39),
    .A1(\src_data_reg[10] ),
    .S(_068_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _083_ (.A0(net40),
    .A1(\src_data_reg[11] ),
    .S(_068_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _084_ (.A0(net41),
    .A1(\src_data_reg[12] ),
    .S(_068_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _085_ (.A0(net42),
    .A1(\src_data_reg[13] ),
    .S(_068_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _086_ (.A0(net43),
    .A1(\src_data_reg[14] ),
    .S(_068_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _087_ (.A0(net44),
    .A1(\src_data_reg[15] ),
    .S(_068_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _088_ (.A0(net45),
    .A1(\src_data_reg[16] ),
    .S(_068_),
    .X(_008_));
 sky130_fd_sc_hd__buf_6 _089_ (.A(_067_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _090_ (.A0(net46),
    .A1(\src_data_reg[17] ),
    .S(_069_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _091_ (.A0(net47),
    .A1(\src_data_reg[18] ),
    .S(_069_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _092_ (.A0(net48),
    .A1(\src_data_reg[19] ),
    .S(_069_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _093_ (.A0(net49),
    .A1(\src_data_reg[1] ),
    .S(_069_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _094_ (.A0(net50),
    .A1(\src_data_reg[20] ),
    .S(_069_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _095_ (.A0(net51),
    .A1(\src_data_reg[21] ),
    .S(_069_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _096_ (.A0(net52),
    .A1(\src_data_reg[22] ),
    .S(_069_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _097_ (.A0(net53),
    .A1(\src_data_reg[23] ),
    .S(_069_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _098_ (.A0(net54),
    .A1(\src_data_reg[24] ),
    .S(_069_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _099_ (.A0(net55),
    .A1(\src_data_reg[25] ),
    .S(_069_),
    .X(_018_));
 sky130_fd_sc_hd__buf_6 _100_ (.A(_067_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _101_ (.A0(net56),
    .A1(\src_data_reg[26] ),
    .S(_070_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(net57),
    .A1(\src_data_reg[27] ),
    .S(_070_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _103_ (.A0(net58),
    .A1(\src_data_reg[28] ),
    .S(_070_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _104_ (.A0(net59),
    .A1(\src_data_reg[29] ),
    .S(_070_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _105_ (.A0(net60),
    .A1(\src_data_reg[2] ),
    .S(_070_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _106_ (.A0(net61),
    .A1(\src_data_reg[30] ),
    .S(_070_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _107_ (.A0(net62),
    .A1(\src_data_reg[31] ),
    .S(_070_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _108_ (.A0(net63),
    .A1(\src_data_reg[3] ),
    .S(_070_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _109_ (.A0(net64),
    .A1(\src_data_reg[4] ),
    .S(_070_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _110_ (.A0(net65),
    .A1(\src_data_reg[5] ),
    .S(_070_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _111_ (.A0(net66),
    .A1(\src_data_reg[6] ),
    .S(_067_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _112_ (.A0(net67),
    .A1(\src_data_reg[7] ),
    .S(_067_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _113_ (.A0(net68),
    .A1(\src_data_reg[8] ),
    .S(_067_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _114_ (.A0(net69),
    .A1(\src_data_reg[9] ),
    .S(_067_),
    .X(_032_));
 sky130_fd_sc_hd__inv_1 _115_ (.A(net3),
    .Y(_071_));
 sky130_fd_sc_hd__a21o_1 _116_ (.A1(_071_),
    .A2(net70),
    .B1(_068_),
    .X(_033_));
 sky130_fd_sc_hd__nand2_2 _117_ (.A(net37),
    .B(net71),
    .Y(_072_));
 sky130_fd_sc_hd__buf_6 _118_ (.A(_072_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _119_ (.A0(net5),
    .A1(\src_data_reg[0] ),
    .S(_073_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _120_ (.A0(net6),
    .A1(\src_data_reg[10] ),
    .S(_073_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _121_ (.A0(net7),
    .A1(\src_data_reg[11] ),
    .S(_073_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(net8),
    .A1(\src_data_reg[12] ),
    .S(_073_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _123_ (.A0(net9),
    .A1(\src_data_reg[13] ),
    .S(_073_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _124_ (.A0(net10),
    .A1(\src_data_reg[14] ),
    .S(_073_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _125_ (.A0(net11),
    .A1(\src_data_reg[15] ),
    .S(_073_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _126_ (.A0(net12),
    .A1(\src_data_reg[16] ),
    .S(_073_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _127_ (.A0(net13),
    .A1(\src_data_reg[17] ),
    .S(_073_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _128_ (.A0(net14),
    .A1(\src_data_reg[18] ),
    .S(_073_),
    .X(_043_));
 sky130_fd_sc_hd__buf_6 _129_ (.A(_072_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _130_ (.A0(net15),
    .A1(\src_data_reg[19] ),
    .S(_074_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _131_ (.A0(net16),
    .A1(\src_data_reg[1] ),
    .S(_074_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _132_ (.A0(net17),
    .A1(\src_data_reg[20] ),
    .S(_074_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _133_ (.A0(net18),
    .A1(\src_data_reg[21] ),
    .S(_074_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _134_ (.A0(net19),
    .A1(\src_data_reg[22] ),
    .S(_074_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _135_ (.A0(net20),
    .A1(\src_data_reg[23] ),
    .S(_074_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _136_ (.A0(net21),
    .A1(\src_data_reg[24] ),
    .S(_074_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _137_ (.A0(net22),
    .A1(\src_data_reg[25] ),
    .S(_074_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _138_ (.A0(net23),
    .A1(\src_data_reg[26] ),
    .S(_074_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _139_ (.A0(net24),
    .A1(\src_data_reg[27] ),
    .S(_074_),
    .X(_053_));
 sky130_fd_sc_hd__buf_6 _140_ (.A(_072_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _141_ (.A0(net25),
    .A1(\src_data_reg[28] ),
    .S(_075_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _142_ (.A0(net26),
    .A1(\src_data_reg[29] ),
    .S(_075_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _143_ (.A0(net27),
    .A1(\src_data_reg[2] ),
    .S(_075_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _144_ (.A0(net28),
    .A1(\src_data_reg[30] ),
    .S(_075_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _145_ (.A0(net29),
    .A1(\src_data_reg[31] ),
    .S(_075_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _146_ (.A0(net30),
    .A1(\src_data_reg[3] ),
    .S(_075_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _147_ (.A0(net31),
    .A1(\src_data_reg[4] ),
    .S(_075_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _148_ (.A0(net32),
    .A1(\src_data_reg[5] ),
    .S(_075_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _149_ (.A0(net33),
    .A1(\src_data_reg[6] ),
    .S(_075_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(net34),
    .A1(\src_data_reg[7] ),
    .S(_075_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _151_ (.A0(net35),
    .A1(\src_data_reg[8] ),
    .S(_072_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _152_ (.A0(net36),
    .A1(\src_data_reg[9] ),
    .S(_072_),
    .X(_065_));
 sky130_fd_sc_hd__nor2_1 _153_ (.A(net37),
    .B(src_req),
    .Y(_076_));
 sky130_fd_sc_hd__a21oi_1 _154_ (.A1(net37),
    .A2(src_ack),
    .B1(_076_),
    .Y(_066_));
 sky130_fd_sc_hd__edfxtp_1 \dst_ack$_DFFE_PP_  (.D(\dst_req_sync[1] ),
    .DE(_000_),
    .Q(dst_ack),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[0]$_DFFE_PN0P_  (.D(_001_),
    .Q(net38),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[10]$_DFFE_PN0P_  (.D(_002_),
    .Q(net39),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[11]$_DFFE_PN0P_  (.D(_003_),
    .Q(net40),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[12]$_DFFE_PN0P_  (.D(_004_),
    .Q(net41),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[13]$_DFFE_PN0P_  (.D(_005_),
    .Q(net42),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[14]$_DFFE_PN0P_  (.D(_006_),
    .Q(net43),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[15]$_DFFE_PN0P_  (.D(_007_),
    .Q(net44),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[16]$_DFFE_PN0P_  (.D(_008_),
    .Q(net45),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[17]$_DFFE_PN0P_  (.D(_009_),
    .Q(net46),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[18]$_DFFE_PN0P_  (.D(_010_),
    .Q(net47),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[19]$_DFFE_PN0P_  (.D(_011_),
    .Q(net48),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[1]$_DFFE_PN0P_  (.D(_012_),
    .Q(net49),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[20]$_DFFE_PN0P_  (.D(_013_),
    .Q(net50),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[21]$_DFFE_PN0P_  (.D(_014_),
    .Q(net51),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[22]$_DFFE_PN0P_  (.D(_015_),
    .Q(net52),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[23]$_DFFE_PN0P_  (.D(_016_),
    .Q(net53),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[24]$_DFFE_PN0P_  (.D(_017_),
    .Q(net54),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[25]$_DFFE_PN0P_  (.D(_018_),
    .Q(net55),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[26]$_DFFE_PN0P_  (.D(_019_),
    .Q(net56),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[27]$_DFFE_PN0P_  (.D(_020_),
    .Q(net57),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[28]$_DFFE_PN0P_  (.D(_021_),
    .Q(net58),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[29]$_DFFE_PN0P_  (.D(_022_),
    .Q(net59),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[2]$_DFFE_PN0P_  (.D(_023_),
    .Q(net60),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[30]$_DFFE_PN0P_  (.D(_024_),
    .Q(net61),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[31]$_DFFE_PN0P_  (.D(_025_),
    .Q(net62),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[3]$_DFFE_PN0P_  (.D(_026_),
    .Q(net63),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[4]$_DFFE_PN0P_  (.D(_027_),
    .Q(net64),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[5]$_DFFE_PN0P_  (.D(_028_),
    .Q(net65),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[6]$_DFFE_PN0P_  (.D(_029_),
    .Q(net66),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[7]$_DFFE_PN0P_  (.D(_030_),
    .Q(net67),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[8]$_DFFE_PN0P_  (.D(_031_),
    .Q(net68),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_data[9]$_DFFE_PN0P_  (.D(_032_),
    .Q(net69),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_req_prev$_DFF_PN0_  (.D(\dst_req_sync[1] ),
    .Q(dst_req_prev),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_req_sync[0]$_DFF_PN0_  (.D(src_req),
    .Q(\dst_req_sync[0] ),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_2 \dst_req_sync[1]$_DFF_PN0_  (.D(\dst_req_sync[0] ),
    .Q(\dst_req_sync[1] ),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \dst_valid$_DFFE_PN0P_  (.D(_033_),
    .Q(net70),
    .RESET_B(net4),
    .CLK(net2));
 sky130_fd_sc_hd__dfrtp_1 \src_ack_sync[0]$_DFF_PN0_  (.D(dst_ack),
    .Q(\src_ack_sync[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_ack_sync[1]$_DFF_PN0_  (.D(\src_ack_sync[0] ),
    .Q(src_ack),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[0]$_DFFE_PN0P_  (.D(_034_),
    .Q(\src_data_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[10]$_DFFE_PN0P_  (.D(_035_),
    .Q(\src_data_reg[10] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[11]$_DFFE_PN0P_  (.D(_036_),
    .Q(\src_data_reg[11] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[12]$_DFFE_PN0P_  (.D(_037_),
    .Q(\src_data_reg[12] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[13]$_DFFE_PN0P_  (.D(_038_),
    .Q(\src_data_reg[13] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[14]$_DFFE_PN0P_  (.D(_039_),
    .Q(\src_data_reg[14] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[15]$_DFFE_PN0P_  (.D(_040_),
    .Q(\src_data_reg[15] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[16]$_DFFE_PN0P_  (.D(_041_),
    .Q(\src_data_reg[16] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[17]$_DFFE_PN0P_  (.D(_042_),
    .Q(\src_data_reg[17] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[18]$_DFFE_PN0P_  (.D(_043_),
    .Q(\src_data_reg[18] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[19]$_DFFE_PN0P_  (.D(_044_),
    .Q(\src_data_reg[19] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[1]$_DFFE_PN0P_  (.D(_045_),
    .Q(\src_data_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[20]$_DFFE_PN0P_  (.D(_046_),
    .Q(\src_data_reg[20] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[21]$_DFFE_PN0P_  (.D(_047_),
    .Q(\src_data_reg[21] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[22]$_DFFE_PN0P_  (.D(_048_),
    .Q(\src_data_reg[22] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[23]$_DFFE_PN0P_  (.D(_049_),
    .Q(\src_data_reg[23] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[24]$_DFFE_PN0P_  (.D(_050_),
    .Q(\src_data_reg[24] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[25]$_DFFE_PN0P_  (.D(_051_),
    .Q(\src_data_reg[25] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[26]$_DFFE_PN0P_  (.D(_052_),
    .Q(\src_data_reg[26] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[27]$_DFFE_PN0P_  (.D(_053_),
    .Q(\src_data_reg[27] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[28]$_DFFE_PN0P_  (.D(_054_),
    .Q(\src_data_reg[28] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[29]$_DFFE_PN0P_  (.D(_055_),
    .Q(\src_data_reg[29] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[2]$_DFFE_PN0P_  (.D(_056_),
    .Q(\src_data_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[30]$_DFFE_PN0P_  (.D(_057_),
    .Q(\src_data_reg[30] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[31]$_DFFE_PN0P_  (.D(_058_),
    .Q(\src_data_reg[31] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[3]$_DFFE_PN0P_  (.D(_059_),
    .Q(\src_data_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[4]$_DFFE_PN0P_  (.D(_060_),
    .Q(\src_data_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[5]$_DFFE_PN0P_  (.D(_061_),
    .Q(\src_data_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[6]$_DFFE_PN0P_  (.D(_062_),
    .Q(\src_data_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[7]$_DFFE_PN0P_  (.D(_063_),
    .Q(\src_data_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[8]$_DFFE_PN0P_  (.D(_064_),
    .Q(\src_data_reg[8] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_data_reg[9]$_DFFE_PN0P_  (.D(_065_),
    .Q(\src_data_reg[9] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__dfrtp_1 \src_req$_DFFE_PN0P_  (.D(_066_),
    .Q(src_req),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net72),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_76 ();
 sky130_fd_sc_hd__buf_16 input1 (.A(dst_clk),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dst_ready),
    .X(net3));
 sky130_fd_sc_hd__buf_12 input3 (.A(dst_rst_n),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(src_data[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(src_data[10]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(src_data[11]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(src_data[12]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(src_data[13]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(src_data[14]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(src_data[15]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(src_data[16]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(src_data[17]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(src_data[18]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(src_data[19]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(src_data[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(src_data[20]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(src_data[21]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(src_data[22]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(src_data[23]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(src_data[24]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(src_data[25]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(src_data[26]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(src_data[27]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(src_data[28]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(src_data[29]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(src_data[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(src_data[30]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(src_data[31]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(src_data[3]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(src_data[4]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(src_data[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(src_data[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(src_data[7]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(src_data[8]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(src_data[9]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(src_valid),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(dst_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(dst_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(dst_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(dst_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(dst_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(dst_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(dst_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(dst_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(dst_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(dst_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(dst_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(dst_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(dst_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(dst_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(dst_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(dst_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(dst_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net55),
    .X(dst_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net56),
    .X(dst_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net57),
    .X(dst_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net58),
    .X(dst_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net59),
    .X(dst_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net60),
    .X(dst_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net61),
    .X(dst_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net62),
    .X(dst_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net63),
    .X(dst_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net64),
    .X(dst_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net65),
    .X(dst_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net66),
    .X(dst_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net67),
    .X(dst_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(dst_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(dst_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(dst_valid));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(src_ready));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_src_clk (.A(src_clk),
    .X(clknet_0_src_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_src_clk (.A(clknet_0_src_clk),
    .X(clknet_2_0__leaf_src_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_src_clk (.A(clknet_0_src_clk),
    .X(clknet_2_1__leaf_src_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_src_clk (.A(clknet_0_src_clk),
    .X(clknet_2_2__leaf_src_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_src_clk (.A(clknet_0_src_clk),
    .X(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_2_3__leaf_src_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(src_rst_n),
    .X(net72));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
endmodule
