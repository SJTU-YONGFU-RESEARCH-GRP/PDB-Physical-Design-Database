module ahb_lite_master (hbusreq,
    hclk,
    hgrant,
    hready,
    hreset,
    hwrite,
    start_trans,
    trans_done,
    trans_write,
    haddr,
    hburst,
    hrdata,
    hresp,
    hsize,
    htrans,
    hwdata,
    read_data,
    trans_addr,
    trans_burst,
    trans_resp,
    trans_size,
    write_data);
 output hbusreq;
 input hclk;
 input hgrant;
 input hready;
 input hreset;
 output hwrite;
 input start_trans;
 output trans_done;
 input trans_write;
 output [31:0] haddr;
 output [2:0] hburst;
 input [31:0] hrdata;
 input [1:0] hresp;
 output [2:0] hsize;
 output [1:0] htrans;
 output [31:0] hwdata;
 output [31:0] read_data;
 input [31:0] trans_addr;
 input [2:0] trans_burst;
 output [1:0] trans_resp;
 input [2:0] trans_size;
 input [31:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire \burst_count[0] ;
 wire \burst_count[1] ;
 wire \burst_count[2] ;
 wire \burst_count[3] ;
 wire \burst_count[4] ;
 wire \burst_count[5] ;
 wire \burst_count[6] ;
 wire \burst_count[7] ;
 wire \burst_total[0] ;
 wire \burst_total[2] ;
 wire \burst_total[3] ;
 wire \burst_total[4] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;

 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _0521_ (.A1(\burst_total[3] ),
    .A2(\burst_total[2] ),
    .A3(\burst_total[0] ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0522_ (.I(\burst_total[4] ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0523_ (.A1(\burst_total[3] ),
    .A2(_0489_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0524_ (.I(net149),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0525_ (.A1(net147),
    .A2(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0526_ (.A1(net148),
    .A2(_0122_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0527_ (.I(_0465_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0528_ (.I(net148),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0529_ (.A1(_0123_),
    .A2(net147),
    .A3(net149),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0530_ (.A1(_0123_),
    .A2(_0122_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0531_ (.A1(net148),
    .A2(net147),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0532_ (.A1(net149),
    .A2(_0124_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0533_ (.A1(_0123_),
    .A2(net147),
    .A3(net149),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0534_ (.A1(_0123_),
    .A2(net147),
    .A3(_0121_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0535_ (.A1(net148),
    .A2(net147),
    .A3(net149),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0536_ (.I(\state[0] ),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _0537_ (.I(\state[1] ),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0538_ (.I(net35),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0539_ (.A1(\state[2] ),
    .A2(_0125_),
    .A3(_0126_),
    .A4(_0127_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0540_ (.I(_0485_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0541_ (.A1(_0492_),
    .A2(_0491_),
    .B(_0486_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0542_ (.A1(\burst_total[0] ),
    .A2(\burst_count[0] ),
    .B(_0494_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0543_ (.A1(_0485_),
    .A2(_0491_),
    .A3(_0493_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0544_ (.A1(_0471_),
    .A2(_0474_),
    .A3(_0477_),
    .A4(_0483_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_4 _0545_ (.A1(_0129_),
    .A2(_0130_),
    .B1(_0131_),
    .B2(_0132_),
    .C(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0546_ (.A1(_0471_),
    .A2(_0474_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0547_ (.A1(_0482_),
    .A2(_0477_),
    .B(_0476_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0548_ (.A1(_0471_),
    .A2(_0473_),
    .B(_0470_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0549_ (.A1(_0135_),
    .A2(_0136_),
    .B(_0137_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0550_ (.I(_0480_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0551_ (.A1(_0134_),
    .A2(_0138_),
    .B(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _0552_ (.A1(_0128_),
    .A2(_0140_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0553_ (.I(\state[1] ),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0554_ (.I0(net2),
    .I1(net35),
    .S(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0555_ (.A1(_0126_),
    .A2(net39),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _0556_ (.A1(_0142_),
    .A2(net35),
    .B(_0144_),
    .C(\state[0] ),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _0557_ (.A1(\state[0] ),
    .A2(_0143_),
    .B(_0145_),
    .C(\state[2] ),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0558_ (.A1(_0141_),
    .A2(_0146_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0559_ (.A1(_0142_),
    .A2(_0127_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0560_ (.A1(\state[0] ),
    .A2(_0126_),
    .A3(net2),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0561_ (.A1(_0147_),
    .A2(_0148_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0562_ (.A1(\state[2] ),
    .A2(_0142_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0563_ (.A1(\state[2] ),
    .A2(_0149_),
    .B1(_0150_),
    .B2(\state[0] ),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0564_ (.I(_0128_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0565_ (.I(net122),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0566_ (.I(_0496_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0567_ (.I(\burst_total[0] ),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0568_ (.I(_0489_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0569_ (.A1(\burst_total[3] ),
    .A2(\burst_total[4] ),
    .A3(_0151_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0570_ (.A1(_0478_),
    .A2(_0479_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0571_ (.A1(_0478_),
    .A2(_0479_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0572_ (.I(\burst_total[2] ),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0573_ (.A1(_0121_),
    .A2(_0124_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _0574_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0575_ (.A1(\state[1] ),
    .A2(net35),
    .A3(_0152_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0576_ (.A1(_0140_),
    .A2(_0153_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0577_ (.A1(\state[1] ),
    .A2(_0152_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _0578_ (.A1(_0127_),
    .A2(_0134_),
    .A3(_0138_),
    .A4(_0155_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__and3_4 _0579_ (.A1(_0126_),
    .A2(net39),
    .A3(_0152_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0580_ (.A1(_0480_),
    .A2(_0153_),
    .B(_0157_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0581_ (.A1(_0156_),
    .A2(_0158_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0582_ (.I0(_0154_),
    .I1(_0159_),
    .S(\burst_count[0] ),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0583_ (.A1(_0142_),
    .A2(_0152_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0584_ (.A1(_0520_),
    .A2(_0160_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0585_ (.A1(_0156_),
    .A2(_0158_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0586_ (.I0(\burst_count[1] ),
    .I1(_0161_),
    .S(_0162_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0587_ (.A1(_0144_),
    .A2(_0152_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0588_ (.I(\burst_count[2] ),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0589_ (.I(_0519_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0590_ (.A1(_0156_),
    .A2(_0158_),
    .B(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0591_ (.A1(_0164_),
    .A2(_0166_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0592_ (.A1(_0163_),
    .A2(_0167_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0593_ (.I(\burst_count[3] ),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0594_ (.A1(\burst_count[2] ),
    .A2(\burst_count[0] ),
    .A3(\burst_count[1] ),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0595_ (.A1(_0156_),
    .A2(_0158_),
    .B(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0596_ (.A1(_0168_),
    .A2(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0597_ (.A1(_0163_),
    .A2(_0171_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0598_ (.I(\burst_count[4] ),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0599_ (.A1(_0164_),
    .A2(_0165_),
    .A3(_0168_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0600_ (.A1(_0156_),
    .A2(_0158_),
    .B(_0173_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0601_ (.A1(_0172_),
    .A2(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0602_ (.A1(_0163_),
    .A2(_0175_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0603_ (.A1(\burst_count[5] ),
    .A2(_0163_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0604_ (.A1(\burst_count[5] ),
    .A2(_0157_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0605_ (.A1(_0172_),
    .A2(_0169_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0606_ (.A1(\burst_count[3] ),
    .A2(_0162_),
    .A3(_0178_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0607_ (.I0(_0176_),
    .I1(_0177_),
    .S(_0179_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0608_ (.A1(\burst_count[4] ),
    .A2(\burst_count[2] ),
    .A3(_0519_),
    .A4(\burst_count[3] ),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0609_ (.A1(\burst_count[5] ),
    .A2(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0610_ (.A1(_0159_),
    .A2(_0181_),
    .B(\burst_count[6] ),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0611_ (.A1(\burst_count[6] ),
    .A2(_0159_),
    .A3(_0181_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0612_ (.A1(_0182_),
    .A2(_0183_),
    .B(_0157_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0613_ (.A1(\burst_count[6] ),
    .A2(\burst_count[5] ),
    .A3(\burst_count[3] ),
    .A4(_0178_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0614_ (.A1(_0159_),
    .A2(_0184_),
    .B(\burst_count[7] ),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0615_ (.A1(\burst_count[7] ),
    .A2(_0159_),
    .A3(_0184_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0616_ (.A1(_0185_),
    .A2(_0186_),
    .B(_0157_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0617_ (.A1(net74),
    .A2(net72),
    .A3(net73),
    .A4(_0163_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0618_ (.A1(_0487_),
    .A2(_0157_),
    .B(_0187_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0619_ (.I(net72),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0620_ (.I(net73),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0621_ (.A1(_0188_),
    .A2(_0189_),
    .B(net74),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0622_ (.I0(\burst_total[2] ),
    .I1(_0190_),
    .S(_0157_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0623_ (.A1(net74),
    .A2(_0189_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0624_ (.I0(\burst_total[3] ),
    .I1(_0191_),
    .S(_0157_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0625_ (.A1(net74),
    .A2(net73),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0626_ (.I0(\burst_total[4] ),
    .I1(_0192_),
    .S(_0157_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0627_ (.I(\state[2] ),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0628_ (.A1(_0193_),
    .A2(\state[0] ),
    .A3(_0126_),
    .A4(net2),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0629_ (.I(_0194_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0630_ (.I0(net143),
    .I1(net72),
    .S(_0195_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0631_ (.I0(net144),
    .I1(net73),
    .S(_0195_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0632_ (.I0(net145),
    .I1(net74),
    .S(_0195_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0633_ (.A1(\state[2] ),
    .A2(_0125_),
    .A3(_0142_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0634_ (.I(_0155_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0635_ (.A1(net39),
    .A2(_0197_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0636_ (.A1(_0196_),
    .A2(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0637_ (.A1(_0125_),
    .A2(net35),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0638_ (.A1(net145),
    .A2(net144),
    .A3(net143),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0639_ (.A1(_0140_),
    .A2(_0160_),
    .A3(_0201_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _0640_ (.A1(_0142_),
    .A2(_0200_),
    .B(_0202_),
    .C(\state[2] ),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0641_ (.I0(net146),
    .I1(_0199_),
    .S(_0203_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0642_ (.I0(net147),
    .I1(net75),
    .S(_0195_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0643_ (.I0(net148),
    .I1(net76),
    .S(_0195_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0644_ (.I0(net149),
    .I1(net77),
    .S(_0195_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0645_ (.I(net150),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0646_ (.A1(_0193_),
    .A2(_0126_),
    .A3(net2),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0647_ (.A1(_0147_),
    .A2(_0152_),
    .B(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0648_ (.A1(net2),
    .A2(_0196_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0649_ (.A1(_0204_),
    .A2(_0206_),
    .B1(_0203_),
    .B2(_0207_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0650_ (.I(net151),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0651_ (.A1(_0208_),
    .A2(_0206_),
    .B1(_0203_),
    .B2(_0196_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0652_ (.A1(net184),
    .A2(_0153_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0653_ (.I(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0654_ (.I0(net152),
    .I1(net79),
    .S(_0210_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0655_ (.I0(net153),
    .I1(net80),
    .S(_0210_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0656_ (.I0(net154),
    .I1(net81),
    .S(_0210_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0657_ (.I0(net155),
    .I1(net82),
    .S(_0210_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0658_ (.I0(net156),
    .I1(net83),
    .S(_0210_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0659_ (.I0(net157),
    .I1(net84),
    .S(_0210_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0660_ (.I0(net158),
    .I1(net85),
    .S(_0210_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0661_ (.I0(net159),
    .I1(net86),
    .S(_0210_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0662_ (.I0(net160),
    .I1(net87),
    .S(_0210_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0663_ (.I0(net161),
    .I1(net88),
    .S(_0210_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0664_ (.I(_0209_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0665_ (.I0(net162),
    .I1(net89),
    .S(_0211_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0666_ (.I0(net163),
    .I1(net90),
    .S(_0211_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0667_ (.I0(net164),
    .I1(net91),
    .S(_0211_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0668_ (.I0(net165),
    .I1(net92),
    .S(_0211_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0669_ (.I0(net166),
    .I1(net93),
    .S(_0211_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0670_ (.I0(net167),
    .I1(net94),
    .S(_0211_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0671_ (.I0(net168),
    .I1(net95),
    .S(_0211_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0672_ (.I0(net169),
    .I1(net96),
    .S(_0211_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0673_ (.I0(net170),
    .I1(net97),
    .S(_0211_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0674_ (.I0(net171),
    .I1(net98),
    .S(_0211_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0675_ (.I(_0209_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0676_ (.I0(net172),
    .I1(net99),
    .S(_0212_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0677_ (.I0(net173),
    .I1(net100),
    .S(_0212_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0678_ (.I0(net174),
    .I1(net101),
    .S(_0212_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0679_ (.I0(net175),
    .I1(net102),
    .S(_0212_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0680_ (.I0(net176),
    .I1(net103),
    .S(_0212_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0681_ (.I0(net177),
    .I1(net104),
    .S(_0212_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0682_ (.I0(net178),
    .I1(net105),
    .S(_0212_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0683_ (.I0(net179),
    .I1(net106),
    .S(_0212_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0684_ (.I0(net180),
    .I1(net107),
    .S(_0212_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0685_ (.I0(net181),
    .I1(net108),
    .S(_0212_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0686_ (.I0(net182),
    .I1(net109),
    .S(_0209_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0687_ (.I0(net183),
    .I1(net110),
    .S(_0209_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0688_ (.I0(net184),
    .I1(net78),
    .S(_0195_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0689_ (.A1(net145),
    .A2(net144),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0690_ (.A1(net143),
    .A2(_0213_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _0691_ (.A1(_0155_),
    .A2(_0214_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0692_ (.I(_0215_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0693_ (.A1(net40),
    .A2(_0197_),
    .B1(_0216_),
    .B2(_0497_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0694_ (.I(_0217_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0695_ (.A1(_0142_),
    .A2(net35),
    .A3(_0152_),
    .A4(_0201_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0696_ (.A1(_0134_),
    .A2(_0138_),
    .A3(_0219_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0697_ (.A1(_0142_),
    .A2(net35),
    .A3(_0152_),
    .A4(_0201_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0698_ (.A1(_0480_),
    .A2(_0221_),
    .B(_0195_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _0699_ (.A1(_0220_),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0700_ (.I0(net111),
    .I1(_0218_),
    .S(_0223_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0701_ (.I(net112),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0702_ (.A1(_0515_),
    .A2(_0514_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0703_ (.A1(_0518_),
    .A2(_0225_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0704_ (.A1(net141),
    .A2(net142),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0705_ (.A1(_0517_),
    .A2(_0226_),
    .B(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0706_ (.A1(_0506_),
    .A2(_0505_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0707_ (.A1(_0509_),
    .A2(_0512_),
    .A3(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0708_ (.I(_0503_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0709_ (.I(_0502_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0710_ (.I(_0505_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _0711_ (.A1(_0467_),
    .A2(_0231_),
    .B(_0232_),
    .C(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0712_ (.A1(_0512_),
    .A2(_0508_),
    .B(_0511_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0713_ (.I(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0714_ (.A1(_0518_),
    .A2(_0514_),
    .B(_0517_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0715_ (.I(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _0716_ (.A1(_0230_),
    .A2(_0234_),
    .B(_0236_),
    .C(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0717_ (.I(_0239_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0718_ (.A1(_0228_),
    .A2(_0240_),
    .B(_0216_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0719_ (.A1(_0223_),
    .A2(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0720_ (.I(_0155_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0721_ (.A1(_0228_),
    .A2(_0239_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0722_ (.A1(_0224_),
    .A2(_0216_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0723_ (.A1(net41),
    .A2(_0243_),
    .B1(_0244_),
    .B2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0724_ (.A1(_0220_),
    .A2(_0222_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0725_ (.I(_0247_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0726_ (.A1(_0224_),
    .A2(_0242_),
    .B1(_0246_),
    .B2(_0248_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0727_ (.I(_0247_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0728_ (.I(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0729_ (.I(_0155_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0730_ (.I(net113),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0731_ (.I(_0511_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0732_ (.A1(_0515_),
    .A2(_0518_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0733_ (.A1(_0512_),
    .A2(_0515_),
    .A3(_0518_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0734_ (.A1(_0509_),
    .A2(_0505_),
    .B(_0508_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0735_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0255_),
    .B2(_0256_),
    .C(_0237_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _0736_ (.A1(_0503_),
    .A2(_0502_),
    .B(_0509_),
    .C(_0506_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _0737_ (.A1(_0496_),
    .A2(_0500_),
    .B(_0499_),
    .C(_0502_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0738_ (.A1(_0255_),
    .A2(_0258_),
    .A3(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0739_ (.A1(_0257_),
    .A2(_0260_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0740_ (.I(_0261_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0741_ (.I(_0227_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0742_ (.A1(net112),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0743_ (.A1(_0252_),
    .A2(_0216_),
    .A3(_0262_),
    .A4(_0264_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0744_ (.A1(net42),
    .A2(_0251_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0745_ (.I(_0247_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__or2_4 _0746_ (.A1(_0155_),
    .A2(_0214_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0747_ (.A1(_0262_),
    .A2(_0264_),
    .B(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0748_ (.A1(_0267_),
    .A2(_0269_),
    .B(net113),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0749_ (.A1(_0250_),
    .A2(_0266_),
    .B(_0270_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0750_ (.I(net114),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _0751_ (.A1(_0230_),
    .A2(_0234_),
    .B(_0236_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0752_ (.A1(_0515_),
    .A2(_0518_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0753_ (.A1(net112),
    .A2(net113),
    .A3(_0263_),
    .A4(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0754_ (.A1(net112),
    .A2(net113),
    .A3(_0263_),
    .A4(_0238_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _0755_ (.A1(_0272_),
    .A2(_0274_),
    .B(_0275_),
    .C(_0216_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0756_ (.A1(_0223_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0757_ (.A1(_0272_),
    .A2(_0274_),
    .B(_0275_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0758_ (.I(_0215_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0759_ (.A1(_0271_),
    .A2(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0760_ (.A1(net43),
    .A2(_0243_),
    .B1(_0278_),
    .B2(_0280_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0761_ (.A1(_0271_),
    .A2(_0277_),
    .B1(_0281_),
    .B2(_0248_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0762_ (.A1(net112),
    .A2(net113),
    .A3(net114),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0763_ (.A1(_0215_),
    .A2(_0263_),
    .A3(_0261_),
    .A4(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0764_ (.I(net115),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0765_ (.A1(net44),
    .A2(_0251_),
    .B1(_0283_),
    .B2(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0766_ (.I(_0215_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0767_ (.A1(_0263_),
    .A2(_0262_),
    .A3(_0282_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0768_ (.A1(_0286_),
    .A2(_0287_),
    .B(_0249_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0769_ (.A1(_0250_),
    .A2(_0285_),
    .B1(_0288_),
    .B2(_0284_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0770_ (.I(net116),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0771_ (.A1(net115),
    .A2(_0289_),
    .A3(_0215_),
    .A4(_0282_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0772_ (.A1(net45),
    .A2(_0251_),
    .B1(_0244_),
    .B2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0773_ (.A1(net115),
    .A2(_0244_),
    .A3(_0282_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0774_ (.A1(net116),
    .A2(_0286_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0775_ (.A1(net116),
    .A2(_0267_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0776_ (.A1(_0250_),
    .A2(_0291_),
    .B1(_0292_),
    .B2(_0293_),
    .C(_0294_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0777_ (.I(net117),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _0778_ (.I(_0216_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0779_ (.A1(net115),
    .A2(net116),
    .A3(_0227_),
    .A4(_0282_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0780_ (.A1(_0262_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0781_ (.I(_0247_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0782_ (.A1(_0296_),
    .A2(_0298_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0783_ (.A1(_0295_),
    .A2(_0279_),
    .A3(_0262_),
    .A4(_0297_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0784_ (.A1(net46),
    .A2(_0251_),
    .B(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0785_ (.A1(_0295_),
    .A2(_0300_),
    .B1(_0302_),
    .B2(_0248_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0786_ (.I(net118),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0787_ (.A1(net115),
    .A2(net116),
    .A3(net117),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0788_ (.A1(_0282_),
    .A2(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _0789_ (.A1(_0517_),
    .A2(_0226_),
    .B(_0305_),
    .C(_0227_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _0790_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0791_ (.A1(_0240_),
    .A2(_0307_),
    .B(_0216_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0792_ (.A1(_0223_),
    .A2(_0308_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_4 _0793_ (.A1(_0268_),
    .A2(_0239_),
    .A3(_0306_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0794_ (.A1(net47),
    .A2(_0243_),
    .B1(_0310_),
    .B2(_0303_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0795_ (.A1(_0303_),
    .A2(_0309_),
    .B1(_0311_),
    .B2(_0248_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0796_ (.A1(_0263_),
    .A2(_0261_),
    .A3(_0282_),
    .A4(_0304_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0797_ (.A1(_0303_),
    .A2(net119),
    .A3(_0268_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0798_ (.A1(net48),
    .A2(_0251_),
    .B1(_0312_),
    .B2(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0799_ (.A1(net118),
    .A2(_0312_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0800_ (.A1(net119),
    .A2(_0286_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0801_ (.A1(net119),
    .A2(_0267_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0802_ (.A1(_0250_),
    .A2(_0314_),
    .B1(_0315_),
    .B2(_0316_),
    .C(_0317_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0803_ (.A1(net118),
    .A2(net119),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0804_ (.A1(net120),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0805_ (.A1(net49),
    .A2(_0251_),
    .B1(_0310_),
    .B2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0806_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0318_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0807_ (.A1(_0286_),
    .A2(_0321_),
    .B(_0249_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0808_ (.I(net120),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0809_ (.A1(_0250_),
    .A2(_0320_),
    .B1(_0322_),
    .B2(_0323_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0810_ (.I(net121),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0811_ (.A1(_0323_),
    .A2(_0318_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0812_ (.A1(_0263_),
    .A2(_0262_),
    .A3(_0305_),
    .A4(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0813_ (.A1(_0296_),
    .A2(_0326_),
    .B(_0299_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0814_ (.A1(_0263_),
    .A2(_0261_),
    .A3(_0305_),
    .A4(_0325_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0815_ (.A1(_0324_),
    .A2(_0279_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0816_ (.A1(net50),
    .A2(_0243_),
    .B1(_0328_),
    .B2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0817_ (.A1(_0324_),
    .A2(_0327_),
    .B1(_0330_),
    .B2(_0248_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _0818_ (.A1(net51),
    .A2(_0197_),
    .B1(_0286_),
    .B2(_0468_),
    .C(_0249_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0819_ (.A1(_0464_),
    .A2(_0250_),
    .B(_0331_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0820_ (.I(net123),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0821_ (.A1(net118),
    .A2(net119),
    .A3(net120),
    .A4(net121),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0822_ (.I(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0823_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0334_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0824_ (.A1(_0296_),
    .A2(_0335_),
    .B(_0299_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _0825_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0334_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0826_ (.A1(_0332_),
    .A2(_0279_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0827_ (.A1(net52),
    .A2(_0243_),
    .B1(_0337_),
    .B2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0828_ (.A1(_0332_),
    .A2(_0336_),
    .B1(_0339_),
    .B2(_0248_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0829_ (.I(net124),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0830_ (.A1(net123),
    .A2(_0340_),
    .A3(_0304_),
    .A4(_0333_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0831_ (.A1(net53),
    .A2(_0251_),
    .B1(_0283_),
    .B2(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0832_ (.A1(net123),
    .A2(_0312_),
    .A3(_0333_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0833_ (.A1(net124),
    .A2(_0286_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0834_ (.A1(net124),
    .A2(_0299_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0835_ (.A1(_0250_),
    .A2(_0342_),
    .B1(_0343_),
    .B2(_0344_),
    .C(_0345_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0836_ (.I(net125),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0837_ (.A1(net123),
    .A2(net124),
    .A3(_0333_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0838_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0839_ (.A1(_0296_),
    .A2(_0348_),
    .B(_0299_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0840_ (.A1(net125),
    .A2(_0347_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0841_ (.A1(net54),
    .A2(_0243_),
    .B1(_0310_),
    .B2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0842_ (.A1(_0346_),
    .A2(_0349_),
    .B1(_0351_),
    .B2(_0248_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0843_ (.I(net126),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0844_ (.A1(net123),
    .A2(net124),
    .A3(net125),
    .A4(_0333_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _0845_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_2 _0846_ (.A1(_0263_),
    .A2(_0262_),
    .A3(_0305_),
    .A4(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0847_ (.A1(_0296_),
    .A2(_0355_),
    .B(_0299_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0848_ (.A1(_0263_),
    .A2(_0261_),
    .A3(_0305_),
    .A4(_0354_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0849_ (.A1(_0352_),
    .A2(_0279_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0850_ (.A1(net55),
    .A2(_0243_),
    .B1(_0357_),
    .B2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0851_ (.A1(_0352_),
    .A2(_0356_),
    .B1(_0359_),
    .B2(_0248_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0852_ (.I(net127),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0853_ (.A1(_0346_),
    .A2(_0347_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0854_ (.A1(_0352_),
    .A2(_0240_),
    .A3(_0307_),
    .A4(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0855_ (.A1(_0296_),
    .A2(_0362_),
    .B(_0299_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0856_ (.A1(net126),
    .A2(_0360_),
    .A3(_0354_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0857_ (.A1(net56),
    .A2(_0243_),
    .B1(_0310_),
    .B2(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0858_ (.A1(_0360_),
    .A2(_0363_),
    .B1(_0365_),
    .B2(_0248_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0859_ (.A1(net126),
    .A2(net127),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0860_ (.A1(_0312_),
    .A2(_0354_),
    .A3(_0366_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0861_ (.A1(net128),
    .A2(_0286_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0862_ (.I(net128),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0863_ (.A1(_0369_),
    .A2(_0215_),
    .A3(_0354_),
    .A4(_0366_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0864_ (.A1(net57),
    .A2(_0197_),
    .B1(_0312_),
    .B2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0865_ (.A1(net128),
    .A2(_0299_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0866_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0371_),
    .B2(_0267_),
    .C(_0372_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0867_ (.I(net129),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0868_ (.A1(net128),
    .A2(_0366_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0869_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0361_),
    .A4(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0870_ (.A1(_0296_),
    .A2(_0375_),
    .B(_0249_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0871_ (.A1(net128),
    .A2(_0373_),
    .A3(_0354_),
    .A4(_0366_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0872_ (.A1(net58),
    .A2(_0197_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0873_ (.A1(_0310_),
    .A2(_0377_),
    .B(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0874_ (.A1(_0373_),
    .A2(_0376_),
    .B1(_0379_),
    .B2(_0267_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0875_ (.I(net130),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0876_ (.A1(net126),
    .A2(net127),
    .A3(net128),
    .A4(net129),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0877_ (.A1(_0380_),
    .A2(_0279_),
    .A3(_0381_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0878_ (.A1(net59),
    .A2(_0243_),
    .B1(_0357_),
    .B2(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0879_ (.A1(_0357_),
    .A2(_0381_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0880_ (.A1(net130),
    .A2(_0286_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0881_ (.A1(net130),
    .A2(_0299_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0882_ (.A1(_0250_),
    .A2(_0383_),
    .B1(_0384_),
    .B2(_0385_),
    .C(_0386_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0883_ (.I(net131),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0884_ (.A1(net130),
    .A2(_0381_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0885_ (.A1(_0240_),
    .A2(_0307_),
    .A3(_0361_),
    .A4(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0886_ (.A1(_0296_),
    .A2(_0389_),
    .B(_0249_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0887_ (.A1(net130),
    .A2(_0387_),
    .A3(_0354_),
    .A4(_0381_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0888_ (.A1(net60),
    .A2(_0197_),
    .B1(_0310_),
    .B2(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0889_ (.A1(_0387_),
    .A2(_0390_),
    .B1(_0392_),
    .B2(_0267_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0890_ (.I(net132),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0891_ (.A1(net130),
    .A2(net131),
    .A3(_0381_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0892_ (.A1(_0393_),
    .A2(_0279_),
    .A3(_0354_),
    .A4(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0893_ (.A1(net61),
    .A2(_0243_),
    .B1(_0312_),
    .B2(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0894_ (.A1(_0312_),
    .A2(_0354_),
    .A3(_0394_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0895_ (.A1(net132),
    .A2(_0286_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0896_ (.A1(net132),
    .A2(_0299_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__oai221_2 _0897_ (.A1(_0248_),
    .A2(_0396_),
    .B1(_0397_),
    .B2(_0398_),
    .C(_0399_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0898_ (.A1(_0467_),
    .A2(_0503_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0899_ (.A1(net62),
    .A2(_0197_),
    .B1(_0216_),
    .B2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0900_ (.I(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0901_ (.I0(net133),
    .I1(_0402_),
    .S(_0223_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0902_ (.I(net134),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0903_ (.A1(_0354_),
    .A2(_0394_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _0904_ (.A1(_0393_),
    .A2(_0239_),
    .A3(_0307_),
    .A4(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0905_ (.A1(_0296_),
    .A2(_0405_),
    .B(_0249_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _0906_ (.A1(_0393_),
    .A2(_0240_),
    .A3(_0307_),
    .A4(_0404_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _0907_ (.A1(_0403_),
    .A2(_0279_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0908_ (.A1(net63),
    .A2(_0197_),
    .B1(_0407_),
    .B2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0909_ (.A1(_0403_),
    .A2(_0406_),
    .B1(_0409_),
    .B2(_0267_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0910_ (.I(net135),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0911_ (.A1(net132),
    .A2(net134),
    .A3(_0227_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0912_ (.A1(_0305_),
    .A2(_0353_),
    .A3(_0394_),
    .A4(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0913_ (.A1(_0262_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0914_ (.A1(_0296_),
    .A2(_0413_),
    .B(_0249_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0915_ (.A1(_0410_),
    .A2(_0279_),
    .A3(_0262_),
    .A4(_0412_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0916_ (.A1(net64),
    .A2(_0251_),
    .B(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0917_ (.A1(_0410_),
    .A2(_0414_),
    .B1(_0416_),
    .B2(_0267_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0918_ (.A1(_0496_),
    .A2(_0500_),
    .B(_0499_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0919_ (.A1(_0231_),
    .A2(_0417_),
    .B(_0232_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0920_ (.A1(_0506_),
    .A2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0921_ (.A1(net65),
    .A2(_0155_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0922_ (.A1(_0268_),
    .A2(_0419_),
    .B(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0923_ (.I0(net136),
    .I1(_0421_),
    .S(_0223_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0924_ (.A1(_0467_),
    .A2(_0231_),
    .B(_0232_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0925_ (.A1(_0506_),
    .A2(_0422_),
    .B(_0505_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _0926_ (.A1(_0509_),
    .A2(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0927_ (.A1(net66),
    .A2(_0155_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0928_ (.A1(_0268_),
    .A2(_0424_),
    .B(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0929_ (.I0(net137),
    .I1(_0426_),
    .S(_0223_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0930_ (.A1(_0258_),
    .A2(_0259_),
    .B(_0256_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _0931_ (.A1(_0512_),
    .A2(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0932_ (.A1(net67),
    .A2(_0197_),
    .B1(_0216_),
    .B2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0933_ (.I(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0934_ (.I0(net138),
    .I1(_0430_),
    .S(_0223_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _0935_ (.A1(_0509_),
    .A2(_0512_),
    .A3(_0229_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0936_ (.I(_0467_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _0937_ (.A1(_0432_),
    .A2(_0503_),
    .B(_0502_),
    .C(_0505_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0938_ (.A1(_0431_),
    .A2(_0433_),
    .B(_0235_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _0939_ (.A1(_0515_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0940_ (.A1(net68),
    .A2(_0155_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0941_ (.A1(_0268_),
    .A2(_0435_),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0942_ (.I0(net139),
    .I1(_0437_),
    .S(_0223_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0943_ (.I(net140),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0944_ (.A1(_0511_),
    .A2(_0514_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _0945_ (.A1(_0258_),
    .A2(_0259_),
    .B(_0439_),
    .C(_0256_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _0946_ (.A1(_0512_),
    .A2(_0511_),
    .A3(_0514_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _0947_ (.A1(_0225_),
    .A2(_0440_),
    .A3(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _0948_ (.A1(_0518_),
    .A2(_0442_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _0949_ (.A1(net69),
    .A2(_0197_),
    .B1(_0216_),
    .B2(_0443_),
    .C(_0249_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0950_ (.A1(_0438_),
    .A2(_0250_),
    .B(_0444_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0951_ (.A1(_0272_),
    .A2(_0254_),
    .B(_0237_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _0952_ (.A1(net141),
    .A2(_0268_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _0953_ (.A1(net70),
    .A2(_0251_),
    .B1(_0445_),
    .B2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _0954_ (.A1(_0434_),
    .A2(_0273_),
    .B(_0268_),
    .C(_0238_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0955_ (.A1(_0267_),
    .A2(_0448_),
    .B(net141),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _0956_ (.A1(_0250_),
    .A2(_0447_),
    .B(_0449_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _0957_ (.I(net142),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _0958_ (.A1(net141),
    .A2(_0262_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0959_ (.A1(_0286_),
    .A2(_0451_),
    .B(_0249_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _0960_ (.A1(net141),
    .A2(_0450_),
    .A3(_0279_),
    .A4(_0261_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _0961_ (.A1(net71),
    .A2(_0251_),
    .B(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _0962_ (.A1(_0450_),
    .A2(_0452_),
    .B1(_0454_),
    .B2(_0267_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _0963_ (.A1(net184),
    .A2(_0128_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0964_ (.I(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0965_ (.I0(net3),
    .I1(net185),
    .S(_0456_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0966_ (.I0(net4),
    .I1(net186),
    .S(_0456_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0967_ (.I0(net5),
    .I1(net187),
    .S(_0456_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0968_ (.I0(net6),
    .I1(net188),
    .S(_0456_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0969_ (.I0(net7),
    .I1(net189),
    .S(_0456_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0970_ (.I0(net8),
    .I1(net190),
    .S(_0456_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0971_ (.I0(net9),
    .I1(net191),
    .S(_0456_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0972_ (.I0(net10),
    .I1(net192),
    .S(_0456_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0973_ (.I0(net11),
    .I1(net193),
    .S(_0456_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0974_ (.I0(net12),
    .I1(net194),
    .S(_0456_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0975_ (.I(_0455_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0976_ (.I0(net13),
    .I1(net195),
    .S(_0457_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0977_ (.I0(net14),
    .I1(net196),
    .S(_0457_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0978_ (.I0(net15),
    .I1(net197),
    .S(_0457_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0979_ (.I0(net16),
    .I1(net198),
    .S(_0457_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0980_ (.I0(net17),
    .I1(net199),
    .S(_0457_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0981_ (.I0(net18),
    .I1(net200),
    .S(_0457_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0982_ (.I0(net19),
    .I1(net201),
    .S(_0457_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0983_ (.I0(net20),
    .I1(net202),
    .S(_0457_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0984_ (.I0(net21),
    .I1(net203),
    .S(_0457_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0985_ (.I0(net22),
    .I1(net204),
    .S(_0457_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _0986_ (.I(_0455_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0987_ (.I0(net23),
    .I1(net205),
    .S(_0458_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0988_ (.I0(net24),
    .I1(net206),
    .S(_0458_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0989_ (.I0(net25),
    .I1(net207),
    .S(_0458_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0990_ (.I0(net26),
    .I1(net208),
    .S(_0458_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0991_ (.I0(net27),
    .I1(net209),
    .S(_0458_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0992_ (.I0(net28),
    .I1(net210),
    .S(_0458_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0993_ (.I0(net29),
    .I1(net211),
    .S(_0458_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0994_ (.I0(net30),
    .I1(net212),
    .S(_0458_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0995_ (.I0(net31),
    .I1(net213),
    .S(_0458_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0996_ (.I0(net32),
    .I1(net214),
    .S(_0458_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0997_ (.I0(net33),
    .I1(net215),
    .S(_0455_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _0998_ (.I0(net34),
    .I1(net216),
    .S(_0455_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _0999_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _1000_ (.A1(net217),
    .A2(_0141_),
    .B1(_0459_),
    .B2(_0142_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1001_ (.I(_0460_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1002_ (.I0(net218),
    .I1(net37),
    .S(_0141_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1003_ (.I0(net219),
    .I1(net38),
    .S(_0141_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__addf_4 _1004_ (.A(_0464_),
    .B(_0465_),
    .CI(_0466_),
    .CO(_0467_),
    .S(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1005_ (.A(\burst_count[7] ),
    .B(_0469_),
    .CO(_0470_),
    .S(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1006_ (.A(\burst_count[6] ),
    .B(_0472_),
    .CO(_0473_),
    .S(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1007_ (.A(\burst_count[5] ),
    .B(_0475_),
    .CO(_0476_),
    .S(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1008_ (.A(_0478_),
    .B(_0479_),
    .CO(_0480_),
    .S(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1009_ (.A(\burst_count[4] ),
    .B(_0481_),
    .CO(_0482_),
    .S(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1010_ (.A(\burst_count[3] ),
    .B(_0484_),
    .CO(_0485_),
    .S(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1011_ (.A(_0487_),
    .B(_0488_),
    .CO(_0489_),
    .S(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1012_ (.A(\burst_count[2] ),
    .B(_0490_),
    .CO(_0491_),
    .S(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1013_ (.A(\burst_count[1] ),
    .B(\burst_total[0] ),
    .CO(_0493_),
    .S(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1014_ (.A(net111),
    .B(_0495_),
    .CO(_0496_),
    .S(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1015_ (.A(net122),
    .B(_0498_),
    .CO(_0499_),
    .S(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1016_ (.A(net133),
    .B(_0501_),
    .CO(_0502_),
    .S(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1017_ (.A(net136),
    .B(_0504_),
    .CO(_0505_),
    .S(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1018_ (.A(net137),
    .B(_0507_),
    .CO(_0508_),
    .S(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1019_ (.A(net138),
    .B(_0510_),
    .CO(_0511_),
    .S(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1020_ (.A(net139),
    .B(_0513_),
    .CO(_0514_),
    .S(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _1021_ (.A(net140),
    .B(_0516_),
    .CO(_0517_),
    .S(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _1022_ (.A(\burst_count[0] ),
    .B(\burst_count[1] ),
    .CO(_0519_),
    .S(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[0]$_DFFE_PN0P_  (.D(_0000_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[1]$_DFFE_PN0P_  (.D(_0001_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[2]$_DFFE_PN0P_  (.D(_0002_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[3]$_DFFE_PN0P_  (.D(_0003_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[4]$_DFFE_PN0P_  (.D(_0004_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[5]$_DFFE_PN0P_  (.D(_0005_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[6]$_DFFE_PN0P_  (.D(_0006_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_count[7]$_DFFE_PN0P_  (.D(_0007_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_count[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_total[0]$_DFFE_PN0P_  (.D(_0008_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_total[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_total[2]$_DFFE_PN0P_  (.D(_0009_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_total[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_total[3]$_DFFE_PN0P_  (.D(_0010_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_total[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \burst_total[4]$_DFFE_PN0P_  (.D(_0011_),
    .RN(net36),
    .CLK(net1),
    .Q(\burst_total[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hburst[0]$_DFFE_PN0P_  (.D(_0012_),
    .RN(net36),
    .CLK(net1),
    .Q(net143));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hburst[1]$_DFFE_PN0P_  (.D(_0013_),
    .RN(net36),
    .CLK(net1),
    .Q(net144));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hburst[2]$_DFFE_PN0P_  (.D(_0014_),
    .RN(net36),
    .CLK(net1),
    .Q(net145));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hbusreq$_DFFE_PN0P_  (.D(_0015_),
    .RN(net36),
    .CLK(net1),
    .Q(net146));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hsize[0]$_DFFE_PN0P_  (.D(_0016_),
    .RN(net36),
    .CLK(net1),
    .Q(net147));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hsize[1]$_DFFE_PN0P_  (.D(_0017_),
    .RN(net36),
    .CLK(net1),
    .Q(net148));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hsize[2]$_DFFE_PN0P_  (.D(_0018_),
    .RN(net36),
    .CLK(net1),
    .Q(net149));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \htrans[0]$_DFFE_PN0P_  (.D(_0019_),
    .RN(net36),
    .CLK(net1),
    .Q(net150));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \htrans[1]$_DFFE_PN0P_  (.D(_0020_),
    .RN(net36),
    .CLK(net1),
    .Q(net151));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[0]$_DFFE_PN0P_  (.D(_0021_),
    .RN(net36),
    .CLK(net1),
    .Q(net152));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[10]$_DFFE_PN0P_  (.D(_0022_),
    .RN(net36),
    .CLK(net1),
    .Q(net153));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[11]$_DFFE_PN0P_  (.D(_0023_),
    .RN(net36),
    .CLK(net1),
    .Q(net154));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[12]$_DFFE_PN0P_  (.D(_0024_),
    .RN(net36),
    .CLK(net1),
    .Q(net155));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[13]$_DFFE_PN0P_  (.D(_0025_),
    .RN(net36),
    .CLK(net1),
    .Q(net156));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[14]$_DFFE_PN0P_  (.D(_0026_),
    .RN(net36),
    .CLK(net1),
    .Q(net157));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[15]$_DFFE_PN0P_  (.D(_0027_),
    .RN(net36),
    .CLK(net1),
    .Q(net158));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[16]$_DFFE_PN0P_  (.D(_0028_),
    .RN(net36),
    .CLK(net1),
    .Q(net159));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[17]$_DFFE_PN0P_  (.D(_0029_),
    .RN(net36),
    .CLK(net1),
    .Q(net160));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[18]$_DFFE_PN0P_  (.D(_0030_),
    .RN(net36),
    .CLK(net1),
    .Q(net161));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[19]$_DFFE_PN0P_  (.D(_0031_),
    .RN(net36),
    .CLK(net1),
    .Q(net162));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[1]$_DFFE_PN0P_  (.D(_0032_),
    .RN(net36),
    .CLK(net1),
    .Q(net163));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[20]$_DFFE_PN0P_  (.D(_0033_),
    .RN(net36),
    .CLK(net1),
    .Q(net164));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[21]$_DFFE_PN0P_  (.D(_0034_),
    .RN(net36),
    .CLK(net1),
    .Q(net165));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[22]$_DFFE_PN0P_  (.D(_0035_),
    .RN(net36),
    .CLK(net1),
    .Q(net166));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[23]$_DFFE_PN0P_  (.D(_0036_),
    .RN(net36),
    .CLK(net1),
    .Q(net167));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[24]$_DFFE_PN0P_  (.D(_0037_),
    .RN(net36),
    .CLK(net1),
    .Q(net168));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[25]$_DFFE_PN0P_  (.D(_0038_),
    .RN(net36),
    .CLK(net1),
    .Q(net169));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[26]$_DFFE_PN0P_  (.D(_0039_),
    .RN(net36),
    .CLK(net1),
    .Q(net170));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[27]$_DFFE_PN0P_  (.D(_0040_),
    .RN(net36),
    .CLK(net1),
    .Q(net171));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[28]$_DFFE_PN0P_  (.D(_0041_),
    .RN(net36),
    .CLK(net1),
    .Q(net172));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[29]$_DFFE_PN0P_  (.D(_0042_),
    .RN(net36),
    .CLK(net1),
    .Q(net173));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[2]$_DFFE_PN0P_  (.D(_0043_),
    .RN(net36),
    .CLK(net1),
    .Q(net174));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[30]$_DFFE_PN0P_  (.D(_0044_),
    .RN(net36),
    .CLK(net1),
    .Q(net175));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[31]$_DFFE_PN0P_  (.D(_0045_),
    .RN(net36),
    .CLK(net1),
    .Q(net176));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[3]$_DFFE_PN0P_  (.D(_0046_),
    .RN(net36),
    .CLK(net1),
    .Q(net177));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[4]$_DFFE_PN0P_  (.D(_0047_),
    .RN(net36),
    .CLK(net1),
    .Q(net178));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[5]$_DFFE_PN0P_  (.D(_0048_),
    .RN(net36),
    .CLK(net1),
    .Q(net179));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[6]$_DFFE_PN0P_  (.D(_0049_),
    .RN(net36),
    .CLK(net1),
    .Q(net180));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[7]$_DFFE_PN0P_  (.D(_0050_),
    .RN(net36),
    .CLK(net1),
    .Q(net181));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[8]$_DFFE_PN0P_  (.D(_0051_),
    .RN(net36),
    .CLK(net1),
    .Q(net182));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwdata[9]$_DFFE_PN0P_  (.D(_0052_),
    .RN(net36),
    .CLK(net1),
    .Q(net183));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \hwrite$_DFFE_PN0P_  (.D(_0053_),
    .RN(net36),
    .CLK(net1),
    .Q(net184));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[0]$_DFFE_PN0P_  (.D(_0054_),
    .RN(net36),
    .CLK(net1),
    .Q(net111));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[10]$_DFFE_PN0P_  (.D(_0055_),
    .RN(net36),
    .CLK(net1),
    .Q(net112));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[11]$_DFFE_PN0P_  (.D(_0056_),
    .RN(net36),
    .CLK(net1),
    .Q(net113));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[12]$_DFFE_PN0P_  (.D(_0057_),
    .RN(net36),
    .CLK(net1),
    .Q(net114));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[13]$_DFFE_PN0P_  (.D(_0058_),
    .RN(net36),
    .CLK(net1),
    .Q(net115));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[14]$_DFFE_PN0P_  (.D(_0059_),
    .RN(net36),
    .CLK(net1),
    .Q(net116));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[15]$_DFFE_PN0P_  (.D(_0060_),
    .RN(net36),
    .CLK(net1),
    .Q(net117));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[16]$_DFFE_PN0P_  (.D(_0061_),
    .RN(net36),
    .CLK(net1),
    .Q(net118));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[17]$_DFFE_PN0P_  (.D(_0062_),
    .RN(net36),
    .CLK(net1),
    .Q(net119));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[18]$_DFFE_PN0P_  (.D(_0063_),
    .RN(net36),
    .CLK(net1),
    .Q(net120));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[19]$_DFFE_PN0P_  (.D(_0064_),
    .RN(net36),
    .CLK(net1),
    .Q(net121));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[1]$_DFFE_PN0P_  (.D(_0065_),
    .RN(net36),
    .CLK(net1),
    .Q(net122));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[20]$_DFFE_PN0P_  (.D(_0066_),
    .RN(net36),
    .CLK(net1),
    .Q(net123));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[21]$_DFFE_PN0P_  (.D(_0067_),
    .RN(net36),
    .CLK(net1),
    .Q(net124));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[22]$_DFFE_PN0P_  (.D(_0068_),
    .RN(net36),
    .CLK(net1),
    .Q(net125));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[23]$_DFFE_PN0P_  (.D(_0069_),
    .RN(net36),
    .CLK(net1),
    .Q(net126));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[24]$_DFFE_PN0P_  (.D(_0070_),
    .RN(net36),
    .CLK(net1),
    .Q(net127));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[25]$_DFFE_PN0P_  (.D(_0071_),
    .RN(net36),
    .CLK(net1),
    .Q(net128));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[26]$_DFFE_PN0P_  (.D(_0072_),
    .RN(net36),
    .CLK(net1),
    .Q(net129));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[27]$_DFFE_PN0P_  (.D(_0073_),
    .RN(net36),
    .CLK(net1),
    .Q(net130));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[28]$_DFFE_PN0P_  (.D(_0074_),
    .RN(net36),
    .CLK(net1),
    .Q(net131));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[29]$_DFFE_PN0P_  (.D(_0075_),
    .RN(net36),
    .CLK(net1),
    .Q(net132));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[2]$_DFFE_PN0P_  (.D(_0076_),
    .RN(net36),
    .CLK(net1),
    .Q(net133));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[30]$_DFFE_PN0P_  (.D(_0077_),
    .RN(net36),
    .CLK(net1),
    .Q(net134));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[31]$_DFFE_PN0P_  (.D(_0078_),
    .RN(net36),
    .CLK(net1),
    .Q(net135));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[3]$_DFFE_PN0P_  (.D(_0079_),
    .RN(net36),
    .CLK(net1),
    .Q(net136));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[4]$_DFFE_PN0P_  (.D(_0080_),
    .RN(net36),
    .CLK(net1),
    .Q(net137));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[5]$_DFFE_PN0P_  (.D(_0081_),
    .RN(net36),
    .CLK(net1),
    .Q(net138));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[6]$_DFFE_PN0P_  (.D(_0082_),
    .RN(net36),
    .CLK(net1),
    .Q(net139));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[7]$_DFFE_PN0P_  (.D(_0083_),
    .RN(net36),
    .CLK(net1),
    .Q(net140));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[8]$_DFFE_PN0P_  (.D(_0084_),
    .RN(net36),
    .CLK(net1),
    .Q(net141));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \next_addr[9]$_DFFE_PN0P_  (.D(_0085_),
    .RN(net36),
    .CLK(net1),
    .Q(net142));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[0]$_DFFE_PN0P_  (.D(_0086_),
    .RN(net36),
    .CLK(net1),
    .Q(net185));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[10]$_DFFE_PN0P_  (.D(_0087_),
    .RN(net36),
    .CLK(net1),
    .Q(net186));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[11]$_DFFE_PN0P_  (.D(_0088_),
    .RN(net36),
    .CLK(net1),
    .Q(net187));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[12]$_DFFE_PN0P_  (.D(_0089_),
    .RN(net36),
    .CLK(net1),
    .Q(net188));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[13]$_DFFE_PN0P_  (.D(_0090_),
    .RN(net36),
    .CLK(net1),
    .Q(net189));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[14]$_DFFE_PN0P_  (.D(_0091_),
    .RN(net36),
    .CLK(net1),
    .Q(net190));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[15]$_DFFE_PN0P_  (.D(_0092_),
    .RN(net36),
    .CLK(net1),
    .Q(net191));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[16]$_DFFE_PN0P_  (.D(_0093_),
    .RN(net36),
    .CLK(net1),
    .Q(net192));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[17]$_DFFE_PN0P_  (.D(_0094_),
    .RN(net36),
    .CLK(net1),
    .Q(net193));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[18]$_DFFE_PN0P_  (.D(_0095_),
    .RN(net36),
    .CLK(net1),
    .Q(net194));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[19]$_DFFE_PN0P_  (.D(_0096_),
    .RN(net36),
    .CLK(net1),
    .Q(net195));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[1]$_DFFE_PN0P_  (.D(_0097_),
    .RN(net36),
    .CLK(net1),
    .Q(net196));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[20]$_DFFE_PN0P_  (.D(_0098_),
    .RN(net36),
    .CLK(net1),
    .Q(net197));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[21]$_DFFE_PN0P_  (.D(_0099_),
    .RN(net36),
    .CLK(net1),
    .Q(net198));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[22]$_DFFE_PN0P_  (.D(_0100_),
    .RN(net36),
    .CLK(net1),
    .Q(net199));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[23]$_DFFE_PN0P_  (.D(_0101_),
    .RN(net36),
    .CLK(net1),
    .Q(net200));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[24]$_DFFE_PN0P_  (.D(_0102_),
    .RN(net36),
    .CLK(net1),
    .Q(net201));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[25]$_DFFE_PN0P_  (.D(_0103_),
    .RN(net36),
    .CLK(net1),
    .Q(net202));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[26]$_DFFE_PN0P_  (.D(_0104_),
    .RN(net36),
    .CLK(net1),
    .Q(net203));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[27]$_DFFE_PN0P_  (.D(_0105_),
    .RN(net36),
    .CLK(net1),
    .Q(net204));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[28]$_DFFE_PN0P_  (.D(_0106_),
    .RN(net36),
    .CLK(net1),
    .Q(net205));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[29]$_DFFE_PN0P_  (.D(_0107_),
    .RN(net36),
    .CLK(net1),
    .Q(net206));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[2]$_DFFE_PN0P_  (.D(_0108_),
    .RN(net36),
    .CLK(net1),
    .Q(net207));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[30]$_DFFE_PN0P_  (.D(_0109_),
    .RN(net36),
    .CLK(net1),
    .Q(net208));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[31]$_DFFE_PN0P_  (.D(_0110_),
    .RN(net36),
    .CLK(net1),
    .Q(net209));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[3]$_DFFE_PN0P_  (.D(_0111_),
    .RN(net36),
    .CLK(net1),
    .Q(net210));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[4]$_DFFE_PN0P_  (.D(_0112_),
    .RN(net36),
    .CLK(net1),
    .Q(net211));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[5]$_DFFE_PN0P_  (.D(_0113_),
    .RN(net36),
    .CLK(net1),
    .Q(net212));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[6]$_DFFE_PN0P_  (.D(_0114_),
    .RN(net36),
    .CLK(net1),
    .Q(net213));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[7]$_DFFE_PN0P_  (.D(_0115_),
    .RN(net36),
    .CLK(net1),
    .Q(net214));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[8]$_DFFE_PN0P_  (.D(_0116_),
    .RN(net36),
    .CLK(net1),
    .Q(net215));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \read_data[9]$_DFFE_PN0P_  (.D(_0117_),
    .RN(net36),
    .CLK(net1),
    .Q(net216));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFF_PN0_  (.D(_0461_),
    .RN(net36),
    .CLK(net1),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \state[1]$_DFF_PN0_  (.D(_0462_),
    .RN(net36),
    .CLK(net1),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[2]$_DFF_PN0_  (.D(_0463_),
    .RN(net36),
    .CLK(net1),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \trans_done$_DFFE_PN0P_  (.D(_0118_),
    .RN(net36),
    .CLK(net1),
    .Q(net217));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \trans_resp[0]$_DFFE_PN0P_  (.D(_0119_),
    .RN(net36),
    .CLK(net1),
    .Q(net218));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \trans_resp[1]$_DFFE_PN0P_  (.D(_0120_),
    .RN(net36),
    .CLK(net1),
    .Q(net219));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_106 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_107 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_108 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_109 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_110 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_111 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_112 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_113 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_114 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_115 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_116 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_117 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_118 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_119 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_120 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_121 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_122 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_123 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_124 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_125 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_126 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_127 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_128 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_160 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input1 (.I(hclk),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(hgrant),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(hrdata[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(hrdata[10]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(hrdata[11]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(hrdata[12]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(hrdata[13]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(hrdata[14]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(hrdata[15]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(hrdata[16]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(hrdata[17]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input12 (.I(hrdata[18]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(hrdata[19]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(hrdata[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(hrdata[20]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(hrdata[21]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(hrdata[22]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(hrdata[23]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(hrdata[24]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(hrdata[25]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(hrdata[26]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(hrdata[27]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input23 (.I(hrdata[28]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(hrdata[29]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(hrdata[2]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(hrdata[30]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(hrdata[31]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(hrdata[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(hrdata[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(hrdata[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(hrdata[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(hrdata[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input33 (.I(hrdata[8]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(hrdata[9]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input35 (.I(hready),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input36 (.I(hreset),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(hresp[0]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(hresp[1]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input39 (.I(start_trans),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input40 (.I(trans_addr[0]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(trans_addr[10]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(trans_addr[11]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(trans_addr[12]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input44 (.I(trans_addr[13]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(trans_addr[14]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(trans_addr[15]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(trans_addr[16]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(trans_addr[17]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(trans_addr[18]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input50 (.I(trans_addr[19]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(trans_addr[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(trans_addr[20]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(trans_addr[21]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(trans_addr[22]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input55 (.I(trans_addr[23]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(trans_addr[24]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(trans_addr[25]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(trans_addr[26]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(trans_addr[27]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input60 (.I(trans_addr[28]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input61 (.I(trans_addr[29]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(trans_addr[2]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(trans_addr[30]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(trans_addr[31]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input65 (.I(trans_addr[3]),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input66 (.I(trans_addr[4]),
    .Z(net66));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input67 (.I(trans_addr[5]),
    .Z(net67));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input68 (.I(trans_addr[6]),
    .Z(net68));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input69 (.I(trans_addr[7]),
    .Z(net69));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input70 (.I(trans_addr[8]),
    .Z(net70));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input71 (.I(trans_addr[9]),
    .Z(net71));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input72 (.I(trans_burst[0]),
    .Z(net72));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input73 (.I(trans_burst[1]),
    .Z(net73));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input74 (.I(trans_burst[2]),
    .Z(net74));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input75 (.I(trans_size[0]),
    .Z(net75));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input76 (.I(trans_size[1]),
    .Z(net76));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input77 (.I(trans_size[2]),
    .Z(net77));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input78 (.I(trans_write),
    .Z(net78));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input79 (.I(write_data[0]),
    .Z(net79));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input80 (.I(write_data[10]),
    .Z(net80));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input81 (.I(write_data[11]),
    .Z(net81));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input82 (.I(write_data[12]),
    .Z(net82));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input83 (.I(write_data[13]),
    .Z(net83));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input84 (.I(write_data[14]),
    .Z(net84));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input85 (.I(write_data[15]),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input86 (.I(write_data[16]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input87 (.I(write_data[17]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input88 (.I(write_data[18]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input89 (.I(write_data[19]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input90 (.I(write_data[1]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input91 (.I(write_data[20]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input92 (.I(write_data[21]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input93 (.I(write_data[22]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input94 (.I(write_data[23]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input95 (.I(write_data[24]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input96 (.I(write_data[25]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input97 (.I(write_data[26]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input98 (.I(write_data[27]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input99 (.I(write_data[28]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input100 (.I(write_data[29]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input101 (.I(write_data[2]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input102 (.I(write_data[30]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input103 (.I(write_data[31]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input104 (.I(write_data[3]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input105 (.I(write_data[4]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input106 (.I(write_data[5]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input107 (.I(write_data[6]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input108 (.I(write_data[7]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input109 (.I(write_data[8]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input110 (.I(write_data[9]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output111 (.I(net111),
    .Z(haddr[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output112 (.I(net112),
    .Z(haddr[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output113 (.I(net113),
    .Z(haddr[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output114 (.I(net114),
    .Z(haddr[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output115 (.I(net115),
    .Z(haddr[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output116 (.I(net116),
    .Z(haddr[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output117 (.I(net117),
    .Z(haddr[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output118 (.I(net118),
    .Z(haddr[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output119 (.I(net119),
    .Z(haddr[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output120 (.I(net120),
    .Z(haddr[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output121 (.I(net121),
    .Z(haddr[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output122 (.I(net122),
    .Z(haddr[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output123 (.I(net123),
    .Z(haddr[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output124 (.I(net124),
    .Z(haddr[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output125 (.I(net125),
    .Z(haddr[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output126 (.I(net126),
    .Z(haddr[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output127 (.I(net127),
    .Z(haddr[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output128 (.I(net128),
    .Z(haddr[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output129 (.I(net129),
    .Z(haddr[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output130 (.I(net130),
    .Z(haddr[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output131 (.I(net131),
    .Z(haddr[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output132 (.I(net132),
    .Z(haddr[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output133 (.I(net133),
    .Z(haddr[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output134 (.I(net134),
    .Z(haddr[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output135 (.I(net135),
    .Z(haddr[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output136 (.I(net136),
    .Z(haddr[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output137 (.I(net137),
    .Z(haddr[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output138 (.I(net138),
    .Z(haddr[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output139 (.I(net139),
    .Z(haddr[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output140 (.I(net140),
    .Z(haddr[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output141 (.I(net141),
    .Z(haddr[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output142 (.I(net142),
    .Z(haddr[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output143 (.I(net143),
    .Z(hburst[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output144 (.I(net144),
    .Z(hburst[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output145 (.I(net145),
    .Z(hburst[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output146 (.I(net146),
    .Z(hbusreq));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output147 (.I(net147),
    .Z(hsize[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output148 (.I(net148),
    .Z(hsize[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output149 (.I(net149),
    .Z(hsize[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output150 (.I(net150),
    .Z(htrans[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output151 (.I(net151),
    .Z(htrans[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output152 (.I(net152),
    .Z(hwdata[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output153 (.I(net153),
    .Z(hwdata[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output154 (.I(net154),
    .Z(hwdata[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output155 (.I(net155),
    .Z(hwdata[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output156 (.I(net156),
    .Z(hwdata[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output157 (.I(net157),
    .Z(hwdata[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output158 (.I(net158),
    .Z(hwdata[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output159 (.I(net159),
    .Z(hwdata[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output160 (.I(net160),
    .Z(hwdata[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output161 (.I(net161),
    .Z(hwdata[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output162 (.I(net162),
    .Z(hwdata[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output163 (.I(net163),
    .Z(hwdata[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output164 (.I(net164),
    .Z(hwdata[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output165 (.I(net165),
    .Z(hwdata[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output166 (.I(net166),
    .Z(hwdata[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output167 (.I(net167),
    .Z(hwdata[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output168 (.I(net168),
    .Z(hwdata[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output169 (.I(net169),
    .Z(hwdata[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output170 (.I(net170),
    .Z(hwdata[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output171 (.I(net171),
    .Z(hwdata[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output172 (.I(net172),
    .Z(hwdata[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output173 (.I(net173),
    .Z(hwdata[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output174 (.I(net174),
    .Z(hwdata[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output175 (.I(net175),
    .Z(hwdata[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output176 (.I(net176),
    .Z(hwdata[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output177 (.I(net177),
    .Z(hwdata[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output178 (.I(net178),
    .Z(hwdata[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output179 (.I(net179),
    .Z(hwdata[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output180 (.I(net180),
    .Z(hwdata[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output181 (.I(net181),
    .Z(hwdata[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output182 (.I(net182),
    .Z(hwdata[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output183 (.I(net183),
    .Z(hwdata[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output184 (.I(net184),
    .Z(hwrite));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output185 (.I(net185),
    .Z(read_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output186 (.I(net186),
    .Z(read_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output187 (.I(net187),
    .Z(read_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output188 (.I(net188),
    .Z(read_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output189 (.I(net189),
    .Z(read_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output190 (.I(net190),
    .Z(read_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output191 (.I(net191),
    .Z(read_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output192 (.I(net192),
    .Z(read_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output193 (.I(net193),
    .Z(read_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output194 (.I(net194),
    .Z(read_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output195 (.I(net195),
    .Z(read_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output196 (.I(net196),
    .Z(read_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output197 (.I(net197),
    .Z(read_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output198 (.I(net198),
    .Z(read_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output199 (.I(net199),
    .Z(read_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output200 (.I(net200),
    .Z(read_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output201 (.I(net201),
    .Z(read_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output202 (.I(net202),
    .Z(read_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output203 (.I(net203),
    .Z(read_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output204 (.I(net204),
    .Z(read_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output205 (.I(net205),
    .Z(read_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output206 (.I(net206),
    .Z(read_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output207 (.I(net207),
    .Z(read_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output208 (.I(net208),
    .Z(read_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output209 (.I(net209),
    .Z(read_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output210 (.I(net210),
    .Z(read_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output211 (.I(net211),
    .Z(read_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output212 (.I(net212),
    .Z(read_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output213 (.I(net213),
    .Z(read_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output214 (.I(net214),
    .Z(read_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output215 (.I(net215),
    .Z(read_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output216 (.I(net216),
    .Z(read_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output217 (.I(net217),
    .Z(trans_done));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output218 (.I(net218),
    .Z(trans_resp[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output219 (.I(net219),
    .Z(trans_resp[1]));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_397 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_68 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_59 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_12 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_43 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_19 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_486 ();
endmodule
