module network_interface (clk,
    mem_read,
    mem_ready,
    mem_write,
    router_in_ready,
    router_in_valid,
    router_out_ready,
    router_out_valid,
    rst_n,
    dest_id,
    mem_addr,
    mem_rdata,
    mem_wdata,
    msg_type,
    router_in_data,
    router_out_data);
 input clk;
 input mem_read;
 output mem_ready;
 input mem_write;
 input router_in_ready;
 output router_in_valid;
 output router_out_ready;
 input router_out_valid;
 input rst_n;
 input [7:0] dest_id;
 input [31:0] mem_addr;
 output [31:0] mem_rdata;
 input [31:0] mem_wdata;
 input [2:0] msg_type;
 output [31:0] router_in_data;
 input [31:0] router_out_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire first_write_done;
 wire is_write_op;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 BUF_X2 _374_ (.A(rst_n),
    .Z(_073_));
 BUF_X2 _375_ (.A(_073_),
    .Z(_074_));
 BUF_X2 _376_ (.A(_074_),
    .Z(_075_));
 BUF_X4 _377_ (.A(\state[2] ),
    .Z(_076_));
 BUF_X4 _378_ (.A(_076_),
    .Z(_077_));
 INV_X4 _379_ (.A(_077_),
    .ZN(_078_));
 BUF_X4 _380_ (.A(_078_),
    .Z(_079_));
 NAND2_X1 _381_ (.A1(net165),
    .A2(net66),
    .ZN(_080_));
 BUF_X4 _382_ (.A(\state[1] ),
    .Z(_081_));
 NAND3_X2 _383_ (.A1(net165),
    .A2(net66),
    .A3(is_write_op),
    .ZN(_082_));
 NAND2_X1 _384_ (.A1(_081_),
    .A2(_082_),
    .ZN(_083_));
 OAI22_X1 _385_ (.A1(_079_),
    .A2(_080_),
    .B1(_083_),
    .B2(net99),
    .ZN(_084_));
 AND2_X1 _386_ (.A1(_075_),
    .A2(_084_),
    .ZN(_002_));
 INV_X1 _387_ (.A(_073_),
    .ZN(_085_));
 BUF_X4 _388_ (.A(_085_),
    .Z(_086_));
 CLKBUF_X3 _389_ (.A(_086_),
    .Z(_087_));
 CLKBUF_X3 _390_ (.A(_076_),
    .Z(_088_));
 CLKBUF_X3 _391_ (.A(_088_),
    .Z(_089_));
 NAND2_X1 _392_ (.A1(_089_),
    .A2(_080_),
    .ZN(_090_));
 BUF_X4 _393_ (.A(\state[0] ),
    .Z(_091_));
 BUF_X4 _394_ (.A(mem_write),
    .Z(_092_));
 OAI21_X1 _395_ (.A(_091_),
    .B1(_092_),
    .B2(net30),
    .ZN(_093_));
 AOI21_X1 _396_ (.A(_087_),
    .B1(_090_),
    .B2(_093_),
    .ZN(_003_));
 AND3_X1 _397_ (.A1(net165),
    .A2(net66),
    .A3(is_write_op),
    .ZN(_094_));
 NAND2_X1 _398_ (.A1(_081_),
    .A2(_094_),
    .ZN(_095_));
 INV_X2 _399_ (.A(_091_),
    .ZN(_096_));
 OR3_X2 _400_ (.A1(_096_),
    .A2(_092_),
    .A3(net30),
    .ZN(_097_));
 NOR2_X1 _401_ (.A1(_087_),
    .A2(\state[3] ),
    .ZN(_098_));
 NAND3_X1 _402_ (.A1(_095_),
    .A2(_097_),
    .A3(_098_),
    .ZN(_001_));
 NAND3_X4 _403_ (.A1(net99),
    .A2(_081_),
    .A3(_082_),
    .ZN(_099_));
 BUF_X8 _404_ (.A(_099_),
    .Z(_100_));
 NOR2_X1 _405_ (.A1(_087_),
    .A2(_100_),
    .ZN(_000_));
 MUX2_X1 _406_ (.A(net67),
    .B(net100),
    .S(_100_),
    .Z(_101_));
 AND2_X1 _407_ (.A1(_075_),
    .A2(_101_),
    .ZN(_005_));
 MUX2_X1 _408_ (.A(net68),
    .B(net101),
    .S(_100_),
    .Z(_102_));
 AND2_X1 _409_ (.A1(_075_),
    .A2(_102_),
    .ZN(_006_));
 MUX2_X1 _410_ (.A(net69),
    .B(net102),
    .S(_100_),
    .Z(_103_));
 AND2_X1 _411_ (.A1(_075_),
    .A2(_103_),
    .ZN(_007_));
 MUX2_X1 _412_ (.A(net70),
    .B(net103),
    .S(_100_),
    .Z(_104_));
 AND2_X1 _413_ (.A1(_075_),
    .A2(_104_),
    .ZN(_008_));
 MUX2_X1 _414_ (.A(net71),
    .B(net104),
    .S(_100_),
    .Z(_105_));
 AND2_X1 _415_ (.A1(_075_),
    .A2(_105_),
    .ZN(_009_));
 MUX2_X1 _416_ (.A(net72),
    .B(net105),
    .S(_100_),
    .Z(_106_));
 AND2_X1 _417_ (.A1(_075_),
    .A2(_106_),
    .ZN(_010_));
 MUX2_X1 _418_ (.A(net73),
    .B(net106),
    .S(_100_),
    .Z(_107_));
 AND2_X1 _419_ (.A1(_075_),
    .A2(_107_),
    .ZN(_011_));
 MUX2_X1 _420_ (.A(net74),
    .B(net107),
    .S(_100_),
    .Z(_108_));
 AND2_X1 _421_ (.A1(_075_),
    .A2(_108_),
    .ZN(_012_));
 MUX2_X1 _422_ (.A(net75),
    .B(net108),
    .S(_100_),
    .Z(_109_));
 AND2_X1 _423_ (.A1(_075_),
    .A2(_109_),
    .ZN(_013_));
 CLKBUF_X2 _424_ (.A(_074_),
    .Z(_110_));
 BUF_X8 _425_ (.A(_099_),
    .Z(_111_));
 MUX2_X1 _426_ (.A(net76),
    .B(net109),
    .S(_111_),
    .Z(_112_));
 AND2_X1 _427_ (.A1(_110_),
    .A2(_112_),
    .ZN(_014_));
 MUX2_X1 _428_ (.A(net77),
    .B(net110),
    .S(_111_),
    .Z(_113_));
 AND2_X1 _429_ (.A1(_110_),
    .A2(_113_),
    .ZN(_015_));
 MUX2_X1 _430_ (.A(net78),
    .B(net111),
    .S(_111_),
    .Z(_114_));
 AND2_X1 _431_ (.A1(_110_),
    .A2(_114_),
    .ZN(_016_));
 MUX2_X1 _432_ (.A(net79),
    .B(net112),
    .S(_111_),
    .Z(_115_));
 AND2_X1 _433_ (.A1(_110_),
    .A2(_115_),
    .ZN(_017_));
 MUX2_X1 _434_ (.A(net80),
    .B(net113),
    .S(_111_),
    .Z(_116_));
 AND2_X1 _435_ (.A1(_110_),
    .A2(_116_),
    .ZN(_018_));
 MUX2_X1 _436_ (.A(net81),
    .B(net114),
    .S(_111_),
    .Z(_117_));
 AND2_X1 _437_ (.A1(_110_),
    .A2(_117_),
    .ZN(_019_));
 MUX2_X1 _438_ (.A(net82),
    .B(net115),
    .S(_111_),
    .Z(_118_));
 AND2_X1 _439_ (.A1(_110_),
    .A2(_118_),
    .ZN(_020_));
 MUX2_X1 _440_ (.A(net83),
    .B(net116),
    .S(_111_),
    .Z(_119_));
 AND2_X1 _441_ (.A1(_110_),
    .A2(_119_),
    .ZN(_021_));
 MUX2_X1 _442_ (.A(net84),
    .B(net117),
    .S(_111_),
    .Z(_120_));
 AND2_X1 _443_ (.A1(_110_),
    .A2(_120_),
    .ZN(_022_));
 MUX2_X1 _444_ (.A(net85),
    .B(net118),
    .S(_111_),
    .Z(_121_));
 AND2_X1 _445_ (.A1(_110_),
    .A2(_121_),
    .ZN(_023_));
 CLKBUF_X2 _446_ (.A(_074_),
    .Z(_122_));
 BUF_X8 _447_ (.A(_099_),
    .Z(_123_));
 MUX2_X1 _448_ (.A(net86),
    .B(net119),
    .S(_123_),
    .Z(_124_));
 AND2_X1 _449_ (.A1(_122_),
    .A2(_124_),
    .ZN(_024_));
 MUX2_X1 _450_ (.A(net87),
    .B(net120),
    .S(_123_),
    .Z(_125_));
 AND2_X1 _451_ (.A1(_122_),
    .A2(_125_),
    .ZN(_025_));
 MUX2_X1 _452_ (.A(net88),
    .B(net121),
    .S(_123_),
    .Z(_126_));
 AND2_X1 _453_ (.A1(_122_),
    .A2(_126_),
    .ZN(_026_));
 MUX2_X1 _454_ (.A(net89),
    .B(net122),
    .S(_123_),
    .Z(_127_));
 AND2_X1 _455_ (.A1(_122_),
    .A2(_127_),
    .ZN(_027_));
 MUX2_X1 _456_ (.A(net90),
    .B(net123),
    .S(_123_),
    .Z(_128_));
 AND2_X1 _457_ (.A1(_122_),
    .A2(_128_),
    .ZN(_028_));
 MUX2_X1 _458_ (.A(net91),
    .B(net124),
    .S(_123_),
    .Z(_129_));
 AND2_X1 _459_ (.A1(_122_),
    .A2(_129_),
    .ZN(_029_));
 MUX2_X1 _460_ (.A(net92),
    .B(net125),
    .S(_123_),
    .Z(_130_));
 AND2_X1 _461_ (.A1(_122_),
    .A2(_130_),
    .ZN(_030_));
 MUX2_X1 _462_ (.A(net93),
    .B(net126),
    .S(_123_),
    .Z(_131_));
 AND2_X1 _463_ (.A1(_122_),
    .A2(_131_),
    .ZN(_031_));
 MUX2_X1 _464_ (.A(net94),
    .B(net127),
    .S(_123_),
    .Z(_132_));
 AND2_X1 _465_ (.A1(_122_),
    .A2(_132_),
    .ZN(_032_));
 MUX2_X1 _466_ (.A(net95),
    .B(net128),
    .S(_123_),
    .Z(_133_));
 AND2_X1 _467_ (.A1(_122_),
    .A2(_133_),
    .ZN(_033_));
 MUX2_X1 _468_ (.A(net96),
    .B(net129),
    .S(_099_),
    .Z(_134_));
 AND2_X1 _469_ (.A1(_074_),
    .A2(_134_),
    .ZN(_034_));
 MUX2_X1 _470_ (.A(net97),
    .B(net130),
    .S(_099_),
    .Z(_135_));
 AND2_X1 _471_ (.A1(_074_),
    .A2(_135_),
    .ZN(_035_));
 MUX2_X1 _472_ (.A(net98),
    .B(net131),
    .S(_099_),
    .Z(_136_));
 AND2_X1 _473_ (.A1(_074_),
    .A2(_136_),
    .ZN(_036_));
 NOR2_X1 _474_ (.A1(\state[3] ),
    .A2(_091_),
    .ZN(_137_));
 NAND3_X1 _475_ (.A1(_073_),
    .A2(_081_),
    .A3(_137_),
    .ZN(_138_));
 BUF_X2 _476_ (.A(_073_),
    .Z(_139_));
 NAND3_X1 _477_ (.A1(_139_),
    .A2(_081_),
    .A3(net132),
    .ZN(_140_));
 NOR2_X1 _478_ (.A1(net99),
    .A2(_094_),
    .ZN(_141_));
 MUX2_X1 _479_ (.A(_138_),
    .B(_140_),
    .S(_141_),
    .Z(_142_));
 NAND3_X1 _480_ (.A1(_074_),
    .A2(net132),
    .A3(_137_),
    .ZN(_143_));
 NAND2_X1 _481_ (.A1(_142_),
    .A2(_143_),
    .ZN(_037_));
 INV_X1 _482_ (.A(net31),
    .ZN(_144_));
 INV_X4 _483_ (.A(_092_),
    .ZN(_145_));
 BUF_X1 _484_ (.A(first_write_done),
    .Z(_146_));
 OR2_X1 _485_ (.A1(_145_),
    .A2(_146_),
    .ZN(_147_));
 BUF_X4 _486_ (.A(_147_),
    .Z(_148_));
 BUF_X4 _487_ (.A(_076_),
    .Z(_149_));
 NOR2_X1 _488_ (.A1(_149_),
    .A2(net9),
    .ZN(_150_));
 AOI221_X1 _489_ (.A(_086_),
    .B1(_088_),
    .B2(_144_),
    .C1(_148_),
    .C2(_150_),
    .ZN(_151_));
 AND2_X1 _490_ (.A1(_074_),
    .A2(net133),
    .ZN(_152_));
 MUX2_X1 _491_ (.A(_091_),
    .B(_094_),
    .S(_076_),
    .Z(_153_));
 NAND2_X4 _492_ (.A1(_097_),
    .A2(_153_),
    .ZN(_154_));
 BUF_X8 _493_ (.A(_154_),
    .Z(_155_));
 MUX2_X1 _494_ (.A(_151_),
    .B(_152_),
    .S(_155_),
    .Z(_038_));
 INV_X1 _495_ (.A(net32),
    .ZN(_156_));
 NOR2_X1 _496_ (.A1(_149_),
    .A2(net10),
    .ZN(_157_));
 AOI221_X1 _497_ (.A(_086_),
    .B1(_088_),
    .B2(_156_),
    .C1(_148_),
    .C2(_157_),
    .ZN(_158_));
 AND2_X1 _498_ (.A1(_074_),
    .A2(net134),
    .ZN(_159_));
 MUX2_X1 _499_ (.A(_158_),
    .B(_159_),
    .S(_155_),
    .Z(_039_));
 NAND2_X1 _500_ (.A1(_089_),
    .A2(net33),
    .ZN(_160_));
 BUF_X4 _501_ (.A(_146_),
    .Z(_161_));
 BUF_X4 _502_ (.A(_161_),
    .Z(_162_));
 BUF_X4 _503_ (.A(_145_),
    .Z(_163_));
 OAI211_X2 _504_ (.A(_079_),
    .B(net11),
    .C1(_162_),
    .C2(_163_),
    .ZN(_164_));
 AOI21_X1 _505_ (.A(_087_),
    .B1(_160_),
    .B2(_164_),
    .ZN(_165_));
 AND2_X1 _506_ (.A1(_074_),
    .A2(net135),
    .ZN(_166_));
 MUX2_X1 _507_ (.A(_165_),
    .B(_166_),
    .S(_155_),
    .Z(_040_));
 NAND2_X1 _508_ (.A1(_089_),
    .A2(net34),
    .ZN(_167_));
 OAI211_X2 _509_ (.A(_079_),
    .B(net12),
    .C1(_162_),
    .C2(_163_),
    .ZN(_168_));
 AOI21_X1 _510_ (.A(_087_),
    .B1(_167_),
    .B2(_168_),
    .ZN(_169_));
 BUF_X2 _511_ (.A(_073_),
    .Z(_170_));
 AND2_X1 _512_ (.A1(_170_),
    .A2(net136),
    .ZN(_171_));
 MUX2_X1 _513_ (.A(_169_),
    .B(_171_),
    .S(_155_),
    .Z(_041_));
 NAND2_X1 _514_ (.A1(_089_),
    .A2(net35),
    .ZN(_172_));
 OAI211_X2 _515_ (.A(_079_),
    .B(net13),
    .C1(_162_),
    .C2(_163_),
    .ZN(_173_));
 AOI21_X1 _516_ (.A(_087_),
    .B1(_172_),
    .B2(_173_),
    .ZN(_174_));
 AND2_X1 _517_ (.A1(_170_),
    .A2(net137),
    .ZN(_175_));
 MUX2_X1 _518_ (.A(_174_),
    .B(_175_),
    .S(_155_),
    .Z(_042_));
 INV_X1 _519_ (.A(net36),
    .ZN(_176_));
 NOR2_X1 _520_ (.A1(_149_),
    .A2(net14),
    .ZN(_177_));
 AOI221_X1 _521_ (.A(_086_),
    .B1(_088_),
    .B2(_176_),
    .C1(_148_),
    .C2(_177_),
    .ZN(_178_));
 AND2_X1 _522_ (.A1(_170_),
    .A2(net138),
    .ZN(_179_));
 MUX2_X1 _523_ (.A(_178_),
    .B(_179_),
    .S(_155_),
    .Z(_043_));
 CLKBUF_X3 _524_ (.A(_086_),
    .Z(_180_));
 NAND2_X1 _525_ (.A1(_089_),
    .A2(net37),
    .ZN(_181_));
 OAI211_X2 _526_ (.A(_079_),
    .B(net15),
    .C1(_162_),
    .C2(_163_),
    .ZN(_182_));
 AOI21_X1 _527_ (.A(_180_),
    .B1(_181_),
    .B2(_182_),
    .ZN(_183_));
 AND2_X1 _528_ (.A1(_170_),
    .A2(net139),
    .ZN(_184_));
 MUX2_X1 _529_ (.A(_183_),
    .B(_184_),
    .S(_155_),
    .Z(_044_));
 CLKBUF_X3 _530_ (.A(_085_),
    .Z(_185_));
 INV_X1 _531_ (.A(net38),
    .ZN(_186_));
 NOR2_X1 _532_ (.A1(_149_),
    .A2(net16),
    .ZN(_187_));
 AOI221_X1 _533_ (.A(_185_),
    .B1(_088_),
    .B2(_186_),
    .C1(_148_),
    .C2(_187_),
    .ZN(_188_));
 AND2_X1 _534_ (.A1(_170_),
    .A2(net140),
    .ZN(_189_));
 MUX2_X1 _535_ (.A(_188_),
    .B(_189_),
    .S(_155_),
    .Z(_045_));
 INV_X1 _536_ (.A(net39),
    .ZN(_190_));
 NOR2_X1 _537_ (.A1(_149_),
    .A2(net17),
    .ZN(_191_));
 AOI221_X1 _538_ (.A(_185_),
    .B1(_088_),
    .B2(_190_),
    .C1(_148_),
    .C2(_191_),
    .ZN(_192_));
 AND2_X1 _539_ (.A1(_170_),
    .A2(net141),
    .ZN(_193_));
 MUX2_X1 _540_ (.A(_192_),
    .B(_193_),
    .S(_155_),
    .Z(_046_));
 NAND2_X1 _541_ (.A1(_089_),
    .A2(net40),
    .ZN(_194_));
 OAI211_X2 _542_ (.A(_079_),
    .B(net18),
    .C1(_162_),
    .C2(_163_),
    .ZN(_195_));
 AOI21_X1 _543_ (.A(_180_),
    .B1(_194_),
    .B2(_195_),
    .ZN(_196_));
 AND2_X1 _544_ (.A1(_170_),
    .A2(net142),
    .ZN(_197_));
 MUX2_X1 _545_ (.A(_196_),
    .B(_197_),
    .S(_155_),
    .Z(_047_));
 INV_X1 _546_ (.A(net41),
    .ZN(_198_));
 NOR2_X1 _547_ (.A1(_077_),
    .A2(net19),
    .ZN(_199_));
 AOI221_X1 _548_ (.A(_185_),
    .B1(_088_),
    .B2(_198_),
    .C1(_148_),
    .C2(_199_),
    .ZN(_200_));
 AND2_X1 _549_ (.A1(_170_),
    .A2(net143),
    .ZN(_201_));
 BUF_X8 _550_ (.A(_154_),
    .Z(_202_));
 MUX2_X1 _551_ (.A(_200_),
    .B(_201_),
    .S(_202_),
    .Z(_048_));
 INV_X1 _552_ (.A(net42),
    .ZN(_203_));
 NOR2_X1 _553_ (.A1(_077_),
    .A2(net20),
    .ZN(_204_));
 AOI221_X1 _554_ (.A(_185_),
    .B1(_088_),
    .B2(_203_),
    .C1(_148_),
    .C2(_204_),
    .ZN(_205_));
 AND2_X1 _555_ (.A1(_170_),
    .A2(net144),
    .ZN(_206_));
 MUX2_X1 _556_ (.A(_205_),
    .B(_206_),
    .S(_202_),
    .Z(_049_));
 NOR2_X1 _557_ (.A1(_079_),
    .A2(net43),
    .ZN(_207_));
 CLKBUF_X3 _558_ (.A(_149_),
    .Z(_208_));
 NOR3_X1 _559_ (.A1(_208_),
    .A2(_092_),
    .A3(net21),
    .ZN(_209_));
 NOR3_X1 _560_ (.A1(_087_),
    .A2(_207_),
    .A3(_209_),
    .ZN(_210_));
 AND2_X1 _561_ (.A1(_170_),
    .A2(net145),
    .ZN(_211_));
 MUX2_X1 _562_ (.A(_210_),
    .B(_211_),
    .S(_202_),
    .Z(_050_));
 INV_X1 _563_ (.A(net44),
    .ZN(_212_));
 NOR2_X1 _564_ (.A1(_077_),
    .A2(net63),
    .ZN(_213_));
 AOI221_X1 _565_ (.A(_185_),
    .B1(_088_),
    .B2(_212_),
    .C1(_148_),
    .C2(_213_),
    .ZN(_214_));
 BUF_X2 _566_ (.A(_073_),
    .Z(_215_));
 AND2_X1 _567_ (.A1(_215_),
    .A2(net146),
    .ZN(_216_));
 MUX2_X1 _568_ (.A(_214_),
    .B(_216_),
    .S(_202_),
    .Z(_051_));
 NAND2_X1 _569_ (.A1(_089_),
    .A2(net45),
    .ZN(_217_));
 OAI211_X2 _570_ (.A(_079_),
    .B(net64),
    .C1(_162_),
    .C2(_163_),
    .ZN(_218_));
 AOI21_X1 _571_ (.A(_180_),
    .B1(_217_),
    .B2(_218_),
    .ZN(_219_));
 AND2_X1 _572_ (.A1(_215_),
    .A2(net147),
    .ZN(_220_));
 MUX2_X1 _573_ (.A(_219_),
    .B(_220_),
    .S(_202_),
    .Z(_052_));
 NAND2_X1 _574_ (.A1(_089_),
    .A2(net46),
    .ZN(_221_));
 OAI211_X2 _575_ (.A(_079_),
    .B(net65),
    .C1(_162_),
    .C2(_163_),
    .ZN(_222_));
 AOI21_X1 _576_ (.A(_180_),
    .B1(_221_),
    .B2(_222_),
    .ZN(_223_));
 AND2_X1 _577_ (.A1(_215_),
    .A2(net148),
    .ZN(_224_));
 MUX2_X1 _578_ (.A(_223_),
    .B(_224_),
    .S(_202_),
    .Z(_053_));
 INV_X1 _579_ (.A(net47),
    .ZN(_225_));
 NOR2_X1 _580_ (.A1(_077_),
    .A2(net1),
    .ZN(_226_));
 AOI221_X1 _581_ (.A(_185_),
    .B1(_088_),
    .B2(_225_),
    .C1(_148_),
    .C2(_226_),
    .ZN(_227_));
 AND2_X1 _582_ (.A1(_215_),
    .A2(net149),
    .ZN(_228_));
 MUX2_X1 _583_ (.A(_227_),
    .B(_228_),
    .S(_202_),
    .Z(_054_));
 NAND2_X1 _584_ (.A1(_089_),
    .A2(net48),
    .ZN(_229_));
 OAI211_X2 _585_ (.A(_079_),
    .B(net2),
    .C1(_162_),
    .C2(_163_),
    .ZN(_230_));
 AOI21_X1 _586_ (.A(_180_),
    .B1(_229_),
    .B2(_230_),
    .ZN(_231_));
 AND2_X1 _587_ (.A1(_215_),
    .A2(net150),
    .ZN(_232_));
 MUX2_X1 _588_ (.A(_231_),
    .B(_232_),
    .S(_202_),
    .Z(_055_));
 NAND2_X1 _589_ (.A1(_089_),
    .A2(net49),
    .ZN(_233_));
 BUF_X8 _590_ (.A(_078_),
    .Z(_234_));
 OAI211_X2 _591_ (.A(_234_),
    .B(net3),
    .C1(_162_),
    .C2(_163_),
    .ZN(_235_));
 AOI21_X1 _592_ (.A(_180_),
    .B1(_233_),
    .B2(_235_),
    .ZN(_236_));
 AND2_X1 _593_ (.A1(_215_),
    .A2(net151),
    .ZN(_237_));
 MUX2_X1 _594_ (.A(_236_),
    .B(_237_),
    .S(_202_),
    .Z(_056_));
 NAND2_X1 _595_ (.A1(_208_),
    .A2(net50),
    .ZN(_238_));
 OAI211_X2 _596_ (.A(_234_),
    .B(net4),
    .C1(_161_),
    .C2(_163_),
    .ZN(_239_));
 AOI21_X1 _597_ (.A(_180_),
    .B1(_238_),
    .B2(_239_),
    .ZN(_240_));
 AND2_X1 _598_ (.A1(_215_),
    .A2(net152),
    .ZN(_241_));
 MUX2_X1 _599_ (.A(_240_),
    .B(_241_),
    .S(_202_),
    .Z(_057_));
 NAND2_X1 _600_ (.A1(_208_),
    .A2(net51),
    .ZN(_242_));
 OAI211_X2 _601_ (.A(_234_),
    .B(net5),
    .C1(_161_),
    .C2(_145_),
    .ZN(_243_));
 AOI21_X1 _602_ (.A(_180_),
    .B1(_242_),
    .B2(_243_),
    .ZN(_244_));
 AND2_X1 _603_ (.A1(_215_),
    .A2(net153),
    .ZN(_245_));
 BUF_X8 _604_ (.A(_154_),
    .Z(_246_));
 MUX2_X1 _605_ (.A(_244_),
    .B(_245_),
    .S(_246_),
    .Z(_058_));
 NAND2_X1 _606_ (.A1(_208_),
    .A2(net52),
    .ZN(_247_));
 OAI211_X2 _607_ (.A(_234_),
    .B(net6),
    .C1(_161_),
    .C2(_145_),
    .ZN(_248_));
 AOI21_X1 _608_ (.A(_180_),
    .B1(_247_),
    .B2(_248_),
    .ZN(_249_));
 AND2_X1 _609_ (.A1(_215_),
    .A2(net154),
    .ZN(_250_));
 MUX2_X1 _610_ (.A(_249_),
    .B(_250_),
    .S(_246_),
    .Z(_059_));
 INV_X1 _611_ (.A(net53),
    .ZN(_251_));
 NOR2_X1 _612_ (.A1(_077_),
    .A2(net22),
    .ZN(_252_));
 AOI221_X1 _613_ (.A(_185_),
    .B1(_149_),
    .B2(_251_),
    .C1(_148_),
    .C2(_252_),
    .ZN(_253_));
 AND2_X1 _614_ (.A1(_215_),
    .A2(net155),
    .ZN(_254_));
 MUX2_X1 _615_ (.A(_253_),
    .B(_254_),
    .S(_246_),
    .Z(_060_));
 NAND2_X1 _616_ (.A1(_208_),
    .A2(net54),
    .ZN(_255_));
 OAI211_X2 _617_ (.A(_234_),
    .B(net7),
    .C1(_161_),
    .C2(_145_),
    .ZN(_256_));
 AOI21_X1 _618_ (.A(_180_),
    .B1(_255_),
    .B2(_256_),
    .ZN(_257_));
 AND2_X1 _619_ (.A1(_139_),
    .A2(net156),
    .ZN(_258_));
 MUX2_X1 _620_ (.A(_257_),
    .B(_258_),
    .S(_246_),
    .Z(_061_));
 NAND2_X1 _621_ (.A1(_208_),
    .A2(net55),
    .ZN(_259_));
 OAI211_X2 _622_ (.A(_234_),
    .B(net8),
    .C1(_161_),
    .C2(_145_),
    .ZN(_260_));
 AOI21_X1 _623_ (.A(_086_),
    .B1(_259_),
    .B2(_260_),
    .ZN(_261_));
 AND2_X1 _624_ (.A1(_139_),
    .A2(net157),
    .ZN(_262_));
 MUX2_X1 _625_ (.A(_261_),
    .B(_262_),
    .S(_246_),
    .Z(_062_));
 NAND2_X1 _626_ (.A1(_208_),
    .A2(net56),
    .ZN(_263_));
 OAI211_X2 _627_ (.A(_234_),
    .B(net23),
    .C1(_161_),
    .C2(_145_),
    .ZN(_264_));
 AOI21_X1 _628_ (.A(_086_),
    .B1(_263_),
    .B2(_264_),
    .ZN(_265_));
 AND2_X1 _629_ (.A1(_139_),
    .A2(net158),
    .ZN(_266_));
 MUX2_X1 _630_ (.A(_265_),
    .B(_266_),
    .S(_246_),
    .Z(_063_));
 NAND2_X1 _631_ (.A1(_208_),
    .A2(net57),
    .ZN(_267_));
 OAI211_X2 _632_ (.A(_234_),
    .B(net24),
    .C1(_161_),
    .C2(_145_),
    .ZN(_268_));
 AOI21_X1 _633_ (.A(_086_),
    .B1(_267_),
    .B2(_268_),
    .ZN(_269_));
 AND2_X1 _634_ (.A1(_139_),
    .A2(net159),
    .ZN(_270_));
 MUX2_X1 _635_ (.A(_269_),
    .B(_270_),
    .S(_246_),
    .Z(_064_));
 INV_X1 _636_ (.A(net58),
    .ZN(_271_));
 NOR2_X1 _637_ (.A1(_077_),
    .A2(net25),
    .ZN(_272_));
 AOI221_X1 _638_ (.A(_185_),
    .B1(_149_),
    .B2(_271_),
    .C1(_147_),
    .C2(_272_),
    .ZN(_273_));
 AND2_X1 _639_ (.A1(_139_),
    .A2(net160),
    .ZN(_274_));
 MUX2_X1 _640_ (.A(_273_),
    .B(_274_),
    .S(_246_),
    .Z(_065_));
 INV_X1 _641_ (.A(net59),
    .ZN(_275_));
 NOR2_X1 _642_ (.A1(_077_),
    .A2(net26),
    .ZN(_276_));
 AOI221_X1 _643_ (.A(_185_),
    .B1(_149_),
    .B2(_275_),
    .C1(_147_),
    .C2(_276_),
    .ZN(_277_));
 AND2_X1 _644_ (.A1(_139_),
    .A2(net161),
    .ZN(_278_));
 MUX2_X1 _645_ (.A(_277_),
    .B(_278_),
    .S(_246_),
    .Z(_066_));
 NAND2_X1 _646_ (.A1(_208_),
    .A2(net60),
    .ZN(_279_));
 OAI211_X2 _647_ (.A(_234_),
    .B(net27),
    .C1(_161_),
    .C2(_145_),
    .ZN(_280_));
 AOI21_X1 _648_ (.A(_086_),
    .B1(_279_),
    .B2(_280_),
    .ZN(_281_));
 AND2_X1 _649_ (.A1(_139_),
    .A2(net162),
    .ZN(_282_));
 MUX2_X1 _650_ (.A(_281_),
    .B(_282_),
    .S(_246_),
    .Z(_067_));
 INV_X1 _651_ (.A(net61),
    .ZN(_283_));
 NOR2_X1 _652_ (.A1(_077_),
    .A2(net28),
    .ZN(_284_));
 AOI221_X1 _653_ (.A(_185_),
    .B1(_149_),
    .B2(_283_),
    .C1(_147_),
    .C2(_284_),
    .ZN(_285_));
 AND2_X1 _654_ (.A1(_139_),
    .A2(net163),
    .ZN(_286_));
 MUX2_X1 _655_ (.A(_285_),
    .B(_286_),
    .S(_154_),
    .Z(_068_));
 NAND2_X1 _656_ (.A1(_208_),
    .A2(net62),
    .ZN(_287_));
 OAI211_X2 _657_ (.A(_234_),
    .B(net29),
    .C1(_161_),
    .C2(_145_),
    .ZN(_288_));
 AOI21_X1 _658_ (.A(_086_),
    .B1(_287_),
    .B2(_288_),
    .ZN(_289_));
 AND2_X1 _659_ (.A1(_139_),
    .A2(net164),
    .ZN(_290_));
 MUX2_X1 _660_ (.A(_289_),
    .B(_290_),
    .S(_154_),
    .Z(_069_));
 INV_X1 _661_ (.A(_081_),
    .ZN(_291_));
 NAND3_X1 _662_ (.A1(_291_),
    .A2(_096_),
    .A3(_004_),
    .ZN(_292_));
 OAI21_X1 _663_ (.A(_077_),
    .B1(is_write_op),
    .B2(_080_),
    .ZN(_293_));
 AND3_X1 _664_ (.A1(_097_),
    .A2(_292_),
    .A3(_293_),
    .ZN(_294_));
 OR2_X1 _665_ (.A1(_076_),
    .A2(_081_),
    .ZN(_295_));
 AOI21_X1 _666_ (.A(_295_),
    .B1(_004_),
    .B2(_096_),
    .ZN(_296_));
 AOI22_X1 _667_ (.A1(_081_),
    .A2(_082_),
    .B1(_097_),
    .B2(_296_),
    .ZN(_297_));
 NAND2_X1 _668_ (.A1(_097_),
    .A2(_296_),
    .ZN(_298_));
 INV_X1 _669_ (.A(net165),
    .ZN(_299_));
 AOI221_X1 _670_ (.A(_087_),
    .B1(_294_),
    .B2(_297_),
    .C1(_298_),
    .C2(_299_),
    .ZN(_070_));
 AOI21_X1 _671_ (.A(_162_),
    .B1(_092_),
    .B2(_091_),
    .ZN(_300_));
 NOR2_X1 _672_ (.A1(_087_),
    .A2(_300_),
    .ZN(_071_));
 NAND2_X1 _673_ (.A1(_091_),
    .A2(net30),
    .ZN(_301_));
 AOI22_X1 _674_ (.A1(_091_),
    .A2(_092_),
    .B1(_301_),
    .B2(is_write_op),
    .ZN(_302_));
 NOR2_X1 _675_ (.A1(_087_),
    .A2(_302_),
    .ZN(_072_));
 OR2_X1 _676_ (.A1(_081_),
    .A2(\state[3] ),
    .ZN(net166));
 DFF_X1 \first_write_done$_SDFFE_PN0P_  (.D(_071_),
    .CK(clknet_3_1__leaf_clk),
    .Q(first_write_done),
    .QN(_370_));
 DFF_X2 \is_write_op$_SDFFE_PN0P_  (.D(_072_),
    .CK(clknet_3_0__leaf_clk),
    .Q(is_write_op),
    .QN(_369_));
 DFF_X1 \mem_rdata[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net100),
    .QN(_368_));
 DFF_X1 \mem_rdata[10]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net101),
    .QN(_367_));
 DFF_X1 \mem_rdata[11]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net102),
    .QN(_366_));
 DFF_X1 \mem_rdata[12]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net103),
    .QN(_365_));
 DFF_X1 \mem_rdata[13]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net104),
    .QN(_364_));
 DFF_X1 \mem_rdata[14]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net105),
    .QN(_363_));
 DFF_X1 \mem_rdata[15]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net106),
    .QN(_362_));
 DFF_X1 \mem_rdata[16]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net107),
    .QN(_361_));
 DFF_X1 \mem_rdata[17]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net108),
    .QN(_360_));
 DFF_X1 \mem_rdata[18]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net109),
    .QN(_359_));
 DFF_X1 \mem_rdata[19]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net110),
    .QN(_358_));
 DFF_X1 \mem_rdata[1]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net111),
    .QN(_357_));
 DFF_X1 \mem_rdata[20]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net112),
    .QN(_356_));
 DFF_X1 \mem_rdata[21]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net113),
    .QN(_355_));
 DFF_X1 \mem_rdata[22]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net114),
    .QN(_354_));
 DFF_X1 \mem_rdata[23]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net115),
    .QN(_353_));
 DFF_X1 \mem_rdata[24]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net116),
    .QN(_352_));
 DFF_X1 \mem_rdata[25]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net117),
    .QN(_351_));
 DFF_X1 \mem_rdata[26]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net118),
    .QN(_350_));
 DFF_X1 \mem_rdata[27]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net119),
    .QN(_349_));
 DFF_X1 \mem_rdata[28]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net120),
    .QN(_348_));
 DFF_X1 \mem_rdata[29]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net121),
    .QN(_347_));
 DFF_X1 \mem_rdata[2]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net122),
    .QN(_346_));
 DFF_X1 \mem_rdata[30]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net123),
    .QN(_345_));
 DFF_X1 \mem_rdata[31]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net124),
    .QN(_344_));
 DFF_X1 \mem_rdata[3]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net125),
    .QN(_343_));
 DFF_X1 \mem_rdata[4]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net126),
    .QN(_342_));
 DFF_X1 \mem_rdata[5]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net127),
    .QN(_341_));
 DFF_X1 \mem_rdata[6]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net128),
    .QN(_340_));
 DFF_X1 \mem_rdata[7]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net129),
    .QN(_339_));
 DFF_X1 \mem_rdata[8]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net130),
    .QN(_338_));
 DFF_X1 \mem_rdata[9]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net131),
    .QN(_337_));
 DFF_X1 \mem_ready$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_3_2__leaf_clk),
    .Q(net132),
    .QN(_371_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\state[0] ),
    .QN(_372_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_002_),
    .CK(clknet_3_2__leaf_clk),
    .Q(\state[1] ),
    .QN(_373_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_003_),
    .CK(clknet_3_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_004_));
 DFF_X1 \state[3]$_DFF_P_  (.D(_000_),
    .CK(clknet_3_0__leaf_clk),
    .Q(\state[3] ),
    .QN(_336_));
 DFF_X1 \tx_data[0]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net133),
    .QN(_335_));
 DFF_X1 \tx_data[10]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_3_3__leaf_clk),
    .Q(net134),
    .QN(_334_));
 DFF_X1 \tx_data[11]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_3_6__leaf_clk),
    .Q(net135),
    .QN(_333_));
 DFF_X1 \tx_data[12]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net136),
    .QN(_332_));
 DFF_X1 \tx_data[13]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net137),
    .QN(_331_));
 DFF_X1 \tx_data[14]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net138),
    .QN(_330_));
 DFF_X1 \tx_data[15]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net139),
    .QN(_329_));
 DFF_X1 \tx_data[16]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net140),
    .QN(_328_));
 DFF_X1 \tx_data[17]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net141),
    .QN(_327_));
 DFF_X1 \tx_data[18]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_3_7__leaf_clk),
    .Q(net142),
    .QN(_326_));
 DFF_X1 \tx_data[19]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net143),
    .QN(_325_));
 DFF_X1 \tx_data[1]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net144),
    .QN(_324_));
 DFF_X1 \tx_data[20]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net145),
    .QN(_323_));
 DFF_X1 \tx_data[21]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net146),
    .QN(_322_));
 DFF_X1 \tx_data[22]$_SDFFE_PN0P_  (.D(_052_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net147),
    .QN(_321_));
 DFF_X1 \tx_data[23]$_SDFFE_PN0P_  (.D(_053_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net148),
    .QN(_320_));
 DFF_X1 \tx_data[24]$_SDFFE_PN0P_  (.D(_054_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net149),
    .QN(_319_));
 DFF_X1 \tx_data[25]$_SDFFE_PN0P_  (.D(_055_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net150),
    .QN(_318_));
 DFF_X1 \tx_data[26]$_SDFFE_PN0P_  (.D(_056_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net151),
    .QN(_317_));
 DFF_X1 \tx_data[27]$_SDFFE_PN0P_  (.D(_057_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net152),
    .QN(_316_));
 DFF_X1 \tx_data[28]$_SDFFE_PN0P_  (.D(_058_),
    .CK(clknet_3_5__leaf_clk),
    .Q(net153),
    .QN(_315_));
 DFF_X1 \tx_data[29]$_SDFFE_PN0P_  (.D(_059_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net154),
    .QN(_314_));
 DFF_X1 \tx_data[2]$_SDFFE_PN0P_  (.D(_060_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net155),
    .QN(_313_));
 DFF_X1 \tx_data[30]$_SDFFE_PN0P_  (.D(_061_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net156),
    .QN(_312_));
 DFF_X1 \tx_data[31]$_SDFFE_PN0P_  (.D(_062_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net157),
    .QN(_311_));
 DFF_X1 \tx_data[3]$_SDFFE_PN0P_  (.D(_063_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net158),
    .QN(_310_));
 DFF_X1 \tx_data[4]$_SDFFE_PN0P_  (.D(_064_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net159),
    .QN(_309_));
 DFF_X1 \tx_data[5]$_SDFFE_PN0P_  (.D(_065_),
    .CK(clknet_3_4__leaf_clk),
    .Q(net160),
    .QN(_308_));
 DFF_X1 \tx_data[6]$_SDFFE_PN0P_  (.D(_066_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net161),
    .QN(_307_));
 DFF_X1 \tx_data[7]$_SDFFE_PN0P_  (.D(_067_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net162),
    .QN(_306_));
 DFF_X1 \tx_data[8]$_SDFFE_PN0P_  (.D(_068_),
    .CK(clknet_3_1__leaf_clk),
    .Q(net163),
    .QN(_305_));
 DFF_X1 \tx_data[9]$_SDFFE_PN0P_  (.D(_069_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net164),
    .QN(_304_));
 DFF_X2 \tx_valid$_SDFFE_PN0P_  (.D(_070_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net165),
    .QN(_303_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_53 ();
 BUF_X1 input1 (.A(dest_id[0]),
    .Z(net1));
 BUF_X1 input2 (.A(dest_id[1]),
    .Z(net2));
 BUF_X1 input3 (.A(dest_id[2]),
    .Z(net3));
 BUF_X1 input4 (.A(dest_id[3]),
    .Z(net4));
 BUF_X1 input5 (.A(dest_id[4]),
    .Z(net5));
 BUF_X1 input6 (.A(dest_id[5]),
    .Z(net6));
 BUF_X1 input7 (.A(dest_id[6]),
    .Z(net7));
 BUF_X1 input8 (.A(dest_id[7]),
    .Z(net8));
 BUF_X1 input9 (.A(mem_addr[0]),
    .Z(net9));
 BUF_X1 input10 (.A(mem_addr[10]),
    .Z(net10));
 BUF_X1 input11 (.A(mem_addr[11]),
    .Z(net11));
 BUF_X1 input12 (.A(mem_addr[12]),
    .Z(net12));
 BUF_X1 input13 (.A(mem_addr[13]),
    .Z(net13));
 BUF_X1 input14 (.A(mem_addr[14]),
    .Z(net14));
 BUF_X1 input15 (.A(mem_addr[15]),
    .Z(net15));
 BUF_X1 input16 (.A(mem_addr[16]),
    .Z(net16));
 BUF_X1 input17 (.A(mem_addr[17]),
    .Z(net17));
 BUF_X1 input18 (.A(mem_addr[18]),
    .Z(net18));
 BUF_X1 input19 (.A(mem_addr[19]),
    .Z(net19));
 BUF_X1 input20 (.A(mem_addr[1]),
    .Z(net20));
 BUF_X1 input21 (.A(mem_addr[20]),
    .Z(net21));
 BUF_X1 input22 (.A(mem_addr[2]),
    .Z(net22));
 BUF_X1 input23 (.A(mem_addr[3]),
    .Z(net23));
 BUF_X1 input24 (.A(mem_addr[4]),
    .Z(net24));
 BUF_X1 input25 (.A(mem_addr[5]),
    .Z(net25));
 BUF_X1 input26 (.A(mem_addr[6]),
    .Z(net26));
 BUF_X1 input27 (.A(mem_addr[7]),
    .Z(net27));
 BUF_X1 input28 (.A(mem_addr[8]),
    .Z(net28));
 BUF_X1 input29 (.A(mem_addr[9]),
    .Z(net29));
 BUF_X1 input30 (.A(mem_read),
    .Z(net30));
 BUF_X1 input31 (.A(mem_wdata[0]),
    .Z(net31));
 BUF_X1 input32 (.A(mem_wdata[10]),
    .Z(net32));
 BUF_X1 input33 (.A(mem_wdata[11]),
    .Z(net33));
 BUF_X1 input34 (.A(mem_wdata[12]),
    .Z(net34));
 BUF_X1 input35 (.A(mem_wdata[13]),
    .Z(net35));
 BUF_X1 input36 (.A(mem_wdata[14]),
    .Z(net36));
 BUF_X1 input37 (.A(mem_wdata[15]),
    .Z(net37));
 BUF_X1 input38 (.A(mem_wdata[16]),
    .Z(net38));
 BUF_X1 input39 (.A(mem_wdata[17]),
    .Z(net39));
 BUF_X1 input40 (.A(mem_wdata[18]),
    .Z(net40));
 BUF_X1 input41 (.A(mem_wdata[19]),
    .Z(net41));
 BUF_X1 input42 (.A(mem_wdata[1]),
    .Z(net42));
 BUF_X1 input43 (.A(mem_wdata[20]),
    .Z(net43));
 BUF_X1 input44 (.A(mem_wdata[21]),
    .Z(net44));
 BUF_X1 input45 (.A(mem_wdata[22]),
    .Z(net45));
 BUF_X1 input46 (.A(mem_wdata[23]),
    .Z(net46));
 BUF_X1 input47 (.A(mem_wdata[24]),
    .Z(net47));
 BUF_X1 input48 (.A(mem_wdata[25]),
    .Z(net48));
 BUF_X1 input49 (.A(mem_wdata[26]),
    .Z(net49));
 BUF_X1 input50 (.A(mem_wdata[27]),
    .Z(net50));
 BUF_X1 input51 (.A(mem_wdata[28]),
    .Z(net51));
 BUF_X1 input52 (.A(mem_wdata[29]),
    .Z(net52));
 BUF_X1 input53 (.A(mem_wdata[2]),
    .Z(net53));
 BUF_X1 input54 (.A(mem_wdata[30]),
    .Z(net54));
 BUF_X1 input55 (.A(mem_wdata[31]),
    .Z(net55));
 BUF_X1 input56 (.A(mem_wdata[3]),
    .Z(net56));
 BUF_X1 input57 (.A(mem_wdata[4]),
    .Z(net57));
 BUF_X1 input58 (.A(mem_wdata[5]),
    .Z(net58));
 BUF_X1 input59 (.A(mem_wdata[6]),
    .Z(net59));
 BUF_X1 input60 (.A(mem_wdata[7]),
    .Z(net60));
 BUF_X1 input61 (.A(mem_wdata[8]),
    .Z(net61));
 BUF_X1 input62 (.A(mem_wdata[9]),
    .Z(net62));
 BUF_X1 input63 (.A(msg_type[0]),
    .Z(net63));
 BUF_X1 input64 (.A(msg_type[1]),
    .Z(net64));
 BUF_X1 input65 (.A(msg_type[2]),
    .Z(net65));
 BUF_X1 input66 (.A(router_in_ready),
    .Z(net66));
 BUF_X1 input67 (.A(router_out_data[0]),
    .Z(net67));
 BUF_X1 input68 (.A(router_out_data[10]),
    .Z(net68));
 BUF_X1 input69 (.A(router_out_data[11]),
    .Z(net69));
 BUF_X1 input70 (.A(router_out_data[12]),
    .Z(net70));
 BUF_X1 input71 (.A(router_out_data[13]),
    .Z(net71));
 BUF_X1 input72 (.A(router_out_data[14]),
    .Z(net72));
 BUF_X1 input73 (.A(router_out_data[15]),
    .Z(net73));
 BUF_X1 input74 (.A(router_out_data[16]),
    .Z(net74));
 BUF_X1 input75 (.A(router_out_data[17]),
    .Z(net75));
 BUF_X1 input76 (.A(router_out_data[18]),
    .Z(net76));
 BUF_X1 input77 (.A(router_out_data[19]),
    .Z(net77));
 BUF_X1 input78 (.A(router_out_data[1]),
    .Z(net78));
 BUF_X1 input79 (.A(router_out_data[20]),
    .Z(net79));
 BUF_X1 input80 (.A(router_out_data[21]),
    .Z(net80));
 BUF_X1 input81 (.A(router_out_data[22]),
    .Z(net81));
 BUF_X1 input82 (.A(router_out_data[23]),
    .Z(net82));
 BUF_X1 input83 (.A(router_out_data[24]),
    .Z(net83));
 BUF_X1 input84 (.A(router_out_data[25]),
    .Z(net84));
 BUF_X1 input85 (.A(router_out_data[26]),
    .Z(net85));
 BUF_X1 input86 (.A(router_out_data[27]),
    .Z(net86));
 BUF_X1 input87 (.A(router_out_data[28]),
    .Z(net87));
 BUF_X1 input88 (.A(router_out_data[29]),
    .Z(net88));
 BUF_X1 input89 (.A(router_out_data[2]),
    .Z(net89));
 BUF_X1 input90 (.A(router_out_data[30]),
    .Z(net90));
 BUF_X1 input91 (.A(router_out_data[31]),
    .Z(net91));
 BUF_X1 input92 (.A(router_out_data[3]),
    .Z(net92));
 BUF_X1 input93 (.A(router_out_data[4]),
    .Z(net93));
 BUF_X1 input94 (.A(router_out_data[5]),
    .Z(net94));
 BUF_X1 input95 (.A(router_out_data[6]),
    .Z(net95));
 BUF_X1 input96 (.A(router_out_data[7]),
    .Z(net96));
 BUF_X1 input97 (.A(router_out_data[8]),
    .Z(net97));
 BUF_X1 input98 (.A(router_out_data[9]),
    .Z(net98));
 CLKBUF_X2 input99 (.A(router_out_valid),
    .Z(net99));
 BUF_X1 output100 (.A(net100),
    .Z(mem_rdata[0]));
 BUF_X1 output101 (.A(net101),
    .Z(mem_rdata[10]));
 BUF_X1 output102 (.A(net102),
    .Z(mem_rdata[11]));
 BUF_X1 output103 (.A(net103),
    .Z(mem_rdata[12]));
 BUF_X1 output104 (.A(net104),
    .Z(mem_rdata[13]));
 BUF_X1 output105 (.A(net105),
    .Z(mem_rdata[14]));
 BUF_X1 output106 (.A(net106),
    .Z(mem_rdata[15]));
 BUF_X1 output107 (.A(net107),
    .Z(mem_rdata[16]));
 BUF_X1 output108 (.A(net108),
    .Z(mem_rdata[17]));
 BUF_X1 output109 (.A(net109),
    .Z(mem_rdata[18]));
 BUF_X1 output110 (.A(net110),
    .Z(mem_rdata[19]));
 BUF_X1 output111 (.A(net111),
    .Z(mem_rdata[1]));
 BUF_X1 output112 (.A(net112),
    .Z(mem_rdata[20]));
 BUF_X1 output113 (.A(net113),
    .Z(mem_rdata[21]));
 BUF_X1 output114 (.A(net114),
    .Z(mem_rdata[22]));
 BUF_X1 output115 (.A(net115),
    .Z(mem_rdata[23]));
 BUF_X1 output116 (.A(net116),
    .Z(mem_rdata[24]));
 BUF_X1 output117 (.A(net117),
    .Z(mem_rdata[25]));
 BUF_X1 output118 (.A(net118),
    .Z(mem_rdata[26]));
 BUF_X1 output119 (.A(net119),
    .Z(mem_rdata[27]));
 BUF_X1 output120 (.A(net120),
    .Z(mem_rdata[28]));
 BUF_X1 output121 (.A(net121),
    .Z(mem_rdata[29]));
 BUF_X1 output122 (.A(net122),
    .Z(mem_rdata[2]));
 BUF_X1 output123 (.A(net123),
    .Z(mem_rdata[30]));
 BUF_X1 output124 (.A(net124),
    .Z(mem_rdata[31]));
 BUF_X1 output125 (.A(net125),
    .Z(mem_rdata[3]));
 BUF_X1 output126 (.A(net126),
    .Z(mem_rdata[4]));
 BUF_X1 output127 (.A(net127),
    .Z(mem_rdata[5]));
 BUF_X1 output128 (.A(net128),
    .Z(mem_rdata[6]));
 BUF_X1 output129 (.A(net129),
    .Z(mem_rdata[7]));
 BUF_X1 output130 (.A(net130),
    .Z(mem_rdata[8]));
 BUF_X1 output131 (.A(net131),
    .Z(mem_rdata[9]));
 BUF_X1 output132 (.A(net132),
    .Z(mem_ready));
 BUF_X1 output133 (.A(net133),
    .Z(router_in_data[0]));
 BUF_X1 output134 (.A(net134),
    .Z(router_in_data[10]));
 BUF_X1 output135 (.A(net135),
    .Z(router_in_data[11]));
 BUF_X1 output136 (.A(net136),
    .Z(router_in_data[12]));
 BUF_X1 output137 (.A(net137),
    .Z(router_in_data[13]));
 BUF_X1 output138 (.A(net138),
    .Z(router_in_data[14]));
 BUF_X1 output139 (.A(net139),
    .Z(router_in_data[15]));
 BUF_X1 output140 (.A(net140),
    .Z(router_in_data[16]));
 BUF_X1 output141 (.A(net141),
    .Z(router_in_data[17]));
 BUF_X1 output142 (.A(net142),
    .Z(router_in_data[18]));
 BUF_X1 output143 (.A(net143),
    .Z(router_in_data[19]));
 BUF_X1 output144 (.A(net144),
    .Z(router_in_data[1]));
 BUF_X1 output145 (.A(net145),
    .Z(router_in_data[20]));
 BUF_X1 output146 (.A(net146),
    .Z(router_in_data[21]));
 BUF_X1 output147 (.A(net147),
    .Z(router_in_data[22]));
 BUF_X1 output148 (.A(net148),
    .Z(router_in_data[23]));
 BUF_X1 output149 (.A(net149),
    .Z(router_in_data[24]));
 BUF_X1 output150 (.A(net150),
    .Z(router_in_data[25]));
 BUF_X1 output151 (.A(net151),
    .Z(router_in_data[26]));
 BUF_X1 output152 (.A(net152),
    .Z(router_in_data[27]));
 BUF_X1 output153 (.A(net153),
    .Z(router_in_data[28]));
 BUF_X1 output154 (.A(net154),
    .Z(router_in_data[29]));
 BUF_X1 output155 (.A(net155),
    .Z(router_in_data[2]));
 BUF_X1 output156 (.A(net156),
    .Z(router_in_data[30]));
 BUF_X1 output157 (.A(net157),
    .Z(router_in_data[31]));
 BUF_X1 output158 (.A(net158),
    .Z(router_in_data[3]));
 BUF_X1 output159 (.A(net159),
    .Z(router_in_data[4]));
 BUF_X1 output160 (.A(net160),
    .Z(router_in_data[5]));
 BUF_X1 output161 (.A(net161),
    .Z(router_in_data[6]));
 BUF_X1 output162 (.A(net162),
    .Z(router_in_data[7]));
 BUF_X1 output163 (.A(net163),
    .Z(router_in_data[8]));
 BUF_X1 output164 (.A(net164),
    .Z(router_in_data[9]));
 BUF_X1 output165 (.A(net165),
    .Z(router_in_valid));
 BUF_X1 output166 (.A(net166),
    .Z(router_out_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X2 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X4 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X2 clkload2 (.A(clknet_3_3__leaf_clk));
 INV_X2 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_5__leaf_clk));
 INV_X2 clkload5 (.A(clknet_3_6__leaf_clk));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_24 ();
 FILLCELL_X2 FILLER_0_60 ();
 FILLCELL_X1 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_108 ();
 FILLCELL_X1 FILLER_0_112 ();
 FILLCELL_X1 FILLER_0_116 ();
 FILLCELL_X1 FILLER_0_128 ();
 FILLCELL_X2 FILLER_0_148 ();
 FILLCELL_X8 FILLER_0_167 ();
 FILLCELL_X16 FILLER_0_182 ();
 FILLCELL_X4 FILLER_0_198 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X4 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_21 ();
 FILLCELL_X2 FILLER_1_67 ();
 FILLCELL_X2 FILLER_1_82 ();
 FILLCELL_X2 FILLER_1_90 ();
 FILLCELL_X2 FILLER_1_147 ();
 FILLCELL_X2 FILLER_1_197 ();
 FILLCELL_X16 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_17 ();
 FILLCELL_X2 FILLER_2_25 ();
 FILLCELL_X16 FILLER_2_81 ();
 FILLCELL_X2 FILLER_2_97 ();
 FILLCELL_X1 FILLER_2_99 ();
 FILLCELL_X1 FILLER_2_119 ();
 FILLCELL_X1 FILLER_2_123 ();
 FILLCELL_X8 FILLER_2_130 ();
 FILLCELL_X1 FILLER_2_138 ();
 FILLCELL_X4 FILLER_2_143 ();
 FILLCELL_X2 FILLER_2_150 ();
 FILLCELL_X1 FILLER_2_152 ();
 FILLCELL_X2 FILLER_2_170 ();
 FILLCELL_X1 FILLER_2_172 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X1 FILLER_2_201 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X2 FILLER_3_60 ();
 FILLCELL_X2 FILLER_3_79 ();
 FILLCELL_X2 FILLER_3_89 ();
 FILLCELL_X2 FILLER_3_117 ();
 FILLCELL_X1 FILLER_3_119 ();
 FILLCELL_X4 FILLER_3_138 ();
 FILLCELL_X2 FILLER_3_142 ();
 FILLCELL_X1 FILLER_3_144 ();
 FILLCELL_X2 FILLER_3_149 ();
 FILLCELL_X4 FILLER_3_162 ();
 FILLCELL_X2 FILLER_3_166 ();
 FILLCELL_X1 FILLER_3_168 ();
 FILLCELL_X1 FILLER_3_198 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X1 FILLER_4_29 ();
 FILLCELL_X1 FILLER_4_47 ();
 FILLCELL_X2 FILLER_4_51 ();
 FILLCELL_X2 FILLER_4_58 ();
 FILLCELL_X2 FILLER_4_73 ();
 FILLCELL_X16 FILLER_4_100 ();
 FILLCELL_X8 FILLER_4_116 ();
 FILLCELL_X1 FILLER_4_124 ();
 FILLCELL_X8 FILLER_4_151 ();
 FILLCELL_X2 FILLER_4_159 ();
 FILLCELL_X1 FILLER_4_181 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_39 ();
 FILLCELL_X4 FILLER_5_54 ();
 FILLCELL_X1 FILLER_5_94 ();
 FILLCELL_X4 FILLER_5_101 ();
 FILLCELL_X16 FILLER_5_109 ();
 FILLCELL_X4 FILLER_5_125 ();
 FILLCELL_X2 FILLER_5_131 ();
 FILLCELL_X32 FILLER_5_136 ();
 FILLCELL_X2 FILLER_5_168 ();
 FILLCELL_X1 FILLER_5_170 ();
 FILLCELL_X4 FILLER_5_174 ();
 FILLCELL_X2 FILLER_5_178 ();
 FILLCELL_X1 FILLER_5_180 ();
 FILLCELL_X2 FILLER_5_191 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_17 ();
 FILLCELL_X4 FILLER_6_25 ();
 FILLCELL_X2 FILLER_6_29 ();
 FILLCELL_X32 FILLER_6_48 ();
 FILLCELL_X4 FILLER_6_80 ();
 FILLCELL_X2 FILLER_6_84 ();
 FILLCELL_X8 FILLER_6_92 ();
 FILLCELL_X1 FILLER_6_100 ();
 FILLCELL_X2 FILLER_6_125 ();
 FILLCELL_X1 FILLER_6_127 ();
 FILLCELL_X4 FILLER_6_141 ();
 FILLCELL_X2 FILLER_6_145 ();
 FILLCELL_X4 FILLER_6_151 ();
 FILLCELL_X1 FILLER_6_155 ();
 FILLCELL_X1 FILLER_6_163 ();
 FILLCELL_X2 FILLER_6_170 ();
 FILLCELL_X1 FILLER_6_172 ();
 FILLCELL_X2 FILLER_6_191 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_17 ();
 FILLCELL_X32 FILLER_7_26 ();
 FILLCELL_X2 FILLER_7_58 ();
 FILLCELL_X4 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_72 ();
 FILLCELL_X2 FILLER_7_94 ();
 FILLCELL_X1 FILLER_7_96 ();
 FILLCELL_X8 FILLER_7_104 ();
 FILLCELL_X2 FILLER_7_112 ();
 FILLCELL_X1 FILLER_7_114 ();
 FILLCELL_X8 FILLER_7_122 ();
 FILLCELL_X1 FILLER_7_152 ();
 FILLCELL_X1 FILLER_7_174 ();
 FILLCELL_X2 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_3 ();
 FILLCELL_X8 FILLER_8_29 ();
 FILLCELL_X4 FILLER_8_37 ();
 FILLCELL_X16 FILLER_8_46 ();
 FILLCELL_X1 FILLER_8_62 ();
 FILLCELL_X32 FILLER_8_92 ();
 FILLCELL_X1 FILLER_8_124 ();
 FILLCELL_X4 FILLER_8_130 ();
 FILLCELL_X2 FILLER_8_134 ();
 FILLCELL_X1 FILLER_8_136 ();
 FILLCELL_X16 FILLER_8_140 ();
 FILLCELL_X4 FILLER_8_156 ();
 FILLCELL_X1 FILLER_8_160 ();
 FILLCELL_X4 FILLER_8_171 ();
 FILLCELL_X1 FILLER_8_175 ();
 FILLCELL_X2 FILLER_8_179 ();
 FILLCELL_X1 FILLER_8_181 ();
 FILLCELL_X2 FILLER_8_184 ();
 FILLCELL_X1 FILLER_8_186 ();
 FILLCELL_X2 FILLER_8_193 ();
 FILLCELL_X1 FILLER_8_195 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_5 ();
 FILLCELL_X8 FILLER_9_10 ();
 FILLCELL_X1 FILLER_9_39 ();
 FILLCELL_X8 FILLER_9_67 ();
 FILLCELL_X2 FILLER_9_75 ();
 FILLCELL_X4 FILLER_9_82 ();
 FILLCELL_X2 FILLER_9_86 ();
 FILLCELL_X8 FILLER_9_95 ();
 FILLCELL_X4 FILLER_9_103 ();
 FILLCELL_X2 FILLER_9_107 ();
 FILLCELL_X8 FILLER_9_122 ();
 FILLCELL_X2 FILLER_9_130 ();
 FILLCELL_X8 FILLER_9_140 ();
 FILLCELL_X4 FILLER_9_148 ();
 FILLCELL_X2 FILLER_9_152 ();
 FILLCELL_X1 FILLER_9_154 ();
 FILLCELL_X4 FILLER_9_158 ();
 FILLCELL_X1 FILLER_9_166 ();
 FILLCELL_X2 FILLER_9_169 ();
 FILLCELL_X4 FILLER_9_180 ();
 FILLCELL_X2 FILLER_9_184 ();
 FILLCELL_X1 FILLER_9_186 ();
 FILLCELL_X1 FILLER_10_49 ();
 FILLCELL_X8 FILLER_10_81 ();
 FILLCELL_X2 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_91 ();
 FILLCELL_X4 FILLER_10_99 ();
 FILLCELL_X8 FILLER_10_108 ();
 FILLCELL_X2 FILLER_10_116 ();
 FILLCELL_X4 FILLER_10_146 ();
 FILLCELL_X1 FILLER_10_150 ();
 FILLCELL_X2 FILLER_10_164 ();
 FILLCELL_X1 FILLER_10_177 ();
 FILLCELL_X4 FILLER_10_181 ();
 FILLCELL_X2 FILLER_10_185 ();
 FILLCELL_X1 FILLER_10_187 ();
 FILLCELL_X1 FILLER_10_198 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X4 FILLER_11_10 ();
 FILLCELL_X1 FILLER_11_14 ();
 FILLCELL_X2 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_51 ();
 FILLCELL_X4 FILLER_11_83 ();
 FILLCELL_X2 FILLER_11_99 ();
 FILLCELL_X32 FILLER_11_114 ();
 FILLCELL_X4 FILLER_11_146 ();
 FILLCELL_X2 FILLER_11_184 ();
 FILLCELL_X1 FILLER_11_198 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X2 FILLER_12_13 ();
 FILLCELL_X1 FILLER_12_15 ();
 FILLCELL_X8 FILLER_12_19 ();
 FILLCELL_X2 FILLER_12_30 ();
 FILLCELL_X1 FILLER_12_32 ();
 FILLCELL_X2 FILLER_12_36 ();
 FILLCELL_X1 FILLER_12_51 ();
 FILLCELL_X2 FILLER_12_76 ();
 FILLCELL_X8 FILLER_12_99 ();
 FILLCELL_X1 FILLER_12_107 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X2 FILLER_12_135 ();
 FILLCELL_X1 FILLER_12_137 ();
 FILLCELL_X2 FILLER_12_166 ();
 FILLCELL_X1 FILLER_12_168 ();
 FILLCELL_X1 FILLER_12_198 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_17 ();
 FILLCELL_X8 FILLER_13_38 ();
 FILLCELL_X2 FILLER_13_46 ();
 FILLCELL_X16 FILLER_13_53 ();
 FILLCELL_X8 FILLER_13_69 ();
 FILLCELL_X2 FILLER_13_77 ();
 FILLCELL_X1 FILLER_13_79 ();
 FILLCELL_X32 FILLER_13_84 ();
 FILLCELL_X16 FILLER_13_116 ();
 FILLCELL_X4 FILLER_13_132 ();
 FILLCELL_X2 FILLER_13_136 ();
 FILLCELL_X1 FILLER_13_138 ();
 FILLCELL_X8 FILLER_13_144 ();
 FILLCELL_X4 FILLER_13_152 ();
 FILLCELL_X1 FILLER_13_156 ();
 FILLCELL_X2 FILLER_13_185 ();
 FILLCELL_X2 FILLER_13_196 ();
 FILLCELL_X1 FILLER_13_198 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_6 ();
 FILLCELL_X1 FILLER_14_24 ();
 FILLCELL_X1 FILLER_14_29 ();
 FILLCELL_X4 FILLER_14_37 ();
 FILLCELL_X2 FILLER_14_41 ();
 FILLCELL_X1 FILLER_14_43 ();
 FILLCELL_X32 FILLER_14_57 ();
 FILLCELL_X8 FILLER_14_89 ();
 FILLCELL_X4 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_106 ();
 FILLCELL_X2 FILLER_14_110 ();
 FILLCELL_X1 FILLER_14_112 ();
 FILLCELL_X8 FILLER_14_117 ();
 FILLCELL_X4 FILLER_14_125 ();
 FILLCELL_X1 FILLER_14_129 ();
 FILLCELL_X16 FILLER_14_137 ();
 FILLCELL_X4 FILLER_14_153 ();
 FILLCELL_X2 FILLER_14_157 ();
 FILLCELL_X1 FILLER_14_166 ();
 FILLCELL_X1 FILLER_14_174 ();
 FILLCELL_X1 FILLER_14_179 ();
 FILLCELL_X2 FILLER_14_191 ();
 FILLCELL_X2 FILLER_15_7 ();
 FILLCELL_X1 FILLER_15_16 ();
 FILLCELL_X2 FILLER_15_37 ();
 FILLCELL_X1 FILLER_15_39 ();
 FILLCELL_X32 FILLER_15_64 ();
 FILLCELL_X32 FILLER_15_96 ();
 FILLCELL_X1 FILLER_15_189 ();
 FILLCELL_X8 FILLER_16_22 ();
 FILLCELL_X4 FILLER_16_30 ();
 FILLCELL_X2 FILLER_16_34 ();
 FILLCELL_X1 FILLER_16_36 ();
 FILLCELL_X32 FILLER_16_45 ();
 FILLCELL_X32 FILLER_16_77 ();
 FILLCELL_X16 FILLER_16_109 ();
 FILLCELL_X8 FILLER_16_125 ();
 FILLCELL_X1 FILLER_16_133 ();
 FILLCELL_X4 FILLER_16_138 ();
 FILLCELL_X1 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_166 ();
 FILLCELL_X1 FILLER_16_170 ();
 FILLCELL_X2 FILLER_16_180 ();
 FILLCELL_X1 FILLER_16_182 ();
 FILLCELL_X1 FILLER_16_185 ();
 FILLCELL_X1 FILLER_16_195 ();
 FILLCELL_X2 FILLER_16_199 ();
 FILLCELL_X1 FILLER_16_201 ();
 FILLCELL_X1 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_104 ();
 FILLCELL_X4 FILLER_17_136 ();
 FILLCELL_X2 FILLER_17_140 ();
 FILLCELL_X1 FILLER_17_142 ();
 FILLCELL_X2 FILLER_17_161 ();
 FILLCELL_X1 FILLER_17_163 ();
 FILLCELL_X8 FILLER_17_188 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X4 FILLER_18_17 ();
 FILLCELL_X2 FILLER_18_21 ();
 FILLCELL_X1 FILLER_18_23 ();
 FILLCELL_X32 FILLER_18_41 ();
 FILLCELL_X16 FILLER_18_73 ();
 FILLCELL_X2 FILLER_18_89 ();
 FILLCELL_X1 FILLER_18_91 ();
 FILLCELL_X2 FILLER_18_116 ();
 FILLCELL_X1 FILLER_18_118 ();
 FILLCELL_X16 FILLER_18_123 ();
 FILLCELL_X8 FILLER_18_139 ();
 FILLCELL_X4 FILLER_18_147 ();
 FILLCELL_X2 FILLER_18_172 ();
 FILLCELL_X1 FILLER_18_181 ();
 FILLCELL_X1 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_23 ();
 FILLCELL_X2 FILLER_19_28 ();
 FILLCELL_X1 FILLER_19_30 ();
 FILLCELL_X32 FILLER_19_51 ();
 FILLCELL_X4 FILLER_19_83 ();
 FILLCELL_X2 FILLER_19_87 ();
 FILLCELL_X1 FILLER_19_89 ();
 FILLCELL_X1 FILLER_19_93 ();
 FILLCELL_X2 FILLER_19_104 ();
 FILLCELL_X1 FILLER_19_106 ();
 FILLCELL_X8 FILLER_19_133 ();
 FILLCELL_X1 FILLER_19_147 ();
 FILLCELL_X8 FILLER_19_151 ();
 FILLCELL_X2 FILLER_19_159 ();
 FILLCELL_X8 FILLER_19_163 ();
 FILLCELL_X4 FILLER_19_171 ();
 FILLCELL_X2 FILLER_19_175 ();
 FILLCELL_X2 FILLER_19_183 ();
 FILLCELL_X1 FILLER_19_185 ();
 FILLCELL_X1 FILLER_19_194 ();
 FILLCELL_X4 FILLER_20_21 ();
 FILLCELL_X2 FILLER_20_25 ();
 FILLCELL_X2 FILLER_20_57 ();
 FILLCELL_X1 FILLER_20_59 ();
 FILLCELL_X2 FILLER_20_67 ();
 FILLCELL_X16 FILLER_20_73 ();
 FILLCELL_X2 FILLER_20_89 ();
 FILLCELL_X8 FILLER_20_93 ();
 FILLCELL_X4 FILLER_20_101 ();
 FILLCELL_X2 FILLER_20_105 ();
 FILLCELL_X1 FILLER_20_107 ();
 FILLCELL_X16 FILLER_20_110 ();
 FILLCELL_X8 FILLER_20_126 ();
 FILLCELL_X2 FILLER_20_138 ();
 FILLCELL_X16 FILLER_20_142 ();
 FILLCELL_X8 FILLER_20_158 ();
 FILLCELL_X1 FILLER_20_166 ();
 FILLCELL_X4 FILLER_20_172 ();
 FILLCELL_X2 FILLER_20_176 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_3 ();
 FILLCELL_X4 FILLER_21_14 ();
 FILLCELL_X8 FILLER_21_45 ();
 FILLCELL_X1 FILLER_21_53 ();
 FILLCELL_X4 FILLER_21_58 ();
 FILLCELL_X8 FILLER_21_79 ();
 FILLCELL_X4 FILLER_21_87 ();
 FILLCELL_X1 FILLER_21_91 ();
 FILLCELL_X4 FILLER_21_122 ();
 FILLCELL_X2 FILLER_21_133 ();
 FILLCELL_X8 FILLER_21_153 ();
 FILLCELL_X1 FILLER_21_161 ();
 FILLCELL_X1 FILLER_21_192 ();
 FILLCELL_X1 FILLER_21_196 ();
 FILLCELL_X2 FILLER_21_200 ();
 FILLCELL_X4 FILLER_22_7 ();
 FILLCELL_X2 FILLER_22_11 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X2 FILLER_22_21 ();
 FILLCELL_X4 FILLER_22_57 ();
 FILLCELL_X1 FILLER_22_61 ();
 FILLCELL_X8 FILLER_22_95 ();
 FILLCELL_X4 FILLER_22_103 ();
 FILLCELL_X2 FILLER_22_107 ();
 FILLCELL_X4 FILLER_22_113 ();
 FILLCELL_X2 FILLER_22_124 ();
 FILLCELL_X1 FILLER_22_126 ();
 FILLCELL_X4 FILLER_22_144 ();
 FILLCELL_X2 FILLER_22_148 ();
 FILLCELL_X8 FILLER_22_167 ();
 FILLCELL_X2 FILLER_22_175 ();
 FILLCELL_X2 FILLER_22_181 ();
 FILLCELL_X1 FILLER_22_183 ();
 FILLCELL_X2 FILLER_22_191 ();
 FILLCELL_X1 FILLER_22_193 ();
 FILLCELL_X2 FILLER_22_197 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_40 ();
 FILLCELL_X1 FILLER_23_42 ();
 FILLCELL_X8 FILLER_23_57 ();
 FILLCELL_X4 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_75 ();
 FILLCELL_X4 FILLER_23_107 ();
 FILLCELL_X8 FILLER_23_128 ();
 FILLCELL_X2 FILLER_23_136 ();
 FILLCELL_X1 FILLER_23_138 ();
 FILLCELL_X4 FILLER_23_146 ();
 FILLCELL_X2 FILLER_23_150 ();
 FILLCELL_X1 FILLER_23_163 ();
 FILLCELL_X1 FILLER_23_185 ();
 FILLCELL_X1 FILLER_24_22 ();
 FILLCELL_X1 FILLER_24_30 ();
 FILLCELL_X1 FILLER_24_34 ();
 FILLCELL_X2 FILLER_24_42 ();
 FILLCELL_X1 FILLER_24_44 ();
 FILLCELL_X8 FILLER_24_85 ();
 FILLCELL_X1 FILLER_24_93 ();
 FILLCELL_X2 FILLER_24_115 ();
 FILLCELL_X2 FILLER_24_124 ();
 FILLCELL_X1 FILLER_24_126 ();
 FILLCELL_X1 FILLER_24_144 ();
 FILLCELL_X1 FILLER_24_151 ();
 FILLCELL_X1 FILLER_24_176 ();
 FILLCELL_X1 FILLER_24_180 ();
 FILLCELL_X1 FILLER_24_184 ();
 FILLCELL_X2 FILLER_25_7 ();
 FILLCELL_X1 FILLER_25_30 ();
 FILLCELL_X2 FILLER_25_55 ();
 FILLCELL_X2 FILLER_25_91 ();
 FILLCELL_X1 FILLER_25_100 ();
 FILLCELL_X1 FILLER_25_111 ();
 FILLCELL_X2 FILLER_25_132 ();
 FILLCELL_X2 FILLER_25_159 ();
 FILLCELL_X2 FILLER_25_184 ();
 FILLCELL_X2 FILLER_25_190 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_17 ();
 FILLCELL_X2 FILLER_26_41 ();
 FILLCELL_X2 FILLER_26_66 ();
 FILLCELL_X1 FILLER_26_87 ();
 FILLCELL_X1 FILLER_26_91 ();
 FILLCELL_X2 FILLER_26_98 ();
 FILLCELL_X4 FILLER_26_103 ();
 FILLCELL_X2 FILLER_26_107 ();
 FILLCELL_X8 FILLER_26_187 ();
 FILLCELL_X4 FILLER_26_195 ();
 FILLCELL_X2 FILLER_26_199 ();
 FILLCELL_X1 FILLER_26_201 ();
endmodule
