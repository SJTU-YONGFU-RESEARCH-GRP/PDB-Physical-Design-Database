module configurable_kogge_stone_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 INV_X1 _409_ (.A(net1),
    .ZN(_341_));
 INV_X1 _410_ (.A(net33),
    .ZN(_342_));
 INV_X1 _411_ (.A(net65),
    .ZN(_343_));
 INV_X1 _412_ (.A(_345_),
    .ZN(_000_));
 INV_X1 _413_ (.A(_346_),
    .ZN(_001_));
 CLKBUF_X3 _414_ (.A(_353_),
    .Z(_002_));
 BUF_X1 _415_ (.A(_355_),
    .Z(_003_));
 NOR2_X1 _416_ (.A1(_002_),
    .A2(_003_),
    .ZN(_004_));
 INV_X1 _417_ (.A(_357_),
    .ZN(_005_));
 BUF_X2 _418_ (.A(_358_),
    .Z(_006_));
 CLKBUF_X3 _419_ (.A(_360_),
    .Z(_007_));
 BUF_X2 _420_ (.A(_359_),
    .Z(_008_));
 OAI21_X1 _421_ (.A(_006_),
    .B1(_007_),
    .B2(_008_),
    .ZN(_009_));
 CLKBUF_X2 _422_ (.A(_361_),
    .Z(_010_));
 BUF_X4 _423_ (.A(_370_),
    .Z(_011_));
 AOI21_X2 _424_ (.A(_369_),
    .B1(_371_),
    .B2(_011_),
    .ZN(_012_));
 CLKBUF_X3 _425_ (.A(_372_),
    .Z(_013_));
 NAND2_X2 _426_ (.A1(_011_),
    .A2(_013_),
    .ZN(_014_));
 CLKBUF_X3 _427_ (.A(_374_),
    .Z(_015_));
 AOI21_X2 _428_ (.A(_373_),
    .B1(_375_),
    .B2(_015_),
    .ZN(_016_));
 OAI21_X2 _429_ (.A(_012_),
    .B1(_014_),
    .B2(_016_),
    .ZN(_017_));
 CLKBUF_X3 _430_ (.A(_366_),
    .Z(_018_));
 BUF_X4 _431_ (.A(_368_),
    .Z(_019_));
 NAND2_X2 _432_ (.A1(_018_),
    .A2(_019_),
    .ZN(_020_));
 BUF_X2 _433_ (.A(_362_),
    .Z(_021_));
 CLKBUF_X3 _434_ (.A(_364_),
    .Z(_022_));
 NAND2_X1 _435_ (.A1(_021_),
    .A2(_022_),
    .ZN(_023_));
 NOR2_X1 _436_ (.A1(_020_),
    .A2(_023_),
    .ZN(_024_));
 INV_X1 _437_ (.A(_363_),
    .ZN(_025_));
 AOI21_X1 _438_ (.A(_365_),
    .B1(_367_),
    .B2(_018_),
    .ZN(_026_));
 INV_X1 _439_ (.A(_022_),
    .ZN(_027_));
 OAI21_X1 _440_ (.A(_025_),
    .B1(_026_),
    .B2(_027_),
    .ZN(_028_));
 AOI221_X2 _441_ (.A(_010_),
    .B1(_017_),
    .B2(_024_),
    .C1(_028_),
    .C2(_021_),
    .ZN(_029_));
 NOR3_X1 _442_ (.A1(_014_),
    .A2(_020_),
    .A3(_023_),
    .ZN(_030_));
 NOR3_X1 _443_ (.A1(_357_),
    .A2(_008_),
    .A3(_030_),
    .ZN(_031_));
 AOI22_X2 _444_ (.A1(_005_),
    .A2(_009_),
    .B1(_029_),
    .B2(_031_),
    .ZN(_032_));
 INV_X1 _445_ (.A(_008_),
    .ZN(_033_));
 NAND3_X2 _446_ (.A1(_005_),
    .A2(_033_),
    .A3(_029_),
    .ZN(_034_));
 CLKBUF_X3 _447_ (.A(_376_),
    .Z(_035_));
 NAND2_X1 _448_ (.A1(_015_),
    .A2(_035_),
    .ZN(_036_));
 BUF_X2 _449_ (.A(_377_),
    .Z(_037_));
 BUF_X2 _450_ (.A(_379_),
    .Z(_038_));
 CLKBUF_X3 _451_ (.A(_378_),
    .Z(_039_));
 AOI21_X2 _452_ (.A(_037_),
    .B1(_038_),
    .B2(_039_),
    .ZN(_040_));
 NOR2_X1 _453_ (.A1(_036_),
    .A2(_040_),
    .ZN(_041_));
 CLKBUF_X3 _454_ (.A(_380_),
    .Z(_042_));
 AND4_X2 _455_ (.A1(_015_),
    .A2(_035_),
    .A3(_039_),
    .A4(_042_),
    .ZN(_043_));
 BUF_X2 _456_ (.A(_381_),
    .Z(_044_));
 AOI21_X2 _457_ (.A(_041_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_045_));
 CLKBUF_X3 _458_ (.A(_382_),
    .Z(_046_));
 AND2_X1 _459_ (.A1(_046_),
    .A2(_043_),
    .ZN(_047_));
 CLKBUF_X3 _460_ (.A(_398_),
    .Z(_048_));
 AOI21_X1 _461_ (.A(_397_),
    .B1(_399_),
    .B2(_048_),
    .ZN(_049_));
 CLKBUF_X3 _462_ (.A(_402_),
    .Z(_050_));
 CLKBUF_X3 _463_ (.A(_404_),
    .Z(_051_));
 NAND4_X1 _464_ (.A1(_050_),
    .A2(_048_),
    .A3(_400_),
    .A4(_051_),
    .ZN(_052_));
 BUF_X2 _465_ (.A(_406_),
    .Z(_053_));
 AOI21_X2 _466_ (.A(_405_),
    .B1(_407_),
    .B2(_053_),
    .ZN(_054_));
 NAND2_X1 _467_ (.A1(_048_),
    .A2(_400_),
    .ZN(_055_));
 AOI21_X2 _468_ (.A(_401_),
    .B1(_403_),
    .B2(_050_),
    .ZN(_056_));
 OAI221_X4 _469_ (.A(_049_),
    .B1(_052_),
    .B2(_054_),
    .C1(_055_),
    .C2(_056_),
    .ZN(_057_));
 CLKBUF_X3 _470_ (.A(_383_),
    .Z(_058_));
 NOR2_X1 _471_ (.A1(_058_),
    .A2(_385_),
    .ZN(_059_));
 BUF_X2 _472_ (.A(_391_),
    .Z(_060_));
 BUF_X2 _473_ (.A(_393_),
    .Z(_061_));
 CLKBUF_X3 _474_ (.A(_395_),
    .Z(_062_));
 CLKBUF_X3 _475_ (.A(_394_),
    .Z(_063_));
 AOI211_X2 _476_ (.A(_060_),
    .B(_061_),
    .C1(_062_),
    .C2(_063_),
    .ZN(_064_));
 CLKBUF_X3 _477_ (.A(_386_),
    .Z(_065_));
 INV_X2 _478_ (.A(_065_),
    .ZN(_066_));
 CLKBUF_X3 _479_ (.A(_389_),
    .Z(_067_));
 BUF_X4 _480_ (.A(_388_),
    .Z(_068_));
 AOI21_X2 _481_ (.A(_387_),
    .B1(_067_),
    .B2(_068_),
    .ZN(_069_));
 OAI211_X2 _482_ (.A(_059_),
    .B(_064_),
    .C1(_066_),
    .C2(_069_),
    .ZN(_070_));
 OAI21_X2 _483_ (.A(_047_),
    .B1(_057_),
    .B2(_070_),
    .ZN(_071_));
 BUF_X4 _484_ (.A(_384_),
    .Z(_072_));
 OAI21_X2 _485_ (.A(_059_),
    .B1(_069_),
    .B2(_066_),
    .ZN(_073_));
 NAND2_X1 _486_ (.A1(_065_),
    .A2(_068_),
    .ZN(_074_));
 BUF_X4 _487_ (.A(_390_),
    .Z(_075_));
 CLKBUF_X3 _488_ (.A(_392_),
    .Z(_076_));
 OAI21_X1 _489_ (.A(_075_),
    .B1(_076_),
    .B2(_060_),
    .ZN(_077_));
 CLKBUF_X3 _490_ (.A(_396_),
    .Z(_078_));
 OAI21_X1 _491_ (.A(_063_),
    .B1(_078_),
    .B2(_062_),
    .ZN(_079_));
 NOR2_X1 _492_ (.A1(_060_),
    .A2(_061_),
    .ZN(_080_));
 AOI211_X2 _493_ (.A(_074_),
    .B(_077_),
    .C1(_079_),
    .C2(_080_),
    .ZN(_081_));
 OAI22_X4 _494_ (.A1(_072_),
    .A2(_058_),
    .B1(_073_),
    .B2(_081_),
    .ZN(_082_));
 OAI21_X4 _495_ (.A(_045_),
    .B1(_071_),
    .B2(_082_),
    .ZN(_083_));
 OAI21_X4 _496_ (.A(_032_),
    .B1(_034_),
    .B2(_083_),
    .ZN(_084_));
 BUF_X2 _497_ (.A(_356_),
    .Z(_085_));
 INV_X2 _498_ (.A(_085_),
    .ZN(_086_));
 OAI21_X4 _499_ (.A(_004_),
    .B1(_084_),
    .B2(_086_),
    .ZN(_087_));
 CLKBUF_X3 _500_ (.A(_352_),
    .Z(_088_));
 AND3_X1 _501_ (.A1(_348_),
    .A2(_350_),
    .A3(_088_),
    .ZN(_089_));
 BUF_X4 _502_ (.A(_354_),
    .Z(_090_));
 OAI21_X1 _503_ (.A(_089_),
    .B1(_002_),
    .B2(_090_),
    .ZN(_091_));
 INV_X1 _504_ (.A(_091_),
    .ZN(_092_));
 INV_X1 _505_ (.A(_349_),
    .ZN(_093_));
 INV_X4 _506_ (.A(_351_),
    .ZN(_094_));
 INV_X1 _507_ (.A(_350_),
    .ZN(_095_));
 OAI21_X4 _508_ (.A(_093_),
    .B1(_094_),
    .B2(_095_),
    .ZN(_096_));
 AOI221_X2 _509_ (.A(_347_),
    .B1(_087_),
    .B2(_092_),
    .C1(_096_),
    .C2(_348_),
    .ZN(_097_));
 INV_X1 _510_ (.A(_003_),
    .ZN(_098_));
 OAI21_X1 _511_ (.A(_007_),
    .B1(_021_),
    .B2(_010_),
    .ZN(_099_));
 AOI21_X1 _512_ (.A(_363_),
    .B1(_365_),
    .B2(_022_),
    .ZN(_100_));
 AOI21_X2 _513_ (.A(_367_),
    .B1(_369_),
    .B2(_019_),
    .ZN(_101_));
 NAND2_X1 _514_ (.A1(_022_),
    .A2(_018_),
    .ZN(_102_));
 OAI21_X1 _515_ (.A(_100_),
    .B1(_101_),
    .B2(_102_),
    .ZN(_103_));
 NOR2_X1 _516_ (.A1(_010_),
    .A2(_103_),
    .ZN(_104_));
 NAND4_X4 _517_ (.A1(_022_),
    .A2(_018_),
    .A3(_019_),
    .A4(_011_),
    .ZN(_105_));
 AOI21_X4 _518_ (.A(_371_),
    .B1(_373_),
    .B2(_013_),
    .ZN(_106_));
 NOR2_X1 _519_ (.A1(_105_),
    .A2(_106_),
    .ZN(_107_));
 NAND2_X2 _520_ (.A1(_013_),
    .A2(_015_),
    .ZN(_108_));
 NOR2_X1 _521_ (.A1(_105_),
    .A2(_108_),
    .ZN(_109_));
 AOI21_X2 _522_ (.A(_375_),
    .B1(_037_),
    .B2(_035_),
    .ZN(_110_));
 NAND2_X1 _523_ (.A1(_035_),
    .A2(_039_),
    .ZN(_111_));
 AOI21_X2 _524_ (.A(_038_),
    .B1(_044_),
    .B2(_042_),
    .ZN(_112_));
 OAI21_X4 _525_ (.A(_110_),
    .B1(_111_),
    .B2(_112_),
    .ZN(_113_));
 AOI21_X1 _526_ (.A(_107_),
    .B1(_109_),
    .B2(_113_),
    .ZN(_114_));
 AOI21_X2 _527_ (.A(_099_),
    .B1(_104_),
    .B2(_114_),
    .ZN(_115_));
 AND2_X1 _528_ (.A1(_072_),
    .A2(_385_),
    .ZN(_116_));
 NOR2_X1 _529_ (.A1(_058_),
    .A2(_116_),
    .ZN(_117_));
 NAND2_X1 _530_ (.A1(_072_),
    .A2(_065_),
    .ZN(_118_));
 INV_X1 _531_ (.A(_387_),
    .ZN(_119_));
 OAI21_X1 _532_ (.A(_068_),
    .B1(_075_),
    .B2(_067_),
    .ZN(_120_));
 NAND2_X1 _533_ (.A1(_119_),
    .A2(_120_),
    .ZN(_121_));
 NOR3_X1 _534_ (.A1(_387_),
    .A2(_067_),
    .A3(_060_),
    .ZN(_122_));
 OAI21_X1 _535_ (.A(_076_),
    .B1(_063_),
    .B2(_061_),
    .ZN(_123_));
 AOI211_X2 _536_ (.A(_061_),
    .B(_062_),
    .C1(_397_),
    .C2(_078_),
    .ZN(_124_));
 OAI21_X2 _537_ (.A(_122_),
    .B1(_123_),
    .B2(_124_),
    .ZN(_125_));
 INV_X1 _538_ (.A(_399_),
    .ZN(_126_));
 NAND3_X4 _539_ (.A1(_050_),
    .A2(_400_),
    .A3(_051_),
    .ZN(_127_));
 INV_X1 _540_ (.A(_400_),
    .ZN(_128_));
 OAI221_X2 _541_ (.A(_126_),
    .B1(_054_),
    .B2(_127_),
    .C1(_056_),
    .C2(_128_),
    .ZN(_129_));
 NAND4_X4 _542_ (.A1(_076_),
    .A2(_063_),
    .A3(_078_),
    .A4(_048_),
    .ZN(_130_));
 AOI21_X2 _543_ (.A(_130_),
    .B1(_120_),
    .B2(_119_),
    .ZN(_131_));
 AOI22_X4 _544_ (.A1(_121_),
    .A2(_125_),
    .B1(_129_),
    .B2(_131_),
    .ZN(_132_));
 OAI21_X2 _545_ (.A(_117_),
    .B1(_118_),
    .B2(_132_),
    .ZN(_133_));
 NAND4_X2 _546_ (.A1(_035_),
    .A2(_039_),
    .A3(_042_),
    .A4(_046_),
    .ZN(_134_));
 NAND2_X1 _547_ (.A1(_019_),
    .A2(_011_),
    .ZN(_135_));
 NOR2_X1 _548_ (.A1(_135_),
    .A2(_108_),
    .ZN(_136_));
 NAND4_X2 _549_ (.A1(_007_),
    .A2(_021_),
    .A3(_022_),
    .A4(_018_),
    .ZN(_137_));
 INV_X1 _550_ (.A(_137_),
    .ZN(_138_));
 NAND2_X1 _551_ (.A1(_136_),
    .A2(_138_),
    .ZN(_139_));
 NOR2_X1 _552_ (.A1(_134_),
    .A2(_139_),
    .ZN(_140_));
 AOI211_X2 _553_ (.A(_008_),
    .B(_115_),
    .C1(_133_),
    .C2(_140_),
    .ZN(_141_));
 INV_X1 _554_ (.A(_044_),
    .ZN(_142_));
 OAI21_X2 _555_ (.A(_046_),
    .B1(_070_),
    .B2(_057_),
    .ZN(_143_));
 OAI21_X4 _556_ (.A(_142_),
    .B1(_082_),
    .B2(_143_),
    .ZN(_144_));
 NAND4_X4 _557_ (.A1(_019_),
    .A2(_011_),
    .A3(_013_),
    .A4(_015_),
    .ZN(_145_));
 NOR2_X1 _558_ (.A1(_145_),
    .A2(_137_),
    .ZN(_146_));
 OAI21_X2 _559_ (.A(_101_),
    .B1(_106_),
    .B2(_135_),
    .ZN(_147_));
 AOI22_X2 _560_ (.A1(_113_),
    .A2(_146_),
    .B1(_147_),
    .B2(_138_),
    .ZN(_148_));
 INV_X1 _561_ (.A(_002_),
    .ZN(_149_));
 NAND3_X1 _562_ (.A1(_094_),
    .A2(_149_),
    .A3(_033_),
    .ZN(_150_));
 INV_X1 _563_ (.A(_010_),
    .ZN(_151_));
 INV_X1 _564_ (.A(_021_),
    .ZN(_152_));
 OAI21_X1 _565_ (.A(_151_),
    .B1(_100_),
    .B2(_152_),
    .ZN(_153_));
 OAI21_X1 _566_ (.A(_098_),
    .B1(_005_),
    .B2(_086_),
    .ZN(_154_));
 AOI221_X2 _567_ (.A(_150_),
    .B1(_153_),
    .B2(_007_),
    .C1(_154_),
    .C2(_090_),
    .ZN(_155_));
 INV_X1 _568_ (.A(_090_),
    .ZN(_156_));
 OAI21_X1 _569_ (.A(_085_),
    .B1(_006_),
    .B2(_357_),
    .ZN(_157_));
 AOI21_X1 _570_ (.A(_156_),
    .B1(_098_),
    .B2(_157_),
    .ZN(_158_));
 OAI21_X1 _571_ (.A(_088_),
    .B1(_002_),
    .B2(_158_),
    .ZN(_159_));
 AOI22_X2 _572_ (.A1(_148_),
    .A2(_155_),
    .B1(_159_),
    .B2(_094_),
    .ZN(_160_));
 NAND4_X2 _573_ (.A1(_088_),
    .A2(_090_),
    .A3(_085_),
    .A4(_006_),
    .ZN(_161_));
 NOR4_X2 _574_ (.A1(_134_),
    .A2(_145_),
    .A3(_137_),
    .A4(_161_),
    .ZN(_162_));
 OAI21_X1 _575_ (.A(_162_),
    .B1(_116_),
    .B2(_058_),
    .ZN(_163_));
 NAND3_X1 _576_ (.A1(_072_),
    .A2(_065_),
    .A3(_162_),
    .ZN(_164_));
 OAI21_X2 _577_ (.A(_163_),
    .B1(_164_),
    .B2(_132_),
    .ZN(_165_));
 NAND2_X1 _578_ (.A1(_350_),
    .A2(_088_),
    .ZN(_166_));
 OAI21_X1 _579_ (.A(_090_),
    .B1(_085_),
    .B2(_003_),
    .ZN(_167_));
 AOI21_X1 _580_ (.A(_166_),
    .B1(_167_),
    .B2(_149_),
    .ZN(_168_));
 NOR3_X1 _581_ (.A1(_002_),
    .A2(_003_),
    .A3(_357_),
    .ZN(_169_));
 NAND2_X1 _582_ (.A1(_006_),
    .A2(_008_),
    .ZN(_170_));
 NAND2_X2 _583_ (.A1(_006_),
    .A2(_007_),
    .ZN(_171_));
 AOI21_X1 _584_ (.A(_010_),
    .B1(_363_),
    .B2(_021_),
    .ZN(_172_));
 OAI211_X2 _585_ (.A(_169_),
    .B(_170_),
    .C1(_171_),
    .C2(_172_),
    .ZN(_173_));
 AOI21_X1 _586_ (.A(_096_),
    .B1(_168_),
    .B2(_173_),
    .ZN(_174_));
 NOR2_X1 _587_ (.A1(_023_),
    .A2(_171_),
    .ZN(_175_));
 NAND2_X1 _588_ (.A1(_168_),
    .A2(_175_),
    .ZN(_176_));
 OAI21_X1 _589_ (.A(_026_),
    .B1(_012_),
    .B2(_020_),
    .ZN(_177_));
 OAI21_X2 _590_ (.A(_016_),
    .B1(_036_),
    .B2(_040_),
    .ZN(_178_));
 NOR2_X2 _591_ (.A1(_014_),
    .A2(_020_),
    .ZN(_179_));
 AOI21_X2 _592_ (.A(_177_),
    .B1(_178_),
    .B2(_179_),
    .ZN(_180_));
 OAI21_X1 _593_ (.A(_174_),
    .B1(_176_),
    .B2(_180_),
    .ZN(_181_));
 NOR4_X2 _594_ (.A1(_144_),
    .A2(_160_),
    .A3(_165_),
    .A4(_181_),
    .ZN(_182_));
 NAND4_X2 _595_ (.A1(_098_),
    .A2(_084_),
    .A3(_141_),
    .A4(_182_),
    .ZN(_183_));
 AND4_X2 _596_ (.A1(_035_),
    .A2(_039_),
    .A3(_042_),
    .A4(_046_),
    .ZN(_184_));
 NAND2_X2 _597_ (.A1(_053_),
    .A2(_408_),
    .ZN(_185_));
 NAND4_X2 _598_ (.A1(_072_),
    .A2(_065_),
    .A3(_068_),
    .A4(_075_),
    .ZN(_186_));
 NOR4_X4 _599_ (.A1(_127_),
    .A2(_130_),
    .A3(_185_),
    .A4(_186_),
    .ZN(_187_));
 NAND2_X4 _600_ (.A1(_184_),
    .A2(_187_),
    .ZN(_188_));
 NOR2_X2 _601_ (.A1(_139_),
    .A2(_188_),
    .ZN(_189_));
 INV_X1 _602_ (.A(_180_),
    .ZN(_190_));
 AND2_X1 _603_ (.A1(_043_),
    .A2(_179_),
    .ZN(_191_));
 AOI211_X2 _604_ (.A(_147_),
    .B(_190_),
    .C1(_191_),
    .C2(_144_),
    .ZN(_192_));
 INV_X1 _605_ (.A(_014_),
    .ZN(_193_));
 AOI21_X4 _606_ (.A(_017_),
    .B1(_083_),
    .B2(_193_),
    .ZN(_194_));
 INV_X1 _607_ (.A(_385_),
    .ZN(_195_));
 OAI21_X4 _608_ (.A(_195_),
    .B1(_132_),
    .B2(_066_),
    .ZN(_196_));
 AND2_X2 _609_ (.A1(_063_),
    .A2(_078_),
    .ZN(_197_));
 NOR2_X2 _610_ (.A1(_127_),
    .A2(_185_),
    .ZN(_198_));
 NAND3_X2 _611_ (.A1(_048_),
    .A2(_197_),
    .A3(_198_),
    .ZN(_199_));
 NAND2_X1 _612_ (.A1(_050_),
    .A2(_403_),
    .ZN(_200_));
 NAND3_X1 _613_ (.A1(_050_),
    .A2(_051_),
    .A3(_405_),
    .ZN(_201_));
 NAND2_X1 _614_ (.A1(_200_),
    .A2(_201_),
    .ZN(_202_));
 OR3_X1 _615_ (.A1(_062_),
    .A2(_399_),
    .A3(_401_),
    .ZN(_203_));
 INV_X1 _616_ (.A(_407_),
    .ZN(_204_));
 INV_X1 _617_ (.A(_408_),
    .ZN(_205_));
 OAI21_X2 _618_ (.A(_204_),
    .B1(_344_),
    .B2(_205_),
    .ZN(_206_));
 NAND3_X2 _619_ (.A1(_050_),
    .A2(_053_),
    .A3(_051_),
    .ZN(_207_));
 INV_X1 _620_ (.A(_207_),
    .ZN(_208_));
 AOI211_X2 _621_ (.A(_202_),
    .B(_203_),
    .C1(_206_),
    .C2(_208_),
    .ZN(_209_));
 INV_X1 _622_ (.A(_057_),
    .ZN(_210_));
 AOI21_X4 _623_ (.A(_199_),
    .B1(_209_),
    .B2(_210_),
    .ZN(_211_));
 INV_X2 _624_ (.A(_067_),
    .ZN(_212_));
 NAND2_X1 _625_ (.A1(_063_),
    .A2(_062_),
    .ZN(_213_));
 NAND2_X1 _626_ (.A1(_080_),
    .A2(_213_),
    .ZN(_214_));
 AOI21_X4 _627_ (.A(_214_),
    .B1(_057_),
    .B2(_197_),
    .ZN(_215_));
 NOR2_X1 _628_ (.A1(_044_),
    .A2(_058_),
    .ZN(_216_));
 NAND4_X2 _629_ (.A1(_212_),
    .A2(_132_),
    .A3(_215_),
    .A4(_216_),
    .ZN(_217_));
 NOR3_X4 _630_ (.A1(_196_),
    .A2(_211_),
    .A3(_217_),
    .ZN(_218_));
 AND2_X1 _631_ (.A1(_046_),
    .A2(_187_),
    .ZN(_219_));
 NAND3_X2 _632_ (.A1(_193_),
    .A2(_043_),
    .A3(_219_),
    .ZN(_220_));
 OAI211_X4 _633_ (.A(_192_),
    .B(_194_),
    .C1(_218_),
    .C2(_220_),
    .ZN(_221_));
 AOI21_X4 _634_ (.A(_183_),
    .B1(_189_),
    .B2(_221_),
    .ZN(_222_));
 OR2_X1 _635_ (.A1(_108_),
    .A2(_188_),
    .ZN(_223_));
 NAND2_X1 _636_ (.A1(_085_),
    .A2(_021_),
    .ZN(_224_));
 NOR4_X4 _637_ (.A1(_105_),
    .A2(_171_),
    .A3(_223_),
    .A4(_224_),
    .ZN(_225_));
 NAND3_X1 _638_ (.A1(_090_),
    .A2(_089_),
    .A3(_225_),
    .ZN(_226_));
 OR2_X1 _639_ (.A1(_001_),
    .A2(_226_),
    .ZN(_227_));
 OAI221_X1 _640_ (.A(_000_),
    .B1(_001_),
    .B2(_097_),
    .C1(_222_),
    .C2(_227_),
    .ZN(net66));
 AND3_X2 _641_ (.A1(_048_),
    .A2(_197_),
    .A3(_198_),
    .ZN(_228_));
 AND2_X1 _642_ (.A1(_200_),
    .A2(_201_),
    .ZN(_229_));
 NOR2_X1 _643_ (.A1(_399_),
    .A2(_401_),
    .ZN(_230_));
 INV_X1 _644_ (.A(_344_),
    .ZN(_231_));
 AOI21_X2 _645_ (.A(_407_),
    .B1(_231_),
    .B2(_408_),
    .ZN(_232_));
 OAI211_X4 _646_ (.A(_229_),
    .B(_230_),
    .C1(_232_),
    .C2(_207_),
    .ZN(_233_));
 OR2_X1 _647_ (.A1(_062_),
    .A2(_057_),
    .ZN(_234_));
 OAI21_X2 _648_ (.A(_228_),
    .B1(_233_),
    .B2(_234_),
    .ZN(_235_));
 NAND3_X2 _649_ (.A1(_075_),
    .A2(_076_),
    .A3(_228_),
    .ZN(_236_));
 OR2_X1 _650_ (.A1(_077_),
    .A2(_215_),
    .ZN(_237_));
 AOI22_X2 _651_ (.A1(_235_),
    .A2(_215_),
    .B1(_236_),
    .B2(_237_),
    .ZN(_238_));
 NOR2_X2 _652_ (.A1(_067_),
    .A2(_238_),
    .ZN(_239_));
 XNOR2_X2 _653_ (.A(_068_),
    .B(_239_),
    .ZN(net68));
 NAND4_X2 _654_ (.A1(_068_),
    .A2(_075_),
    .A3(_076_),
    .A4(_228_),
    .ZN(_240_));
 OAI21_X4 _655_ (.A(_132_),
    .B1(_239_),
    .B2(_240_),
    .ZN(_241_));
 XNOR2_X2 _656_ (.A(_066_),
    .B(_241_),
    .ZN(net69));
 AND2_X1 _657_ (.A1(_048_),
    .A2(_198_),
    .ZN(_242_));
 AOI21_X2 _658_ (.A(_234_),
    .B1(_233_),
    .B2(_242_),
    .ZN(_243_));
 AND3_X1 _659_ (.A1(_212_),
    .A2(_132_),
    .A3(_215_),
    .ZN(_244_));
 AOI211_X2 _660_ (.A(_074_),
    .B(_236_),
    .C1(_243_),
    .C2(_244_),
    .ZN(_245_));
 NOR2_X1 _661_ (.A1(_196_),
    .A2(_245_),
    .ZN(_246_));
 XNOR2_X2 _662_ (.A(_072_),
    .B(_246_),
    .ZN(net70));
 AOI21_X2 _663_ (.A(_058_),
    .B1(_196_),
    .B2(_072_),
    .ZN(_247_));
 INV_X1 _664_ (.A(_187_),
    .ZN(_248_));
 OAI21_X1 _665_ (.A(_247_),
    .B1(_248_),
    .B2(_246_),
    .ZN(_249_));
 XOR2_X2 _666_ (.A(_046_),
    .B(_249_),
    .Z(net71));
 INV_X1 _667_ (.A(_144_),
    .ZN(_250_));
 NAND2_X1 _668_ (.A1(_046_),
    .A2(_187_),
    .ZN(_251_));
 NOR3_X2 _669_ (.A1(_058_),
    .A2(_196_),
    .A3(_245_),
    .ZN(_252_));
 OAI21_X2 _670_ (.A(_250_),
    .B1(_251_),
    .B2(_252_),
    .ZN(_253_));
 XOR2_X2 _671_ (.A(_042_),
    .B(_253_),
    .Z(net72));
 AOI21_X2 _672_ (.A(_038_),
    .B1(_253_),
    .B2(_042_),
    .ZN(_254_));
 XNOR2_X2 _673_ (.A(_039_),
    .B(_254_),
    .ZN(net73));
 NOR3_X1 _674_ (.A1(_037_),
    .A2(_038_),
    .A3(_144_),
    .ZN(_255_));
 OAI21_X1 _675_ (.A(_255_),
    .B1(_252_),
    .B2(_251_),
    .ZN(_256_));
 OR2_X1 _676_ (.A1(_042_),
    .A2(_037_),
    .ZN(_257_));
 OAI221_X2 _677_ (.A(_256_),
    .B1(_257_),
    .B2(_038_),
    .C1(_037_),
    .C2(_039_),
    .ZN(_258_));
 XNOR2_X2 _678_ (.A(_035_),
    .B(_258_),
    .ZN(net74));
 AND2_X1 _679_ (.A1(_046_),
    .A2(_058_),
    .ZN(_259_));
 NOR4_X1 _680_ (.A1(_044_),
    .A2(_196_),
    .A3(_259_),
    .A4(_245_),
    .ZN(_260_));
 OAI21_X1 _681_ (.A(_247_),
    .B1(_248_),
    .B2(_260_),
    .ZN(_261_));
 INV_X1 _682_ (.A(_188_),
    .ZN(_262_));
 AOI221_X2 _683_ (.A(_113_),
    .B1(_184_),
    .B2(_261_),
    .C1(_262_),
    .C2(_144_),
    .ZN(_263_));
 XNOR2_X2 _684_ (.A(_015_),
    .B(_263_),
    .ZN(net75));
 OR2_X1 _685_ (.A1(_178_),
    .A2(_219_),
    .ZN(_264_));
 OAI22_X1 _686_ (.A1(_043_),
    .A2(_178_),
    .B1(_264_),
    .B2(_144_),
    .ZN(_265_));
 NOR3_X1 _687_ (.A1(_144_),
    .A2(_113_),
    .A3(_178_),
    .ZN(_266_));
 OR3_X1 _688_ (.A1(_058_),
    .A2(_144_),
    .A3(_196_),
    .ZN(_267_));
 OAI21_X1 _689_ (.A(_184_),
    .B1(_245_),
    .B2(_267_),
    .ZN(_268_));
 AOI21_X2 _690_ (.A(_265_),
    .B1(_266_),
    .B2(_268_),
    .ZN(_269_));
 XOR2_X2 _691_ (.A(_013_),
    .B(_269_),
    .Z(net76));
 AOI21_X1 _692_ (.A(_113_),
    .B1(_133_),
    .B2(_184_),
    .ZN(_270_));
 OAI21_X2 _693_ (.A(_106_),
    .B1(_108_),
    .B2(_270_),
    .ZN(_271_));
 NOR2_X1 _694_ (.A1(_108_),
    .A2(_188_),
    .ZN(_272_));
 AOI21_X2 _695_ (.A(_271_),
    .B1(_269_),
    .B2(_272_),
    .ZN(_273_));
 XNOR2_X2 _696_ (.A(_011_),
    .B(_273_),
    .ZN(net77));
 XNOR2_X1 _697_ (.A(_053_),
    .B(_344_),
    .ZN(net78));
 OAI21_X1 _698_ (.A(_194_),
    .B1(_218_),
    .B2(_220_),
    .ZN(_274_));
 XOR2_X2 _699_ (.A(_019_),
    .B(_274_),
    .Z(net79));
 NOR2_X1 _700_ (.A1(_134_),
    .A2(_145_),
    .ZN(_275_));
 AOI221_X2 _701_ (.A(_147_),
    .B1(_275_),
    .B2(_133_),
    .C1(_136_),
    .C2(_113_),
    .ZN(_276_));
 NOR3_X2 _702_ (.A1(_145_),
    .A2(_188_),
    .A3(_194_),
    .ZN(_277_));
 NOR4_X2 _703_ (.A1(_145_),
    .A2(_188_),
    .A3(_218_),
    .A4(_220_),
    .ZN(_278_));
 NOR2_X1 _704_ (.A1(_277_),
    .A2(_278_),
    .ZN(_279_));
 NAND2_X1 _705_ (.A1(_276_),
    .A2(_279_),
    .ZN(_280_));
 XOR2_X2 _706_ (.A(_018_),
    .B(_280_),
    .Z(net80));
 NAND2_X2 _707_ (.A1(_043_),
    .A2(_179_),
    .ZN(_281_));
 NOR2_X1 _708_ (.A1(_281_),
    .A2(_251_),
    .ZN(_282_));
 OAI21_X1 _709_ (.A(_180_),
    .B1(_281_),
    .B2(_250_),
    .ZN(_283_));
 OAI21_X1 _710_ (.A(_221_),
    .B1(_282_),
    .B2(_283_),
    .ZN(_284_));
 XNOR2_X2 _711_ (.A(_022_),
    .B(_284_),
    .ZN(net81));
 INV_X1 _712_ (.A(_103_),
    .ZN(_285_));
 AOI21_X1 _713_ (.A(_190_),
    .B1(_191_),
    .B2(_144_),
    .ZN(_286_));
 NAND2_X1 _714_ (.A1(_286_),
    .A2(_276_),
    .ZN(_287_));
 NOR4_X2 _715_ (.A1(_287_),
    .A2(_271_),
    .A3(_277_),
    .A4(_278_),
    .ZN(_288_));
 INV_X1 _716_ (.A(_105_),
    .ZN(_289_));
 INV_X1 _717_ (.A(_282_),
    .ZN(_290_));
 AOI21_X1 _718_ (.A(_223_),
    .B1(_290_),
    .B2(_286_),
    .ZN(_291_));
 OAI21_X1 _719_ (.A(_289_),
    .B1(_271_),
    .B2(_291_),
    .ZN(_292_));
 OAI21_X1 _720_ (.A(_285_),
    .B1(_288_),
    .B2(_292_),
    .ZN(_293_));
 XNOR2_X2 _721_ (.A(_152_),
    .B(_293_),
    .ZN(net82));
 INV_X1 _722_ (.A(_029_),
    .ZN(_294_));
 AOI21_X1 _723_ (.A(_294_),
    .B1(_083_),
    .B2(_030_),
    .ZN(_295_));
 NOR2_X1 _724_ (.A1(_023_),
    .A2(_290_),
    .ZN(_296_));
 OAI21_X1 _725_ (.A(_296_),
    .B1(_291_),
    .B2(_271_),
    .ZN(_297_));
 OAI21_X1 _726_ (.A(_295_),
    .B1(_288_),
    .B2(_297_),
    .ZN(_298_));
 XOR2_X2 _727_ (.A(_007_),
    .B(_298_),
    .Z(net83));
 NOR2_X1 _728_ (.A1(_008_),
    .A2(_115_),
    .ZN(_299_));
 NAND2_X1 _729_ (.A1(_184_),
    .A2(_146_),
    .ZN(_300_));
 OAI21_X2 _730_ (.A(_299_),
    .B1(_247_),
    .B2(_300_),
    .ZN(_301_));
 AOI21_X2 _731_ (.A(_301_),
    .B1(_189_),
    .B2(_221_),
    .ZN(_302_));
 XNOR2_X2 _732_ (.A(_006_),
    .B(_302_),
    .ZN(net84));
 NAND2_X1 _733_ (.A1(_175_),
    .A2(_282_),
    .ZN(_303_));
 OAI21_X1 _734_ (.A(_084_),
    .B1(_302_),
    .B2(_303_),
    .ZN(_304_));
 XNOR2_X2 _735_ (.A(_086_),
    .B(_304_),
    .ZN(net85));
 NAND2_X1 _736_ (.A1(_098_),
    .A2(_084_),
    .ZN(_305_));
 AOI211_X2 _737_ (.A(_305_),
    .B(_301_),
    .C1(_189_),
    .C2(_221_),
    .ZN(_306_));
 NOR2_X1 _738_ (.A1(_086_),
    .A2(_084_),
    .ZN(_307_));
 OR2_X1 _739_ (.A1(_003_),
    .A2(_225_),
    .ZN(_308_));
 NOR2_X1 _740_ (.A1(_307_),
    .A2(_308_),
    .ZN(_309_));
 NOR2_X1 _741_ (.A1(_306_),
    .A2(_309_),
    .ZN(_310_));
 XNOR2_X2 _742_ (.A(_156_),
    .B(_310_),
    .ZN(net86));
 OAI21_X1 _743_ (.A(_087_),
    .B1(_002_),
    .B2(_090_),
    .ZN(_311_));
 NAND2_X1 _744_ (.A1(_090_),
    .A2(_085_),
    .ZN(_312_));
 INV_X1 _745_ (.A(_175_),
    .ZN(_313_));
 NOR3_X1 _746_ (.A1(_312_),
    .A2(_313_),
    .A3(_290_),
    .ZN(_314_));
 OAI21_X1 _747_ (.A(_314_),
    .B1(_308_),
    .B2(_307_),
    .ZN(_315_));
 OAI21_X1 _748_ (.A(_311_),
    .B1(_306_),
    .B2(_315_),
    .ZN(_316_));
 XOR2_X2 _749_ (.A(_088_),
    .B(_316_),
    .Z(net87));
 NOR2_X1 _750_ (.A1(_160_),
    .A2(_165_),
    .ZN(_317_));
 OR3_X2 _751_ (.A1(_300_),
    .A2(_161_),
    .A3(_248_),
    .ZN(_318_));
 OAI21_X4 _752_ (.A(_317_),
    .B1(_306_),
    .B2(_318_),
    .ZN(_319_));
 XNOR2_X1 _753_ (.A(_095_),
    .B(_319_),
    .ZN(net88));
 AOI21_X1 _754_ (.A(_405_),
    .B1(_206_),
    .B2(_053_),
    .ZN(_320_));
 XNOR2_X1 _755_ (.A(_051_),
    .B(_320_),
    .ZN(net89));
 NOR4_X2 _756_ (.A1(_166_),
    .A2(_312_),
    .A3(_313_),
    .A4(_281_),
    .ZN(_321_));
 OAI21_X2 _757_ (.A(_321_),
    .B1(_219_),
    .B2(_144_),
    .ZN(_322_));
 OR2_X1 _758_ (.A1(_180_),
    .A2(_176_),
    .ZN(_323_));
 AND2_X1 _759_ (.A1(_323_),
    .A2(_174_),
    .ZN(_324_));
 AOI21_X4 _760_ (.A(_222_),
    .B1(_322_),
    .B2(_324_),
    .ZN(_325_));
 XOR2_X1 _761_ (.A(_348_),
    .B(_325_),
    .Z(net90));
 OAI21_X1 _762_ (.A(_097_),
    .B1(_222_),
    .B2(_226_),
    .ZN(_326_));
 XNOR2_X1 _763_ (.A(_001_),
    .B(_326_),
    .ZN(net91));
 OAI21_X1 _764_ (.A(_229_),
    .B1(_207_),
    .B2(_232_),
    .ZN(_327_));
 NOR2_X1 _765_ (.A1(_050_),
    .A2(_403_),
    .ZN(_328_));
 INV_X1 _766_ (.A(_051_),
    .ZN(_329_));
 OR2_X1 _767_ (.A1(_329_),
    .A2(_320_),
    .ZN(_330_));
 AOI21_X1 _768_ (.A(_327_),
    .B1(_328_),
    .B2(_330_),
    .ZN(net92));
 OR2_X1 _769_ (.A1(_401_),
    .A2(_327_),
    .ZN(_331_));
 XNOR2_X1 _770_ (.A(_128_),
    .B(_331_),
    .ZN(net93));
 AOI21_X1 _771_ (.A(_129_),
    .B1(_198_),
    .B2(_331_),
    .ZN(_332_));
 XNOR2_X1 _772_ (.A(_048_),
    .B(_332_),
    .ZN(net94));
 NAND2_X1 _773_ (.A1(_242_),
    .A2(_233_),
    .ZN(_333_));
 NAND2_X1 _774_ (.A1(_210_),
    .A2(_333_),
    .ZN(_334_));
 XOR2_X1 _775_ (.A(_078_),
    .B(_334_),
    .Z(net95));
 AOI21_X1 _776_ (.A(_062_),
    .B1(_334_),
    .B2(_078_),
    .ZN(_335_));
 XNOR2_X1 _777_ (.A(_063_),
    .B(_335_),
    .ZN(net96));
 AOI221_X1 _778_ (.A(_061_),
    .B1(_057_),
    .B2(_197_),
    .C1(_062_),
    .C2(_063_),
    .ZN(_336_));
 NAND2_X1 _779_ (.A1(_235_),
    .A2(_336_),
    .ZN(_337_));
 XOR2_X1 _780_ (.A(_076_),
    .B(_337_),
    .Z(net97));
 INV_X1 _781_ (.A(_060_),
    .ZN(_338_));
 AOI21_X1 _782_ (.A(_129_),
    .B1(_198_),
    .B2(_337_),
    .ZN(_339_));
 OAI221_X1 _783_ (.A(_338_),
    .B1(_124_),
    .B2(_123_),
    .C1(_130_),
    .C2(_339_),
    .ZN(_340_));
 XOR2_X1 _784_ (.A(_075_),
    .B(_340_),
    .Z(net98));
 FA_X1 _785_ (.A(_341_),
    .B(_342_),
    .CI(_343_),
    .CO(_344_),
    .S(net67));
 HA_X1 _786_ (.A(net25),
    .B(net57),
    .CO(_345_),
    .S(_346_));
 HA_X1 _787_ (.A(net24),
    .B(net56),
    .CO(_347_),
    .S(_348_));
 HA_X1 _788_ (.A(net22),
    .B(net54),
    .CO(_349_),
    .S(_350_));
 HA_X1 _789_ (.A(net21),
    .B(net53),
    .CO(_351_),
    .S(_352_));
 HA_X1 _790_ (.A(net20),
    .B(net52),
    .CO(_353_),
    .S(_354_));
 HA_X1 _791_ (.A(net19),
    .B(net51),
    .CO(_355_),
    .S(_356_));
 HA_X1 _792_ (.A(net18),
    .B(net50),
    .CO(_357_),
    .S(_358_));
 HA_X1 _793_ (.A(net17),
    .B(net49),
    .CO(_359_),
    .S(_360_));
 HA_X1 _794_ (.A(net16),
    .B(net48),
    .CO(_361_),
    .S(_362_));
 HA_X1 _795_ (.A(net15),
    .B(net47),
    .CO(_363_),
    .S(_364_));
 HA_X1 _796_ (.A(net14),
    .B(net46),
    .CO(_365_),
    .S(_366_));
 HA_X1 _797_ (.A(net13),
    .B(net45),
    .CO(_367_),
    .S(_368_));
 HA_X1 _798_ (.A(net11),
    .B(net43),
    .CO(_369_),
    .S(_370_));
 HA_X1 _799_ (.A(net10),
    .B(net42),
    .CO(_371_),
    .S(_372_));
 HA_X1 _800_ (.A(net9),
    .B(net41),
    .CO(_373_),
    .S(_374_));
 HA_X1 _801_ (.A(net8),
    .B(net40),
    .CO(_375_),
    .S(_376_));
 HA_X1 _802_ (.A(net7),
    .B(net39),
    .CO(_377_),
    .S(_378_));
 HA_X1 _803_ (.A(net6),
    .B(net38),
    .CO(_379_),
    .S(_380_));
 HA_X1 _804_ (.A(net5),
    .B(net37),
    .CO(_381_),
    .S(_382_));
 HA_X1 _805_ (.A(net4),
    .B(net36),
    .CO(_383_),
    .S(_384_));
 HA_X1 _806_ (.A(net3),
    .B(net35),
    .CO(_385_),
    .S(_386_));
 HA_X1 _807_ (.A(net2),
    .B(net34),
    .CO(_387_),
    .S(_388_));
 HA_X1 _808_ (.A(net32),
    .B(net64),
    .CO(_389_),
    .S(_390_));
 HA_X1 _809_ (.A(net31),
    .B(net63),
    .CO(_391_),
    .S(_392_));
 HA_X1 _810_ (.A(net30),
    .B(net62),
    .CO(_393_),
    .S(_394_));
 HA_X1 _811_ (.A(net29),
    .B(net61),
    .CO(_395_),
    .S(_396_));
 HA_X1 _812_ (.A(net28),
    .B(net60),
    .CO(_397_),
    .S(_398_));
 HA_X1 _813_ (.A(net27),
    .B(net59),
    .CO(_399_),
    .S(_400_));
 HA_X1 _814_ (.A(net26),
    .B(net58),
    .CO(_401_),
    .S(_402_));
 HA_X1 _815_ (.A(net23),
    .B(net55),
    .CO(_403_),
    .S(_404_));
 HA_X1 _816_ (.A(net12),
    .B(net44),
    .CO(_405_),
    .S(_406_));
 HA_X1 _817_ (.A(net1),
    .B(net33),
    .CO(_407_),
    .S(_408_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_658 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 BUF_X2 input2 (.A(a[10]),
    .Z(net2));
 BUF_X2 input3 (.A(a[11]),
    .Z(net3));
 BUF_X2 input4 (.A(a[12]),
    .Z(net4));
 BUF_X2 input5 (.A(a[13]),
    .Z(net5));
 BUF_X2 input6 (.A(a[14]),
    .Z(net6));
 BUF_X2 input7 (.A(a[15]),
    .Z(net7));
 BUF_X2 input8 (.A(a[16]),
    .Z(net8));
 BUF_X2 input9 (.A(a[17]),
    .Z(net9));
 BUF_X2 input10 (.A(a[18]),
    .Z(net10));
 BUF_X2 input11 (.A(a[19]),
    .Z(net11));
 BUF_X1 input12 (.A(a[1]),
    .Z(net12));
 BUF_X2 input13 (.A(a[20]),
    .Z(net13));
 BUF_X2 input14 (.A(a[21]),
    .Z(net14));
 BUF_X2 input15 (.A(a[22]),
    .Z(net15));
 BUF_X2 input16 (.A(a[23]),
    .Z(net16));
 BUF_X2 input17 (.A(a[24]),
    .Z(net17));
 BUF_X2 input18 (.A(a[25]),
    .Z(net18));
 BUF_X2 input19 (.A(a[26]),
    .Z(net19));
 BUF_X1 input20 (.A(a[27]),
    .Z(net20));
 BUF_X1 input21 (.A(a[28]),
    .Z(net21));
 BUF_X1 input22 (.A(a[29]),
    .Z(net22));
 BUF_X1 input23 (.A(a[2]),
    .Z(net23));
 BUF_X1 input24 (.A(a[30]),
    .Z(net24));
 BUF_X1 input25 (.A(a[31]),
    .Z(net25));
 BUF_X1 input26 (.A(a[3]),
    .Z(net26));
 BUF_X1 input27 (.A(a[4]),
    .Z(net27));
 BUF_X1 input28 (.A(a[5]),
    .Z(net28));
 BUF_X1 input29 (.A(a[6]),
    .Z(net29));
 BUF_X1 input30 (.A(a[7]),
    .Z(net30));
 BUF_X1 input31 (.A(a[8]),
    .Z(net31));
 BUF_X2 input32 (.A(a[9]),
    .Z(net32));
 BUF_X1 input33 (.A(b[0]),
    .Z(net33));
 BUF_X2 input34 (.A(b[10]),
    .Z(net34));
 BUF_X2 input35 (.A(b[11]),
    .Z(net35));
 BUF_X2 input36 (.A(b[12]),
    .Z(net36));
 BUF_X2 input37 (.A(b[13]),
    .Z(net37));
 BUF_X2 input38 (.A(b[14]),
    .Z(net38));
 BUF_X2 input39 (.A(b[15]),
    .Z(net39));
 BUF_X2 input40 (.A(b[16]),
    .Z(net40));
 BUF_X2 input41 (.A(b[17]),
    .Z(net41));
 BUF_X2 input42 (.A(b[18]),
    .Z(net42));
 BUF_X2 input43 (.A(b[19]),
    .Z(net43));
 BUF_X1 input44 (.A(b[1]),
    .Z(net44));
 BUF_X2 input45 (.A(b[20]),
    .Z(net45));
 BUF_X2 input46 (.A(b[21]),
    .Z(net46));
 BUF_X2 input47 (.A(b[22]),
    .Z(net47));
 BUF_X2 input48 (.A(b[23]),
    .Z(net48));
 BUF_X2 input49 (.A(b[24]),
    .Z(net49));
 BUF_X2 input50 (.A(b[25]),
    .Z(net50));
 BUF_X2 input51 (.A(b[26]),
    .Z(net51));
 BUF_X1 input52 (.A(b[27]),
    .Z(net52));
 BUF_X1 input53 (.A(b[28]),
    .Z(net53));
 BUF_X1 input54 (.A(b[29]),
    .Z(net54));
 BUF_X1 input55 (.A(b[2]),
    .Z(net55));
 BUF_X1 input56 (.A(b[30]),
    .Z(net56));
 BUF_X1 input57 (.A(b[31]),
    .Z(net57));
 BUF_X1 input58 (.A(b[3]),
    .Z(net58));
 BUF_X1 input59 (.A(b[4]),
    .Z(net59));
 BUF_X1 input60 (.A(b[5]),
    .Z(net60));
 BUF_X1 input61 (.A(b[6]),
    .Z(net61));
 BUF_X1 input62 (.A(b[7]),
    .Z(net62));
 BUF_X1 input63 (.A(b[8]),
    .Z(net63));
 BUF_X2 input64 (.A(b[9]),
    .Z(net64));
 BUF_X1 input65 (.A(cin),
    .Z(net65));
 BUF_X1 output66 (.A(net66),
    .Z(cout));
 BUF_X1 output67 (.A(net67),
    .Z(sum[0]));
 BUF_X1 output68 (.A(net68),
    .Z(sum[10]));
 BUF_X1 output69 (.A(net69),
    .Z(sum[11]));
 BUF_X1 output70 (.A(net70),
    .Z(sum[12]));
 BUF_X1 output71 (.A(net71),
    .Z(sum[13]));
 BUF_X1 output72 (.A(net72),
    .Z(sum[14]));
 BUF_X1 output73 (.A(net73),
    .Z(sum[15]));
 BUF_X1 output74 (.A(net74),
    .Z(sum[16]));
 BUF_X1 output75 (.A(net75),
    .Z(sum[17]));
 BUF_X1 output76 (.A(net76),
    .Z(sum[18]));
 BUF_X1 output77 (.A(net77),
    .Z(sum[19]));
 BUF_X1 output78 (.A(net78),
    .Z(sum[1]));
 BUF_X1 output79 (.A(net79),
    .Z(sum[20]));
 BUF_X1 output80 (.A(net80),
    .Z(sum[21]));
 BUF_X1 output81 (.A(net81),
    .Z(sum[22]));
 BUF_X1 output82 (.A(net82),
    .Z(sum[23]));
 BUF_X1 output83 (.A(net83),
    .Z(sum[24]));
 BUF_X1 output84 (.A(net84),
    .Z(sum[25]));
 BUF_X1 output85 (.A(net85),
    .Z(sum[26]));
 BUF_X1 output86 (.A(net86),
    .Z(sum[27]));
 BUF_X1 output87 (.A(net87),
    .Z(sum[28]));
 BUF_X1 output88 (.A(net88),
    .Z(sum[29]));
 BUF_X1 output89 (.A(net89),
    .Z(sum[2]));
 BUF_X1 output90 (.A(net90),
    .Z(sum[30]));
 BUF_X1 output91 (.A(net91),
    .Z(sum[31]));
 BUF_X1 output92 (.A(net92),
    .Z(sum[3]));
 BUF_X1 output93 (.A(net93),
    .Z(sum[4]));
 BUF_X1 output94 (.A(net94),
    .Z(sum[5]));
 BUF_X1 output95 (.A(net95),
    .Z(sum[6]));
 BUF_X1 output96 (.A(net96),
    .Z(sum[7]));
 BUF_X1 output97 (.A(net97),
    .Z(sum[8]));
 BUF_X1 output98 (.A(net98),
    .Z(sum[9]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X16 FILLER_0_792 ();
 FILLCELL_X4 FILLER_0_808 ();
 FILLCELL_X2 FILLER_0_812 ();
 FILLCELL_X1 FILLER_0_818 ();
 FILLCELL_X4 FILLER_0_825 ();
 FILLCELL_X8 FILLER_0_833 ();
 FILLCELL_X2 FILLER_0_841 ();
 FILLCELL_X2 FILLER_0_846 ();
 FILLCELL_X1 FILLER_0_848 ();
 FILLCELL_X16 FILLER_0_853 ();
 FILLCELL_X1 FILLER_0_869 ();
 FILLCELL_X16 FILLER_0_877 ();
 FILLCELL_X4 FILLER_0_901 ();
 FILLCELL_X1 FILLER_0_905 ();
 FILLCELL_X4 FILLER_0_909 ();
 FILLCELL_X2 FILLER_0_913 ();
 FILLCELL_X1 FILLER_0_915 ();
 FILLCELL_X32 FILLER_0_924 ();
 FILLCELL_X32 FILLER_0_956 ();
 FILLCELL_X32 FILLER_0_988 ();
 FILLCELL_X32 FILLER_0_1020 ();
 FILLCELL_X32 FILLER_0_1052 ();
 FILLCELL_X32 FILLER_0_1084 ();
 FILLCELL_X32 FILLER_0_1116 ();
 FILLCELL_X32 FILLER_0_1148 ();
 FILLCELL_X32 FILLER_0_1180 ();
 FILLCELL_X32 FILLER_0_1212 ();
 FILLCELL_X16 FILLER_0_1244 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X16 FILLER_0_1583 ();
 FILLCELL_X8 FILLER_0_1599 ();
 FILLCELL_X4 FILLER_0_1607 ();
 FILLCELL_X2 FILLER_0_1611 ();
 FILLCELL_X1 FILLER_0_1613 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X8 FILLER_1_801 ();
 FILLCELL_X4 FILLER_1_809 ();
 FILLCELL_X2 FILLER_1_813 ();
 FILLCELL_X1 FILLER_1_815 ();
 FILLCELL_X8 FILLER_1_820 ();
 FILLCELL_X2 FILLER_1_828 ();
 FILLCELL_X16 FILLER_1_834 ();
 FILLCELL_X2 FILLER_1_850 ();
 FILLCELL_X1 FILLER_1_852 ();
 FILLCELL_X16 FILLER_1_857 ();
 FILLCELL_X1 FILLER_1_873 ();
 FILLCELL_X32 FILLER_1_878 ();
 FILLCELL_X32 FILLER_1_910 ();
 FILLCELL_X32 FILLER_1_942 ();
 FILLCELL_X32 FILLER_1_974 ();
 FILLCELL_X32 FILLER_1_1006 ();
 FILLCELL_X32 FILLER_1_1038 ();
 FILLCELL_X32 FILLER_1_1070 ();
 FILLCELL_X32 FILLER_1_1102 ();
 FILLCELL_X32 FILLER_1_1134 ();
 FILLCELL_X32 FILLER_1_1166 ();
 FILLCELL_X32 FILLER_1_1198 ();
 FILLCELL_X32 FILLER_1_1230 ();
 FILLCELL_X1 FILLER_1_1262 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X16 FILLER_1_1584 ();
 FILLCELL_X8 FILLER_1_1600 ();
 FILLCELL_X4 FILLER_1_1608 ();
 FILLCELL_X2 FILLER_1_1612 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X16 FILLER_2_1592 ();
 FILLCELL_X4 FILLER_2_1608 ();
 FILLCELL_X2 FILLER_2_1612 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X16 FILLER_3_1584 ();
 FILLCELL_X8 FILLER_3_1600 ();
 FILLCELL_X4 FILLER_3_1608 ();
 FILLCELL_X2 FILLER_3_1612 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X16 FILLER_4_1592 ();
 FILLCELL_X4 FILLER_4_1608 ();
 FILLCELL_X2 FILLER_4_1612 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X16 FILLER_5_1584 ();
 FILLCELL_X8 FILLER_5_1600 ();
 FILLCELL_X4 FILLER_5_1608 ();
 FILLCELL_X2 FILLER_5_1612 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X16 FILLER_6_1592 ();
 FILLCELL_X4 FILLER_6_1608 ();
 FILLCELL_X2 FILLER_6_1612 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X16 FILLER_7_1584 ();
 FILLCELL_X8 FILLER_7_1600 ();
 FILLCELL_X4 FILLER_7_1608 ();
 FILLCELL_X2 FILLER_7_1612 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X16 FILLER_8_1592 ();
 FILLCELL_X4 FILLER_8_1608 ();
 FILLCELL_X2 FILLER_8_1612 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X16 FILLER_9_1584 ();
 FILLCELL_X8 FILLER_9_1600 ();
 FILLCELL_X4 FILLER_9_1608 ();
 FILLCELL_X2 FILLER_9_1612 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X16 FILLER_10_1592 ();
 FILLCELL_X4 FILLER_10_1608 ();
 FILLCELL_X2 FILLER_10_1612 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X16 FILLER_11_1584 ();
 FILLCELL_X8 FILLER_11_1600 ();
 FILLCELL_X4 FILLER_11_1608 ();
 FILLCELL_X2 FILLER_11_1612 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X16 FILLER_12_1592 ();
 FILLCELL_X4 FILLER_12_1608 ();
 FILLCELL_X2 FILLER_12_1612 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X16 FILLER_13_1584 ();
 FILLCELL_X8 FILLER_13_1600 ();
 FILLCELL_X4 FILLER_13_1608 ();
 FILLCELL_X2 FILLER_13_1612 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X16 FILLER_14_1592 ();
 FILLCELL_X4 FILLER_14_1608 ();
 FILLCELL_X2 FILLER_14_1612 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X16 FILLER_15_1584 ();
 FILLCELL_X8 FILLER_15_1600 ();
 FILLCELL_X4 FILLER_15_1608 ();
 FILLCELL_X2 FILLER_15_1612 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X16 FILLER_16_1592 ();
 FILLCELL_X4 FILLER_16_1608 ();
 FILLCELL_X2 FILLER_16_1612 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X16 FILLER_17_1584 ();
 FILLCELL_X8 FILLER_17_1600 ();
 FILLCELL_X4 FILLER_17_1608 ();
 FILLCELL_X2 FILLER_17_1612 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X16 FILLER_18_1592 ();
 FILLCELL_X4 FILLER_18_1608 ();
 FILLCELL_X2 FILLER_18_1612 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X16 FILLER_19_1584 ();
 FILLCELL_X8 FILLER_19_1600 ();
 FILLCELL_X4 FILLER_19_1608 ();
 FILLCELL_X2 FILLER_19_1612 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X16 FILLER_20_1592 ();
 FILLCELL_X4 FILLER_20_1608 ();
 FILLCELL_X2 FILLER_20_1612 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X16 FILLER_21_1584 ();
 FILLCELL_X8 FILLER_21_1600 ();
 FILLCELL_X4 FILLER_21_1608 ();
 FILLCELL_X2 FILLER_21_1612 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X16 FILLER_22_1592 ();
 FILLCELL_X4 FILLER_22_1608 ();
 FILLCELL_X2 FILLER_22_1612 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X16 FILLER_23_1584 ();
 FILLCELL_X8 FILLER_23_1600 ();
 FILLCELL_X4 FILLER_23_1608 ();
 FILLCELL_X2 FILLER_23_1612 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X16 FILLER_24_1592 ();
 FILLCELL_X4 FILLER_24_1608 ();
 FILLCELL_X2 FILLER_24_1612 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X16 FILLER_25_1584 ();
 FILLCELL_X8 FILLER_25_1600 ();
 FILLCELL_X4 FILLER_25_1608 ();
 FILLCELL_X2 FILLER_25_1612 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X16 FILLER_26_1592 ();
 FILLCELL_X4 FILLER_26_1608 ();
 FILLCELL_X2 FILLER_26_1612 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X16 FILLER_27_1584 ();
 FILLCELL_X8 FILLER_27_1600 ();
 FILLCELL_X4 FILLER_27_1608 ();
 FILLCELL_X2 FILLER_27_1612 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X16 FILLER_28_1592 ();
 FILLCELL_X4 FILLER_28_1608 ();
 FILLCELL_X2 FILLER_28_1612 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X16 FILLER_29_1584 ();
 FILLCELL_X8 FILLER_29_1600 ();
 FILLCELL_X4 FILLER_29_1608 ();
 FILLCELL_X2 FILLER_29_1612 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X16 FILLER_30_1592 ();
 FILLCELL_X4 FILLER_30_1608 ();
 FILLCELL_X2 FILLER_30_1612 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X16 FILLER_31_1584 ();
 FILLCELL_X8 FILLER_31_1600 ();
 FILLCELL_X4 FILLER_31_1608 ();
 FILLCELL_X2 FILLER_31_1612 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X16 FILLER_32_1592 ();
 FILLCELL_X4 FILLER_32_1608 ();
 FILLCELL_X2 FILLER_32_1612 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X16 FILLER_33_1584 ();
 FILLCELL_X8 FILLER_33_1600 ();
 FILLCELL_X4 FILLER_33_1608 ();
 FILLCELL_X2 FILLER_33_1612 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X16 FILLER_34_1592 ();
 FILLCELL_X4 FILLER_34_1608 ();
 FILLCELL_X2 FILLER_34_1612 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X16 FILLER_35_1584 ();
 FILLCELL_X8 FILLER_35_1600 ();
 FILLCELL_X4 FILLER_35_1608 ();
 FILLCELL_X2 FILLER_35_1612 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X16 FILLER_36_1592 ();
 FILLCELL_X4 FILLER_36_1608 ();
 FILLCELL_X2 FILLER_36_1612 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X16 FILLER_37_1584 ();
 FILLCELL_X8 FILLER_37_1600 ();
 FILLCELL_X4 FILLER_37_1608 ();
 FILLCELL_X2 FILLER_37_1612 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X16 FILLER_38_1592 ();
 FILLCELL_X4 FILLER_38_1608 ();
 FILLCELL_X2 FILLER_38_1612 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X16 FILLER_39_1584 ();
 FILLCELL_X8 FILLER_39_1600 ();
 FILLCELL_X4 FILLER_39_1608 ();
 FILLCELL_X2 FILLER_39_1612 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X16 FILLER_40_1592 ();
 FILLCELL_X4 FILLER_40_1608 ();
 FILLCELL_X2 FILLER_40_1612 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X16 FILLER_41_1584 ();
 FILLCELL_X8 FILLER_41_1600 ();
 FILLCELL_X4 FILLER_41_1608 ();
 FILLCELL_X2 FILLER_41_1612 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X16 FILLER_42_1592 ();
 FILLCELL_X4 FILLER_42_1608 ();
 FILLCELL_X2 FILLER_42_1612 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X16 FILLER_43_1584 ();
 FILLCELL_X8 FILLER_43_1600 ();
 FILLCELL_X4 FILLER_43_1608 ();
 FILLCELL_X2 FILLER_43_1612 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X16 FILLER_44_1592 ();
 FILLCELL_X4 FILLER_44_1608 ();
 FILLCELL_X2 FILLER_44_1612 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X16 FILLER_45_1584 ();
 FILLCELL_X8 FILLER_45_1600 ();
 FILLCELL_X4 FILLER_45_1608 ();
 FILLCELL_X2 FILLER_45_1612 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X16 FILLER_46_1592 ();
 FILLCELL_X4 FILLER_46_1608 ();
 FILLCELL_X2 FILLER_46_1612 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X16 FILLER_47_1584 ();
 FILLCELL_X8 FILLER_47_1600 ();
 FILLCELL_X4 FILLER_47_1608 ();
 FILLCELL_X2 FILLER_47_1612 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X16 FILLER_48_1592 ();
 FILLCELL_X4 FILLER_48_1608 ();
 FILLCELL_X2 FILLER_48_1612 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X16 FILLER_49_1584 ();
 FILLCELL_X8 FILLER_49_1600 ();
 FILLCELL_X4 FILLER_49_1608 ();
 FILLCELL_X2 FILLER_49_1612 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X16 FILLER_50_1592 ();
 FILLCELL_X4 FILLER_50_1608 ();
 FILLCELL_X2 FILLER_50_1612 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X16 FILLER_51_1584 ();
 FILLCELL_X8 FILLER_51_1600 ();
 FILLCELL_X4 FILLER_51_1608 ();
 FILLCELL_X2 FILLER_51_1612 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X16 FILLER_52_1592 ();
 FILLCELL_X4 FILLER_52_1608 ();
 FILLCELL_X2 FILLER_52_1612 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X16 FILLER_53_1584 ();
 FILLCELL_X8 FILLER_53_1600 ();
 FILLCELL_X4 FILLER_53_1608 ();
 FILLCELL_X2 FILLER_53_1612 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X16 FILLER_54_1592 ();
 FILLCELL_X4 FILLER_54_1608 ();
 FILLCELL_X2 FILLER_54_1612 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X16 FILLER_55_1584 ();
 FILLCELL_X8 FILLER_55_1600 ();
 FILLCELL_X4 FILLER_55_1608 ();
 FILLCELL_X2 FILLER_55_1612 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X16 FILLER_56_1592 ();
 FILLCELL_X4 FILLER_56_1608 ();
 FILLCELL_X2 FILLER_56_1612 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X16 FILLER_57_1584 ();
 FILLCELL_X8 FILLER_57_1600 ();
 FILLCELL_X4 FILLER_57_1608 ();
 FILLCELL_X2 FILLER_57_1612 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X16 FILLER_58_1592 ();
 FILLCELL_X4 FILLER_58_1608 ();
 FILLCELL_X2 FILLER_58_1612 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X16 FILLER_59_1584 ();
 FILLCELL_X8 FILLER_59_1600 ();
 FILLCELL_X4 FILLER_59_1608 ();
 FILLCELL_X2 FILLER_59_1612 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X16 FILLER_60_1592 ();
 FILLCELL_X4 FILLER_60_1608 ();
 FILLCELL_X2 FILLER_60_1612 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X16 FILLER_61_1584 ();
 FILLCELL_X8 FILLER_61_1600 ();
 FILLCELL_X4 FILLER_61_1608 ();
 FILLCELL_X2 FILLER_61_1612 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X16 FILLER_62_1592 ();
 FILLCELL_X4 FILLER_62_1608 ();
 FILLCELL_X2 FILLER_62_1612 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X16 FILLER_63_1584 ();
 FILLCELL_X8 FILLER_63_1600 ();
 FILLCELL_X4 FILLER_63_1608 ();
 FILLCELL_X2 FILLER_63_1612 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X16 FILLER_64_1592 ();
 FILLCELL_X4 FILLER_64_1608 ();
 FILLCELL_X2 FILLER_64_1612 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X16 FILLER_65_1584 ();
 FILLCELL_X8 FILLER_65_1600 ();
 FILLCELL_X4 FILLER_65_1608 ();
 FILLCELL_X2 FILLER_65_1612 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X16 FILLER_66_1592 ();
 FILLCELL_X4 FILLER_66_1608 ();
 FILLCELL_X2 FILLER_66_1612 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X16 FILLER_67_1584 ();
 FILLCELL_X8 FILLER_67_1600 ();
 FILLCELL_X4 FILLER_67_1608 ();
 FILLCELL_X2 FILLER_67_1612 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X16 FILLER_68_1592 ();
 FILLCELL_X4 FILLER_68_1608 ();
 FILLCELL_X2 FILLER_68_1612 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X16 FILLER_69_1584 ();
 FILLCELL_X8 FILLER_69_1600 ();
 FILLCELL_X4 FILLER_69_1608 ();
 FILLCELL_X2 FILLER_69_1612 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X16 FILLER_70_1592 ();
 FILLCELL_X4 FILLER_70_1608 ();
 FILLCELL_X2 FILLER_70_1612 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X16 FILLER_71_1584 ();
 FILLCELL_X8 FILLER_71_1600 ();
 FILLCELL_X4 FILLER_71_1608 ();
 FILLCELL_X2 FILLER_71_1612 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X16 FILLER_72_1592 ();
 FILLCELL_X4 FILLER_72_1608 ();
 FILLCELL_X2 FILLER_72_1612 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X16 FILLER_73_1584 ();
 FILLCELL_X8 FILLER_73_1600 ();
 FILLCELL_X4 FILLER_73_1608 ();
 FILLCELL_X2 FILLER_73_1612 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X16 FILLER_74_1592 ();
 FILLCELL_X4 FILLER_74_1608 ();
 FILLCELL_X2 FILLER_74_1612 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X16 FILLER_75_1584 ();
 FILLCELL_X8 FILLER_75_1600 ();
 FILLCELL_X4 FILLER_75_1608 ();
 FILLCELL_X2 FILLER_75_1612 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X16 FILLER_76_1592 ();
 FILLCELL_X4 FILLER_76_1608 ();
 FILLCELL_X2 FILLER_76_1612 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X16 FILLER_77_1584 ();
 FILLCELL_X8 FILLER_77_1600 ();
 FILLCELL_X4 FILLER_77_1608 ();
 FILLCELL_X2 FILLER_77_1612 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X16 FILLER_78_1592 ();
 FILLCELL_X4 FILLER_78_1608 ();
 FILLCELL_X2 FILLER_78_1612 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X16 FILLER_79_1584 ();
 FILLCELL_X8 FILLER_79_1600 ();
 FILLCELL_X4 FILLER_79_1608 ();
 FILLCELL_X2 FILLER_79_1612 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X16 FILLER_80_1592 ();
 FILLCELL_X4 FILLER_80_1608 ();
 FILLCELL_X2 FILLER_80_1612 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X16 FILLER_81_1584 ();
 FILLCELL_X8 FILLER_81_1600 ();
 FILLCELL_X4 FILLER_81_1608 ();
 FILLCELL_X2 FILLER_81_1612 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X16 FILLER_82_1592 ();
 FILLCELL_X4 FILLER_82_1608 ();
 FILLCELL_X2 FILLER_82_1612 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X16 FILLER_83_1584 ();
 FILLCELL_X8 FILLER_83_1600 ();
 FILLCELL_X4 FILLER_83_1608 ();
 FILLCELL_X2 FILLER_83_1612 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X16 FILLER_84_1592 ();
 FILLCELL_X4 FILLER_84_1608 ();
 FILLCELL_X2 FILLER_84_1612 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X16 FILLER_85_1584 ();
 FILLCELL_X8 FILLER_85_1600 ();
 FILLCELL_X4 FILLER_85_1608 ();
 FILLCELL_X2 FILLER_85_1612 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X16 FILLER_86_1592 ();
 FILLCELL_X4 FILLER_86_1608 ();
 FILLCELL_X2 FILLER_86_1612 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X16 FILLER_87_1584 ();
 FILLCELL_X8 FILLER_87_1600 ();
 FILLCELL_X4 FILLER_87_1608 ();
 FILLCELL_X2 FILLER_87_1612 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X16 FILLER_88_1592 ();
 FILLCELL_X4 FILLER_88_1608 ();
 FILLCELL_X2 FILLER_88_1612 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X16 FILLER_89_1584 ();
 FILLCELL_X8 FILLER_89_1600 ();
 FILLCELL_X4 FILLER_89_1608 ();
 FILLCELL_X2 FILLER_89_1612 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X16 FILLER_90_1592 ();
 FILLCELL_X4 FILLER_90_1608 ();
 FILLCELL_X2 FILLER_90_1612 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X16 FILLER_91_1584 ();
 FILLCELL_X8 FILLER_91_1600 ();
 FILLCELL_X4 FILLER_91_1608 ();
 FILLCELL_X2 FILLER_91_1612 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X16 FILLER_92_1592 ();
 FILLCELL_X4 FILLER_92_1608 ();
 FILLCELL_X2 FILLER_92_1612 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X16 FILLER_93_1584 ();
 FILLCELL_X8 FILLER_93_1600 ();
 FILLCELL_X4 FILLER_93_1608 ();
 FILLCELL_X2 FILLER_93_1612 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X16 FILLER_94_1592 ();
 FILLCELL_X4 FILLER_94_1608 ();
 FILLCELL_X2 FILLER_94_1612 ();
 FILLCELL_X1 FILLER_95_7 ();
 FILLCELL_X32 FILLER_95_18 ();
 FILLCELL_X32 FILLER_95_50 ();
 FILLCELL_X32 FILLER_95_82 ();
 FILLCELL_X32 FILLER_95_114 ();
 FILLCELL_X32 FILLER_95_146 ();
 FILLCELL_X32 FILLER_95_178 ();
 FILLCELL_X32 FILLER_95_210 ();
 FILLCELL_X32 FILLER_95_242 ();
 FILLCELL_X32 FILLER_95_274 ();
 FILLCELL_X32 FILLER_95_306 ();
 FILLCELL_X32 FILLER_95_338 ();
 FILLCELL_X32 FILLER_95_370 ();
 FILLCELL_X32 FILLER_95_402 ();
 FILLCELL_X32 FILLER_95_434 ();
 FILLCELL_X32 FILLER_95_466 ();
 FILLCELL_X32 FILLER_95_498 ();
 FILLCELL_X32 FILLER_95_530 ();
 FILLCELL_X32 FILLER_95_562 ();
 FILLCELL_X32 FILLER_95_594 ();
 FILLCELL_X32 FILLER_95_626 ();
 FILLCELL_X32 FILLER_95_658 ();
 FILLCELL_X32 FILLER_95_690 ();
 FILLCELL_X32 FILLER_95_722 ();
 FILLCELL_X32 FILLER_95_754 ();
 FILLCELL_X32 FILLER_95_786 ();
 FILLCELL_X32 FILLER_95_818 ();
 FILLCELL_X32 FILLER_95_850 ();
 FILLCELL_X32 FILLER_95_882 ();
 FILLCELL_X32 FILLER_95_914 ();
 FILLCELL_X32 FILLER_95_946 ();
 FILLCELL_X32 FILLER_95_978 ();
 FILLCELL_X32 FILLER_95_1010 ();
 FILLCELL_X32 FILLER_95_1042 ();
 FILLCELL_X32 FILLER_95_1074 ();
 FILLCELL_X32 FILLER_95_1106 ();
 FILLCELL_X32 FILLER_95_1138 ();
 FILLCELL_X32 FILLER_95_1170 ();
 FILLCELL_X32 FILLER_95_1202 ();
 FILLCELL_X16 FILLER_95_1234 ();
 FILLCELL_X8 FILLER_95_1250 ();
 FILLCELL_X4 FILLER_95_1258 ();
 FILLCELL_X1 FILLER_95_1262 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X16 FILLER_95_1584 ();
 FILLCELL_X8 FILLER_95_1600 ();
 FILLCELL_X4 FILLER_95_1608 ();
 FILLCELL_X2 FILLER_95_1612 ();
 FILLCELL_X4 FILLER_96_4 ();
 FILLCELL_X1 FILLER_96_8 ();
 FILLCELL_X8 FILLER_96_14 ();
 FILLCELL_X1 FILLER_96_22 ();
 FILLCELL_X8 FILLER_96_31 ();
 FILLCELL_X1 FILLER_96_39 ();
 FILLCELL_X32 FILLER_96_43 ();
 FILLCELL_X32 FILLER_96_75 ();
 FILLCELL_X32 FILLER_96_107 ();
 FILLCELL_X32 FILLER_96_139 ();
 FILLCELL_X32 FILLER_96_171 ();
 FILLCELL_X32 FILLER_96_203 ();
 FILLCELL_X32 FILLER_96_235 ();
 FILLCELL_X32 FILLER_96_267 ();
 FILLCELL_X32 FILLER_96_299 ();
 FILLCELL_X32 FILLER_96_331 ();
 FILLCELL_X32 FILLER_96_363 ();
 FILLCELL_X32 FILLER_96_395 ();
 FILLCELL_X32 FILLER_96_427 ();
 FILLCELL_X32 FILLER_96_459 ();
 FILLCELL_X32 FILLER_96_491 ();
 FILLCELL_X32 FILLER_96_523 ();
 FILLCELL_X32 FILLER_96_555 ();
 FILLCELL_X32 FILLER_96_587 ();
 FILLCELL_X8 FILLER_96_619 ();
 FILLCELL_X4 FILLER_96_627 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X16 FILLER_96_1592 ();
 FILLCELL_X4 FILLER_96_1608 ();
 FILLCELL_X2 FILLER_96_1612 ();
 FILLCELL_X1 FILLER_97_1 ();
 FILLCELL_X4 FILLER_97_8 ();
 FILLCELL_X2 FILLER_97_12 ();
 FILLCELL_X1 FILLER_97_17 ();
 FILLCELL_X1 FILLER_97_21 ();
 FILLCELL_X1 FILLER_97_32 ();
 FILLCELL_X2 FILLER_97_37 ();
 FILLCELL_X4 FILLER_97_43 ();
 FILLCELL_X2 FILLER_97_47 ();
 FILLCELL_X32 FILLER_97_54 ();
 FILLCELL_X32 FILLER_97_86 ();
 FILLCELL_X32 FILLER_97_118 ();
 FILLCELL_X32 FILLER_97_150 ();
 FILLCELL_X32 FILLER_97_182 ();
 FILLCELL_X32 FILLER_97_214 ();
 FILLCELL_X32 FILLER_97_246 ();
 FILLCELL_X32 FILLER_97_278 ();
 FILLCELL_X32 FILLER_97_310 ();
 FILLCELL_X32 FILLER_97_342 ();
 FILLCELL_X32 FILLER_97_374 ();
 FILLCELL_X32 FILLER_97_406 ();
 FILLCELL_X32 FILLER_97_438 ();
 FILLCELL_X32 FILLER_97_470 ();
 FILLCELL_X32 FILLER_97_502 ();
 FILLCELL_X32 FILLER_97_534 ();
 FILLCELL_X32 FILLER_97_566 ();
 FILLCELL_X32 FILLER_97_598 ();
 FILLCELL_X32 FILLER_97_630 ();
 FILLCELL_X32 FILLER_97_662 ();
 FILLCELL_X32 FILLER_97_694 ();
 FILLCELL_X32 FILLER_97_726 ();
 FILLCELL_X32 FILLER_97_758 ();
 FILLCELL_X32 FILLER_97_790 ();
 FILLCELL_X32 FILLER_97_822 ();
 FILLCELL_X16 FILLER_97_854 ();
 FILLCELL_X2 FILLER_97_870 ();
 FILLCELL_X1 FILLER_97_872 ();
 FILLCELL_X8 FILLER_97_883 ();
 FILLCELL_X2 FILLER_97_891 ();
 FILLCELL_X8 FILLER_97_903 ();
 FILLCELL_X4 FILLER_97_911 ();
 FILLCELL_X1 FILLER_97_915 ();
 FILLCELL_X32 FILLER_97_926 ();
 FILLCELL_X32 FILLER_97_958 ();
 FILLCELL_X32 FILLER_97_990 ();
 FILLCELL_X32 FILLER_97_1022 ();
 FILLCELL_X32 FILLER_97_1054 ();
 FILLCELL_X32 FILLER_97_1086 ();
 FILLCELL_X32 FILLER_97_1118 ();
 FILLCELL_X32 FILLER_97_1150 ();
 FILLCELL_X32 FILLER_97_1182 ();
 FILLCELL_X32 FILLER_97_1214 ();
 FILLCELL_X16 FILLER_97_1246 ();
 FILLCELL_X1 FILLER_97_1262 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X16 FILLER_97_1584 ();
 FILLCELL_X8 FILLER_97_1600 ();
 FILLCELL_X4 FILLER_97_1608 ();
 FILLCELL_X2 FILLER_97_1612 ();
 FILLCELL_X2 FILLER_98_4 ();
 FILLCELL_X16 FILLER_98_20 ();
 FILLCELL_X8 FILLER_98_36 ();
 FILLCELL_X4 FILLER_98_51 ();
 FILLCELL_X1 FILLER_98_55 ();
 FILLCELL_X32 FILLER_98_59 ();
 FILLCELL_X32 FILLER_98_91 ();
 FILLCELL_X32 FILLER_98_123 ();
 FILLCELL_X32 FILLER_98_155 ();
 FILLCELL_X32 FILLER_98_187 ();
 FILLCELL_X32 FILLER_98_219 ();
 FILLCELL_X32 FILLER_98_251 ();
 FILLCELL_X32 FILLER_98_283 ();
 FILLCELL_X32 FILLER_98_315 ();
 FILLCELL_X32 FILLER_98_347 ();
 FILLCELL_X32 FILLER_98_379 ();
 FILLCELL_X32 FILLER_98_411 ();
 FILLCELL_X32 FILLER_98_443 ();
 FILLCELL_X32 FILLER_98_475 ();
 FILLCELL_X32 FILLER_98_507 ();
 FILLCELL_X32 FILLER_98_539 ();
 FILLCELL_X32 FILLER_98_571 ();
 FILLCELL_X16 FILLER_98_603 ();
 FILLCELL_X8 FILLER_98_619 ();
 FILLCELL_X4 FILLER_98_627 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X4 FILLER_98_824 ();
 FILLCELL_X2 FILLER_98_828 ();
 FILLCELL_X8 FILLER_98_840 ();
 FILLCELL_X2 FILLER_98_848 ();
 FILLCELL_X1 FILLER_98_850 ();
 FILLCELL_X32 FILLER_98_861 ();
 FILLCELL_X32 FILLER_98_898 ();
 FILLCELL_X32 FILLER_98_930 ();
 FILLCELL_X32 FILLER_98_962 ();
 FILLCELL_X32 FILLER_98_994 ();
 FILLCELL_X32 FILLER_98_1026 ();
 FILLCELL_X32 FILLER_98_1058 ();
 FILLCELL_X32 FILLER_98_1090 ();
 FILLCELL_X32 FILLER_98_1122 ();
 FILLCELL_X32 FILLER_98_1154 ();
 FILLCELL_X32 FILLER_98_1186 ();
 FILLCELL_X32 FILLER_98_1218 ();
 FILLCELL_X32 FILLER_98_1250 ();
 FILLCELL_X32 FILLER_98_1282 ();
 FILLCELL_X32 FILLER_98_1314 ();
 FILLCELL_X32 FILLER_98_1346 ();
 FILLCELL_X32 FILLER_98_1378 ();
 FILLCELL_X32 FILLER_98_1410 ();
 FILLCELL_X32 FILLER_98_1442 ();
 FILLCELL_X32 FILLER_98_1474 ();
 FILLCELL_X32 FILLER_98_1506 ();
 FILLCELL_X32 FILLER_98_1538 ();
 FILLCELL_X32 FILLER_98_1570 ();
 FILLCELL_X8 FILLER_98_1602 ();
 FILLCELL_X4 FILLER_98_1610 ();
 FILLCELL_X2 FILLER_99_1 ();
 FILLCELL_X1 FILLER_99_3 ();
 FILLCELL_X4 FILLER_99_7 ();
 FILLCELL_X2 FILLER_99_14 ();
 FILLCELL_X1 FILLER_99_16 ();
 FILLCELL_X8 FILLER_99_20 ();
 FILLCELL_X4 FILLER_99_28 ();
 FILLCELL_X1 FILLER_99_32 ();
 FILLCELL_X8 FILLER_99_37 ();
 FILLCELL_X2 FILLER_99_45 ();
 FILLCELL_X1 FILLER_99_47 ();
 FILLCELL_X4 FILLER_99_52 ();
 FILLCELL_X32 FILLER_99_63 ();
 FILLCELL_X32 FILLER_99_95 ();
 FILLCELL_X32 FILLER_99_127 ();
 FILLCELL_X32 FILLER_99_159 ();
 FILLCELL_X32 FILLER_99_191 ();
 FILLCELL_X32 FILLER_99_223 ();
 FILLCELL_X32 FILLER_99_255 ();
 FILLCELL_X32 FILLER_99_287 ();
 FILLCELL_X32 FILLER_99_319 ();
 FILLCELL_X32 FILLER_99_351 ();
 FILLCELL_X32 FILLER_99_383 ();
 FILLCELL_X32 FILLER_99_415 ();
 FILLCELL_X32 FILLER_99_447 ();
 FILLCELL_X32 FILLER_99_479 ();
 FILLCELL_X32 FILLER_99_511 ();
 FILLCELL_X32 FILLER_99_543 ();
 FILLCELL_X32 FILLER_99_575 ();
 FILLCELL_X32 FILLER_99_607 ();
 FILLCELL_X32 FILLER_99_639 ();
 FILLCELL_X32 FILLER_99_671 ();
 FILLCELL_X32 FILLER_99_703 ();
 FILLCELL_X32 FILLER_99_735 ();
 FILLCELL_X32 FILLER_99_767 ();
 FILLCELL_X16 FILLER_99_799 ();
 FILLCELL_X1 FILLER_99_815 ();
 FILLCELL_X16 FILLER_99_826 ();
 FILLCELL_X8 FILLER_99_842 ();
 FILLCELL_X1 FILLER_99_850 ();
 FILLCELL_X16 FILLER_99_858 ();
 FILLCELL_X32 FILLER_99_879 ();
 FILLCELL_X4 FILLER_99_911 ();
 FILLCELL_X2 FILLER_99_915 ();
 FILLCELL_X32 FILLER_99_921 ();
 FILLCELL_X32 FILLER_99_953 ();
 FILLCELL_X32 FILLER_99_985 ();
 FILLCELL_X32 FILLER_99_1017 ();
 FILLCELL_X32 FILLER_99_1049 ();
 FILLCELL_X32 FILLER_99_1081 ();
 FILLCELL_X32 FILLER_99_1113 ();
 FILLCELL_X32 FILLER_99_1145 ();
 FILLCELL_X32 FILLER_99_1177 ();
 FILLCELL_X32 FILLER_99_1209 ();
 FILLCELL_X16 FILLER_99_1241 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X16 FILLER_99_1584 ();
 FILLCELL_X8 FILLER_99_1600 ();
 FILLCELL_X4 FILLER_99_1608 ();
 FILLCELL_X2 FILLER_99_1612 ();
 FILLCELL_X4 FILLER_100_1 ();
 FILLCELL_X2 FILLER_100_5 ();
 FILLCELL_X1 FILLER_100_7 ();
 FILLCELL_X1 FILLER_100_10 ();
 FILLCELL_X4 FILLER_100_20 ();
 FILLCELL_X8 FILLER_100_39 ();
 FILLCELL_X4 FILLER_100_47 ();
 FILLCELL_X2 FILLER_100_51 ();
 FILLCELL_X1 FILLER_100_53 ();
 FILLCELL_X2 FILLER_100_61 ();
 FILLCELL_X1 FILLER_100_75 ();
 FILLCELL_X32 FILLER_100_78 ();
 FILLCELL_X32 FILLER_100_110 ();
 FILLCELL_X32 FILLER_100_142 ();
 FILLCELL_X32 FILLER_100_174 ();
 FILLCELL_X32 FILLER_100_206 ();
 FILLCELL_X32 FILLER_100_238 ();
 FILLCELL_X32 FILLER_100_270 ();
 FILLCELL_X32 FILLER_100_302 ();
 FILLCELL_X32 FILLER_100_334 ();
 FILLCELL_X32 FILLER_100_366 ();
 FILLCELL_X32 FILLER_100_398 ();
 FILLCELL_X32 FILLER_100_430 ();
 FILLCELL_X32 FILLER_100_462 ();
 FILLCELL_X32 FILLER_100_494 ();
 FILLCELL_X32 FILLER_100_526 ();
 FILLCELL_X32 FILLER_100_558 ();
 FILLCELL_X32 FILLER_100_590 ();
 FILLCELL_X8 FILLER_100_622 ();
 FILLCELL_X1 FILLER_100_630 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X16 FILLER_100_792 ();
 FILLCELL_X8 FILLER_100_808 ();
 FILLCELL_X1 FILLER_100_816 ();
 FILLCELL_X8 FILLER_100_822 ();
 FILLCELL_X1 FILLER_100_830 ();
 FILLCELL_X16 FILLER_100_838 ();
 FILLCELL_X8 FILLER_100_854 ();
 FILLCELL_X4 FILLER_100_862 ();
 FILLCELL_X32 FILLER_100_875 ();
 FILLCELL_X4 FILLER_100_907 ();
 FILLCELL_X1 FILLER_100_911 ();
 FILLCELL_X8 FILLER_100_914 ();
 FILLCELL_X32 FILLER_100_926 ();
 FILLCELL_X32 FILLER_100_958 ();
 FILLCELL_X32 FILLER_100_990 ();
 FILLCELL_X32 FILLER_100_1022 ();
 FILLCELL_X32 FILLER_100_1054 ();
 FILLCELL_X32 FILLER_100_1086 ();
 FILLCELL_X32 FILLER_100_1118 ();
 FILLCELL_X32 FILLER_100_1150 ();
 FILLCELL_X32 FILLER_100_1182 ();
 FILLCELL_X32 FILLER_100_1214 ();
 FILLCELL_X32 FILLER_100_1246 ();
 FILLCELL_X32 FILLER_100_1278 ();
 FILLCELL_X32 FILLER_100_1310 ();
 FILLCELL_X32 FILLER_100_1342 ();
 FILLCELL_X32 FILLER_100_1374 ();
 FILLCELL_X32 FILLER_100_1406 ();
 FILLCELL_X32 FILLER_100_1438 ();
 FILLCELL_X32 FILLER_100_1470 ();
 FILLCELL_X32 FILLER_100_1502 ();
 FILLCELL_X32 FILLER_100_1534 ();
 FILLCELL_X32 FILLER_100_1566 ();
 FILLCELL_X16 FILLER_100_1598 ();
 FILLCELL_X1 FILLER_101_1 ();
 FILLCELL_X2 FILLER_101_22 ();
 FILLCELL_X1 FILLER_101_24 ();
 FILLCELL_X1 FILLER_101_45 ();
 FILLCELL_X2 FILLER_101_53 ();
 FILLCELL_X2 FILLER_101_59 ();
 FILLCELL_X32 FILLER_101_78 ();
 FILLCELL_X32 FILLER_101_110 ();
 FILLCELL_X32 FILLER_101_142 ();
 FILLCELL_X32 FILLER_101_174 ();
 FILLCELL_X32 FILLER_101_206 ();
 FILLCELL_X32 FILLER_101_238 ();
 FILLCELL_X32 FILLER_101_270 ();
 FILLCELL_X32 FILLER_101_302 ();
 FILLCELL_X32 FILLER_101_334 ();
 FILLCELL_X32 FILLER_101_366 ();
 FILLCELL_X32 FILLER_101_398 ();
 FILLCELL_X32 FILLER_101_430 ();
 FILLCELL_X32 FILLER_101_462 ();
 FILLCELL_X32 FILLER_101_494 ();
 FILLCELL_X32 FILLER_101_526 ();
 FILLCELL_X32 FILLER_101_558 ();
 FILLCELL_X32 FILLER_101_590 ();
 FILLCELL_X32 FILLER_101_622 ();
 FILLCELL_X32 FILLER_101_654 ();
 FILLCELL_X32 FILLER_101_686 ();
 FILLCELL_X32 FILLER_101_718 ();
 FILLCELL_X8 FILLER_101_750 ();
 FILLCELL_X4 FILLER_101_758 ();
 FILLCELL_X2 FILLER_101_762 ();
 FILLCELL_X1 FILLER_101_764 ();
 FILLCELL_X32 FILLER_101_775 ();
 FILLCELL_X32 FILLER_101_807 ();
 FILLCELL_X4 FILLER_101_839 ();
 FILLCELL_X1 FILLER_101_843 ();
 FILLCELL_X4 FILLER_101_853 ();
 FILLCELL_X2 FILLER_101_857 ();
 FILLCELL_X1 FILLER_101_859 ();
 FILLCELL_X8 FILLER_101_867 ();
 FILLCELL_X4 FILLER_101_875 ();
 FILLCELL_X8 FILLER_101_883 ();
 FILLCELL_X4 FILLER_101_898 ();
 FILLCELL_X32 FILLER_101_922 ();
 FILLCELL_X32 FILLER_101_954 ();
 FILLCELL_X32 FILLER_101_986 ();
 FILLCELL_X32 FILLER_101_1018 ();
 FILLCELL_X32 FILLER_101_1050 ();
 FILLCELL_X32 FILLER_101_1082 ();
 FILLCELL_X32 FILLER_101_1114 ();
 FILLCELL_X32 FILLER_101_1146 ();
 FILLCELL_X32 FILLER_101_1178 ();
 FILLCELL_X32 FILLER_101_1210 ();
 FILLCELL_X16 FILLER_101_1242 ();
 FILLCELL_X4 FILLER_101_1258 ();
 FILLCELL_X1 FILLER_101_1262 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X16 FILLER_101_1584 ();
 FILLCELL_X8 FILLER_101_1600 ();
 FILLCELL_X4 FILLER_101_1608 ();
 FILLCELL_X2 FILLER_101_1612 ();
 FILLCELL_X1 FILLER_102_4 ();
 FILLCELL_X4 FILLER_102_12 ();
 FILLCELL_X2 FILLER_102_16 ();
 FILLCELL_X1 FILLER_102_18 ();
 FILLCELL_X4 FILLER_102_29 ();
 FILLCELL_X8 FILLER_102_35 ();
 FILLCELL_X2 FILLER_102_47 ();
 FILLCELL_X1 FILLER_102_49 ();
 FILLCELL_X4 FILLER_102_55 ();
 FILLCELL_X1 FILLER_102_59 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X8 FILLER_102_792 ();
 FILLCELL_X8 FILLER_102_805 ();
 FILLCELL_X2 FILLER_102_813 ();
 FILLCELL_X1 FILLER_102_815 ();
 FILLCELL_X2 FILLER_102_845 ();
 FILLCELL_X1 FILLER_102_847 ();
 FILLCELL_X16 FILLER_102_853 ();
 FILLCELL_X2 FILLER_102_869 ();
 FILLCELL_X16 FILLER_102_876 ();
 FILLCELL_X8 FILLER_102_892 ();
 FILLCELL_X4 FILLER_102_900 ();
 FILLCELL_X1 FILLER_102_904 ();
 FILLCELL_X32 FILLER_102_907 ();
 FILLCELL_X32 FILLER_102_939 ();
 FILLCELL_X32 FILLER_102_971 ();
 FILLCELL_X32 FILLER_102_1003 ();
 FILLCELL_X32 FILLER_102_1035 ();
 FILLCELL_X32 FILLER_102_1067 ();
 FILLCELL_X32 FILLER_102_1099 ();
 FILLCELL_X32 FILLER_102_1131 ();
 FILLCELL_X32 FILLER_102_1163 ();
 FILLCELL_X32 FILLER_102_1195 ();
 FILLCELL_X32 FILLER_102_1227 ();
 FILLCELL_X32 FILLER_102_1259 ();
 FILLCELL_X32 FILLER_102_1291 ();
 FILLCELL_X32 FILLER_102_1323 ();
 FILLCELL_X32 FILLER_102_1355 ();
 FILLCELL_X32 FILLER_102_1387 ();
 FILLCELL_X32 FILLER_102_1419 ();
 FILLCELL_X32 FILLER_102_1451 ();
 FILLCELL_X32 FILLER_102_1483 ();
 FILLCELL_X32 FILLER_102_1515 ();
 FILLCELL_X32 FILLER_102_1547 ();
 FILLCELL_X32 FILLER_102_1579 ();
 FILLCELL_X2 FILLER_102_1611 ();
 FILLCELL_X1 FILLER_102_1613 ();
 FILLCELL_X1 FILLER_103_1 ();
 FILLCELL_X2 FILLER_103_5 ();
 FILLCELL_X16 FILLER_103_10 ();
 FILLCELL_X8 FILLER_103_26 ();
 FILLCELL_X2 FILLER_103_34 ();
 FILLCELL_X1 FILLER_103_36 ();
 FILLCELL_X4 FILLER_103_41 ();
 FILLCELL_X2 FILLER_103_45 ();
 FILLCELL_X1 FILLER_103_47 ();
 FILLCELL_X2 FILLER_103_53 ();
 FILLCELL_X1 FILLER_103_55 ();
 FILLCELL_X32 FILLER_103_69 ();
 FILLCELL_X32 FILLER_103_101 ();
 FILLCELL_X32 FILLER_103_133 ();
 FILLCELL_X32 FILLER_103_165 ();
 FILLCELL_X32 FILLER_103_197 ();
 FILLCELL_X32 FILLER_103_229 ();
 FILLCELL_X32 FILLER_103_261 ();
 FILLCELL_X32 FILLER_103_293 ();
 FILLCELL_X32 FILLER_103_325 ();
 FILLCELL_X32 FILLER_103_357 ();
 FILLCELL_X32 FILLER_103_389 ();
 FILLCELL_X32 FILLER_103_421 ();
 FILLCELL_X32 FILLER_103_453 ();
 FILLCELL_X32 FILLER_103_485 ();
 FILLCELL_X32 FILLER_103_517 ();
 FILLCELL_X32 FILLER_103_549 ();
 FILLCELL_X32 FILLER_103_581 ();
 FILLCELL_X32 FILLER_103_613 ();
 FILLCELL_X32 FILLER_103_645 ();
 FILLCELL_X32 FILLER_103_677 ();
 FILLCELL_X32 FILLER_103_709 ();
 FILLCELL_X32 FILLER_103_741 ();
 FILLCELL_X32 FILLER_103_773 ();
 FILLCELL_X16 FILLER_103_805 ();
 FILLCELL_X2 FILLER_103_821 ();
 FILLCELL_X1 FILLER_103_823 ();
 FILLCELL_X2 FILLER_103_834 ();
 FILLCELL_X2 FILLER_103_841 ();
 FILLCELL_X1 FILLER_103_843 ();
 FILLCELL_X4 FILLER_103_862 ();
 FILLCELL_X1 FILLER_103_876 ();
 FILLCELL_X2 FILLER_103_881 ();
 FILLCELL_X1 FILLER_103_903 ();
 FILLCELL_X32 FILLER_103_908 ();
 FILLCELL_X32 FILLER_103_940 ();
 FILLCELL_X32 FILLER_103_972 ();
 FILLCELL_X32 FILLER_103_1004 ();
 FILLCELL_X32 FILLER_103_1036 ();
 FILLCELL_X32 FILLER_103_1068 ();
 FILLCELL_X32 FILLER_103_1100 ();
 FILLCELL_X32 FILLER_103_1132 ();
 FILLCELL_X32 FILLER_103_1164 ();
 FILLCELL_X32 FILLER_103_1196 ();
 FILLCELL_X32 FILLER_103_1228 ();
 FILLCELL_X2 FILLER_103_1260 ();
 FILLCELL_X1 FILLER_103_1262 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X16 FILLER_103_1584 ();
 FILLCELL_X8 FILLER_103_1600 ();
 FILLCELL_X4 FILLER_103_1608 ();
 FILLCELL_X2 FILLER_103_1612 ();
 FILLCELL_X4 FILLER_104_1 ();
 FILLCELL_X1 FILLER_104_5 ();
 FILLCELL_X2 FILLER_104_16 ();
 FILLCELL_X1 FILLER_104_18 ();
 FILLCELL_X1 FILLER_104_27 ();
 FILLCELL_X8 FILLER_104_32 ();
 FILLCELL_X1 FILLER_104_40 ();
 FILLCELL_X32 FILLER_104_52 ();
 FILLCELL_X32 FILLER_104_84 ();
 FILLCELL_X32 FILLER_104_116 ();
 FILLCELL_X32 FILLER_104_148 ();
 FILLCELL_X32 FILLER_104_180 ();
 FILLCELL_X32 FILLER_104_212 ();
 FILLCELL_X32 FILLER_104_244 ();
 FILLCELL_X32 FILLER_104_276 ();
 FILLCELL_X32 FILLER_104_308 ();
 FILLCELL_X32 FILLER_104_340 ();
 FILLCELL_X32 FILLER_104_372 ();
 FILLCELL_X32 FILLER_104_404 ();
 FILLCELL_X32 FILLER_104_436 ();
 FILLCELL_X32 FILLER_104_468 ();
 FILLCELL_X32 FILLER_104_500 ();
 FILLCELL_X32 FILLER_104_532 ();
 FILLCELL_X32 FILLER_104_564 ();
 FILLCELL_X32 FILLER_104_596 ();
 FILLCELL_X2 FILLER_104_628 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X16 FILLER_104_728 ();
 FILLCELL_X8 FILLER_104_744 ();
 FILLCELL_X4 FILLER_104_752 ();
 FILLCELL_X2 FILLER_104_756 ();
 FILLCELL_X1 FILLER_104_758 ();
 FILLCELL_X32 FILLER_104_769 ();
 FILLCELL_X16 FILLER_104_801 ();
 FILLCELL_X8 FILLER_104_817 ();
 FILLCELL_X2 FILLER_104_825 ();
 FILLCELL_X16 FILLER_104_841 ();
 FILLCELL_X8 FILLER_104_857 ();
 FILLCELL_X4 FILLER_104_865 ();
 FILLCELL_X1 FILLER_104_869 ();
 FILLCELL_X4 FILLER_104_873 ();
 FILLCELL_X8 FILLER_104_883 ();
 FILLCELL_X4 FILLER_104_891 ();
 FILLCELL_X2 FILLER_104_895 ();
 FILLCELL_X1 FILLER_104_897 ();
 FILLCELL_X2 FILLER_104_901 ();
 FILLCELL_X4 FILLER_104_905 ();
 FILLCELL_X1 FILLER_104_909 ();
 FILLCELL_X1 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_925 ();
 FILLCELL_X32 FILLER_104_957 ();
 FILLCELL_X32 FILLER_104_989 ();
 FILLCELL_X32 FILLER_104_1021 ();
 FILLCELL_X32 FILLER_104_1053 ();
 FILLCELL_X32 FILLER_104_1085 ();
 FILLCELL_X32 FILLER_104_1117 ();
 FILLCELL_X32 FILLER_104_1149 ();
 FILLCELL_X32 FILLER_104_1181 ();
 FILLCELL_X32 FILLER_104_1213 ();
 FILLCELL_X32 FILLER_104_1245 ();
 FILLCELL_X32 FILLER_104_1277 ();
 FILLCELL_X32 FILLER_104_1309 ();
 FILLCELL_X32 FILLER_104_1341 ();
 FILLCELL_X32 FILLER_104_1373 ();
 FILLCELL_X32 FILLER_104_1405 ();
 FILLCELL_X32 FILLER_104_1437 ();
 FILLCELL_X32 FILLER_104_1469 ();
 FILLCELL_X32 FILLER_104_1501 ();
 FILLCELL_X32 FILLER_104_1533 ();
 FILLCELL_X32 FILLER_104_1565 ();
 FILLCELL_X16 FILLER_104_1597 ();
 FILLCELL_X1 FILLER_104_1613 ();
 FILLCELL_X1 FILLER_105_1 ();
 FILLCELL_X8 FILLER_105_8 ();
 FILLCELL_X2 FILLER_105_16 ();
 FILLCELL_X4 FILLER_105_22 ();
 FILLCELL_X2 FILLER_105_26 ();
 FILLCELL_X1 FILLER_105_28 ();
 FILLCELL_X8 FILLER_105_33 ();
 FILLCELL_X2 FILLER_105_41 ();
 FILLCELL_X32 FILLER_105_60 ();
 FILLCELL_X32 FILLER_105_92 ();
 FILLCELL_X32 FILLER_105_124 ();
 FILLCELL_X32 FILLER_105_156 ();
 FILLCELL_X32 FILLER_105_188 ();
 FILLCELL_X32 FILLER_105_220 ();
 FILLCELL_X32 FILLER_105_252 ();
 FILLCELL_X32 FILLER_105_284 ();
 FILLCELL_X32 FILLER_105_316 ();
 FILLCELL_X32 FILLER_105_348 ();
 FILLCELL_X32 FILLER_105_380 ();
 FILLCELL_X32 FILLER_105_412 ();
 FILLCELL_X32 FILLER_105_444 ();
 FILLCELL_X32 FILLER_105_476 ();
 FILLCELL_X32 FILLER_105_508 ();
 FILLCELL_X32 FILLER_105_540 ();
 FILLCELL_X32 FILLER_105_572 ();
 FILLCELL_X32 FILLER_105_604 ();
 FILLCELL_X32 FILLER_105_636 ();
 FILLCELL_X32 FILLER_105_668 ();
 FILLCELL_X32 FILLER_105_700 ();
 FILLCELL_X32 FILLER_105_732 ();
 FILLCELL_X16 FILLER_105_764 ();
 FILLCELL_X8 FILLER_105_780 ();
 FILLCELL_X4 FILLER_105_788 ();
 FILLCELL_X1 FILLER_105_792 ();
 FILLCELL_X4 FILLER_105_798 ();
 FILLCELL_X16 FILLER_105_809 ();
 FILLCELL_X4 FILLER_105_825 ();
 FILLCELL_X2 FILLER_105_829 ();
 FILLCELL_X4 FILLER_105_834 ();
 FILLCELL_X2 FILLER_105_838 ();
 FILLCELL_X1 FILLER_105_840 ();
 FILLCELL_X1 FILLER_105_848 ();
 FILLCELL_X8 FILLER_105_868 ();
 FILLCELL_X8 FILLER_105_884 ();
 FILLCELL_X1 FILLER_105_892 ();
 FILLCELL_X1 FILLER_105_900 ();
 FILLCELL_X8 FILLER_105_905 ();
 FILLCELL_X4 FILLER_105_913 ();
 FILLCELL_X2 FILLER_105_917 ();
 FILLCELL_X1 FILLER_105_919 ();
 FILLCELL_X4 FILLER_105_924 ();
 FILLCELL_X4 FILLER_105_932 ();
 FILLCELL_X32 FILLER_105_945 ();
 FILLCELL_X32 FILLER_105_977 ();
 FILLCELL_X32 FILLER_105_1009 ();
 FILLCELL_X32 FILLER_105_1041 ();
 FILLCELL_X32 FILLER_105_1073 ();
 FILLCELL_X32 FILLER_105_1105 ();
 FILLCELL_X32 FILLER_105_1137 ();
 FILLCELL_X32 FILLER_105_1169 ();
 FILLCELL_X32 FILLER_105_1201 ();
 FILLCELL_X16 FILLER_105_1233 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X2 FILLER_105_1584 ();
 FILLCELL_X1 FILLER_105_1586 ();
 FILLCELL_X16 FILLER_105_1590 ();
 FILLCELL_X8 FILLER_105_1606 ();
 FILLCELL_X2 FILLER_106_1 ();
 FILLCELL_X1 FILLER_106_3 ();
 FILLCELL_X1 FILLER_106_14 ();
 FILLCELL_X16 FILLER_106_23 ();
 FILLCELL_X4 FILLER_106_39 ();
 FILLCELL_X2 FILLER_106_43 ();
 FILLCELL_X1 FILLER_106_45 ();
 FILLCELL_X32 FILLER_106_59 ();
 FILLCELL_X32 FILLER_106_91 ();
 FILLCELL_X32 FILLER_106_123 ();
 FILLCELL_X32 FILLER_106_155 ();
 FILLCELL_X32 FILLER_106_187 ();
 FILLCELL_X32 FILLER_106_219 ();
 FILLCELL_X32 FILLER_106_251 ();
 FILLCELL_X32 FILLER_106_283 ();
 FILLCELL_X32 FILLER_106_315 ();
 FILLCELL_X32 FILLER_106_347 ();
 FILLCELL_X32 FILLER_106_379 ();
 FILLCELL_X32 FILLER_106_411 ();
 FILLCELL_X32 FILLER_106_443 ();
 FILLCELL_X32 FILLER_106_475 ();
 FILLCELL_X32 FILLER_106_507 ();
 FILLCELL_X32 FILLER_106_539 ();
 FILLCELL_X32 FILLER_106_571 ();
 FILLCELL_X16 FILLER_106_603 ();
 FILLCELL_X8 FILLER_106_619 ();
 FILLCELL_X4 FILLER_106_627 ();
 FILLCELL_X16 FILLER_106_632 ();
 FILLCELL_X4 FILLER_106_648 ();
 FILLCELL_X32 FILLER_106_662 ();
 FILLCELL_X32 FILLER_106_694 ();
 FILLCELL_X32 FILLER_106_726 ();
 FILLCELL_X32 FILLER_106_758 ();
 FILLCELL_X16 FILLER_106_790 ();
 FILLCELL_X4 FILLER_106_806 ();
 FILLCELL_X1 FILLER_106_810 ();
 FILLCELL_X16 FILLER_106_814 ();
 FILLCELL_X8 FILLER_106_830 ();
 FILLCELL_X4 FILLER_106_838 ();
 FILLCELL_X1 FILLER_106_842 ();
 FILLCELL_X2 FILLER_106_858 ();
 FILLCELL_X1 FILLER_106_860 ();
 FILLCELL_X1 FILLER_106_864 ();
 FILLCELL_X8 FILLER_106_868 ();
 FILLCELL_X4 FILLER_106_876 ();
 FILLCELL_X2 FILLER_106_880 ();
 FILLCELL_X4 FILLER_106_887 ();
 FILLCELL_X1 FILLER_106_891 ();
 FILLCELL_X8 FILLER_106_910 ();
 FILLCELL_X1 FILLER_106_918 ();
 FILLCELL_X2 FILLER_106_923 ();
 FILLCELL_X1 FILLER_106_932 ();
 FILLCELL_X32 FILLER_106_935 ();
 FILLCELL_X32 FILLER_106_967 ();
 FILLCELL_X32 FILLER_106_999 ();
 FILLCELL_X32 FILLER_106_1031 ();
 FILLCELL_X32 FILLER_106_1063 ();
 FILLCELL_X32 FILLER_106_1095 ();
 FILLCELL_X32 FILLER_106_1127 ();
 FILLCELL_X32 FILLER_106_1159 ();
 FILLCELL_X32 FILLER_106_1191 ();
 FILLCELL_X32 FILLER_106_1223 ();
 FILLCELL_X32 FILLER_106_1255 ();
 FILLCELL_X32 FILLER_106_1287 ();
 FILLCELL_X32 FILLER_106_1319 ();
 FILLCELL_X32 FILLER_106_1351 ();
 FILLCELL_X32 FILLER_106_1383 ();
 FILLCELL_X32 FILLER_106_1415 ();
 FILLCELL_X32 FILLER_106_1447 ();
 FILLCELL_X32 FILLER_106_1479 ();
 FILLCELL_X32 FILLER_106_1511 ();
 FILLCELL_X32 FILLER_106_1543 ();
 FILLCELL_X32 FILLER_106_1575 ();
 FILLCELL_X4 FILLER_106_1607 ();
 FILLCELL_X2 FILLER_106_1611 ();
 FILLCELL_X1 FILLER_106_1613 ();
 FILLCELL_X8 FILLER_107_1 ();
 FILLCELL_X2 FILLER_107_12 ();
 FILLCELL_X1 FILLER_107_14 ();
 FILLCELL_X2 FILLER_107_18 ();
 FILLCELL_X1 FILLER_107_20 ();
 FILLCELL_X8 FILLER_107_32 ();
 FILLCELL_X4 FILLER_107_40 ();
 FILLCELL_X1 FILLER_107_44 ();
 FILLCELL_X8 FILLER_107_49 ();
 FILLCELL_X4 FILLER_107_57 ();
 FILLCELL_X2 FILLER_107_61 ();
 FILLCELL_X1 FILLER_107_63 ();
 FILLCELL_X4 FILLER_107_69 ();
 FILLCELL_X1 FILLER_107_73 ();
 FILLCELL_X32 FILLER_107_81 ();
 FILLCELL_X32 FILLER_107_113 ();
 FILLCELL_X32 FILLER_107_145 ();
 FILLCELL_X32 FILLER_107_177 ();
 FILLCELL_X32 FILLER_107_209 ();
 FILLCELL_X32 FILLER_107_241 ();
 FILLCELL_X32 FILLER_107_273 ();
 FILLCELL_X32 FILLER_107_305 ();
 FILLCELL_X32 FILLER_107_337 ();
 FILLCELL_X32 FILLER_107_369 ();
 FILLCELL_X32 FILLER_107_401 ();
 FILLCELL_X32 FILLER_107_433 ();
 FILLCELL_X32 FILLER_107_465 ();
 FILLCELL_X32 FILLER_107_497 ();
 FILLCELL_X32 FILLER_107_529 ();
 FILLCELL_X32 FILLER_107_561 ();
 FILLCELL_X32 FILLER_107_593 ();
 FILLCELL_X32 FILLER_107_625 ();
 FILLCELL_X32 FILLER_107_657 ();
 FILLCELL_X8 FILLER_107_689 ();
 FILLCELL_X4 FILLER_107_697 ();
 FILLCELL_X2 FILLER_107_701 ();
 FILLCELL_X32 FILLER_107_707 ();
 FILLCELL_X32 FILLER_107_739 ();
 FILLCELL_X32 FILLER_107_771 ();
 FILLCELL_X4 FILLER_107_803 ();
 FILLCELL_X2 FILLER_107_810 ();
 FILLCELL_X1 FILLER_107_812 ();
 FILLCELL_X16 FILLER_107_831 ();
 FILLCELL_X2 FILLER_107_847 ();
 FILLCELL_X4 FILLER_107_853 ();
 FILLCELL_X1 FILLER_107_857 ();
 FILLCELL_X8 FILLER_107_867 ();
 FILLCELL_X4 FILLER_107_875 ();
 FILLCELL_X4 FILLER_107_886 ();
 FILLCELL_X2 FILLER_107_890 ();
 FILLCELL_X1 FILLER_107_892 ();
 FILLCELL_X32 FILLER_107_905 ();
 FILLCELL_X32 FILLER_107_937 ();
 FILLCELL_X32 FILLER_107_969 ();
 FILLCELL_X32 FILLER_107_1001 ();
 FILLCELL_X32 FILLER_107_1033 ();
 FILLCELL_X32 FILLER_107_1065 ();
 FILLCELL_X32 FILLER_107_1097 ();
 FILLCELL_X32 FILLER_107_1129 ();
 FILLCELL_X32 FILLER_107_1161 ();
 FILLCELL_X32 FILLER_107_1193 ();
 FILLCELL_X32 FILLER_107_1225 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X16 FILLER_107_1584 ();
 FILLCELL_X2 FILLER_107_1600 ();
 FILLCELL_X8 FILLER_107_1606 ();
 FILLCELL_X4 FILLER_108_1 ();
 FILLCELL_X2 FILLER_108_5 ();
 FILLCELL_X4 FILLER_108_10 ();
 FILLCELL_X2 FILLER_108_14 ();
 FILLCELL_X32 FILLER_108_32 ();
 FILLCELL_X1 FILLER_108_64 ();
 FILLCELL_X1 FILLER_108_71 ();
 FILLCELL_X1 FILLER_108_74 ();
 FILLCELL_X8 FILLER_108_88 ();
 FILLCELL_X1 FILLER_108_96 ();
 FILLCELL_X32 FILLER_108_102 ();
 FILLCELL_X32 FILLER_108_134 ();
 FILLCELL_X32 FILLER_108_166 ();
 FILLCELL_X32 FILLER_108_198 ();
 FILLCELL_X32 FILLER_108_230 ();
 FILLCELL_X32 FILLER_108_262 ();
 FILLCELL_X32 FILLER_108_294 ();
 FILLCELL_X32 FILLER_108_326 ();
 FILLCELL_X32 FILLER_108_358 ();
 FILLCELL_X32 FILLER_108_390 ();
 FILLCELL_X32 FILLER_108_422 ();
 FILLCELL_X32 FILLER_108_454 ();
 FILLCELL_X32 FILLER_108_486 ();
 FILLCELL_X32 FILLER_108_518 ();
 FILLCELL_X32 FILLER_108_550 ();
 FILLCELL_X32 FILLER_108_582 ();
 FILLCELL_X16 FILLER_108_614 ();
 FILLCELL_X1 FILLER_108_630 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X16 FILLER_108_728 ();
 FILLCELL_X4 FILLER_108_744 ();
 FILLCELL_X32 FILLER_108_753 ();
 FILLCELL_X4 FILLER_108_785 ();
 FILLCELL_X2 FILLER_108_796 ();
 FILLCELL_X1 FILLER_108_798 ();
 FILLCELL_X4 FILLER_108_816 ();
 FILLCELL_X8 FILLER_108_829 ();
 FILLCELL_X4 FILLER_108_837 ();
 FILLCELL_X1 FILLER_108_841 ();
 FILLCELL_X4 FILLER_108_866 ();
 FILLCELL_X32 FILLER_108_889 ();
 FILLCELL_X2 FILLER_108_942 ();
 FILLCELL_X2 FILLER_108_964 ();
 FILLCELL_X8 FILLER_108_975 ();
 FILLCELL_X2 FILLER_108_983 ();
 FILLCELL_X1 FILLER_108_985 ();
 FILLCELL_X32 FILLER_108_996 ();
 FILLCELL_X32 FILLER_108_1028 ();
 FILLCELL_X32 FILLER_108_1060 ();
 FILLCELL_X32 FILLER_108_1092 ();
 FILLCELL_X32 FILLER_108_1124 ();
 FILLCELL_X32 FILLER_108_1156 ();
 FILLCELL_X32 FILLER_108_1188 ();
 FILLCELL_X32 FILLER_108_1220 ();
 FILLCELL_X32 FILLER_108_1252 ();
 FILLCELL_X32 FILLER_108_1284 ();
 FILLCELL_X32 FILLER_108_1316 ();
 FILLCELL_X32 FILLER_108_1348 ();
 FILLCELL_X32 FILLER_108_1380 ();
 FILLCELL_X32 FILLER_108_1412 ();
 FILLCELL_X32 FILLER_108_1444 ();
 FILLCELL_X32 FILLER_108_1476 ();
 FILLCELL_X32 FILLER_108_1508 ();
 FILLCELL_X32 FILLER_108_1540 ();
 FILLCELL_X2 FILLER_108_1572 ();
 FILLCELL_X32 FILLER_108_1578 ();
 FILLCELL_X4 FILLER_108_1610 ();
 FILLCELL_X32 FILLER_109_19 ();
 FILLCELL_X1 FILLER_109_51 ();
 FILLCELL_X4 FILLER_109_58 ();
 FILLCELL_X16 FILLER_109_66 ();
 FILLCELL_X4 FILLER_109_88 ();
 FILLCELL_X8 FILLER_109_110 ();
 FILLCELL_X2 FILLER_109_118 ();
 FILLCELL_X1 FILLER_109_120 ();
 FILLCELL_X32 FILLER_109_139 ();
 FILLCELL_X32 FILLER_109_171 ();
 FILLCELL_X32 FILLER_109_203 ();
 FILLCELL_X32 FILLER_109_235 ();
 FILLCELL_X32 FILLER_109_267 ();
 FILLCELL_X32 FILLER_109_299 ();
 FILLCELL_X32 FILLER_109_331 ();
 FILLCELL_X32 FILLER_109_363 ();
 FILLCELL_X32 FILLER_109_395 ();
 FILLCELL_X32 FILLER_109_427 ();
 FILLCELL_X32 FILLER_109_459 ();
 FILLCELL_X32 FILLER_109_491 ();
 FILLCELL_X32 FILLER_109_523 ();
 FILLCELL_X32 FILLER_109_555 ();
 FILLCELL_X32 FILLER_109_587 ();
 FILLCELL_X32 FILLER_109_619 ();
 FILLCELL_X32 FILLER_109_651 ();
 FILLCELL_X32 FILLER_109_683 ();
 FILLCELL_X32 FILLER_109_715 ();
 FILLCELL_X16 FILLER_109_747 ();
 FILLCELL_X1 FILLER_109_763 ();
 FILLCELL_X4 FILLER_109_777 ();
 FILLCELL_X2 FILLER_109_781 ();
 FILLCELL_X16 FILLER_109_823 ();
 FILLCELL_X4 FILLER_109_839 ();
 FILLCELL_X2 FILLER_109_843 ();
 FILLCELL_X16 FILLER_109_855 ();
 FILLCELL_X8 FILLER_109_871 ();
 FILLCELL_X4 FILLER_109_879 ();
 FILLCELL_X8 FILLER_109_888 ();
 FILLCELL_X4 FILLER_109_896 ();
 FILLCELL_X1 FILLER_109_900 ();
 FILLCELL_X16 FILLER_109_911 ();
 FILLCELL_X1 FILLER_109_927 ();
 FILLCELL_X16 FILLER_109_931 ();
 FILLCELL_X1 FILLER_109_947 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X16 FILLER_109_1587 ();
 FILLCELL_X4 FILLER_109_1603 ();
 FILLCELL_X4 FILLER_109_1610 ();
 FILLCELL_X16 FILLER_110_4 ();
 FILLCELL_X8 FILLER_110_20 ();
 FILLCELL_X2 FILLER_110_28 ();
 FILLCELL_X1 FILLER_110_30 ();
 FILLCELL_X16 FILLER_110_35 ();
 FILLCELL_X1 FILLER_110_60 ();
 FILLCELL_X8 FILLER_110_92 ();
 FILLCELL_X4 FILLER_110_100 ();
 FILLCELL_X2 FILLER_110_104 ();
 FILLCELL_X1 FILLER_110_106 ();
 FILLCELL_X2 FILLER_110_111 ();
 FILLCELL_X1 FILLER_110_116 ();
 FILLCELL_X4 FILLER_110_136 ();
 FILLCELL_X1 FILLER_110_140 ();
 FILLCELL_X32 FILLER_110_150 ();
 FILLCELL_X32 FILLER_110_182 ();
 FILLCELL_X32 FILLER_110_214 ();
 FILLCELL_X32 FILLER_110_246 ();
 FILLCELL_X32 FILLER_110_278 ();
 FILLCELL_X32 FILLER_110_310 ();
 FILLCELL_X32 FILLER_110_342 ();
 FILLCELL_X32 FILLER_110_374 ();
 FILLCELL_X32 FILLER_110_406 ();
 FILLCELL_X32 FILLER_110_438 ();
 FILLCELL_X32 FILLER_110_470 ();
 FILLCELL_X32 FILLER_110_502 ();
 FILLCELL_X32 FILLER_110_534 ();
 FILLCELL_X32 FILLER_110_566 ();
 FILLCELL_X32 FILLER_110_598 ();
 FILLCELL_X1 FILLER_110_630 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X8 FILLER_110_696 ();
 FILLCELL_X4 FILLER_110_704 ();
 FILLCELL_X2 FILLER_110_708 ();
 FILLCELL_X32 FILLER_110_724 ();
 FILLCELL_X4 FILLER_110_756 ();
 FILLCELL_X2 FILLER_110_760 ();
 FILLCELL_X1 FILLER_110_762 ();
 FILLCELL_X16 FILLER_110_783 ();
 FILLCELL_X8 FILLER_110_799 ();
 FILLCELL_X2 FILLER_110_807 ();
 FILLCELL_X4 FILLER_110_816 ();
 FILLCELL_X1 FILLER_110_820 ();
 FILLCELL_X4 FILLER_110_830 ();
 FILLCELL_X1 FILLER_110_834 ();
 FILLCELL_X1 FILLER_110_839 ();
 FILLCELL_X16 FILLER_110_842 ();
 FILLCELL_X1 FILLER_110_858 ();
 FILLCELL_X1 FILLER_110_870 ();
 FILLCELL_X2 FILLER_110_873 ();
 FILLCELL_X32 FILLER_110_883 ();
 FILLCELL_X16 FILLER_110_915 ();
 FILLCELL_X4 FILLER_110_931 ();
 FILLCELL_X8 FILLER_110_943 ();
 FILLCELL_X2 FILLER_110_951 ();
 FILLCELL_X1 FILLER_110_953 ();
 FILLCELL_X4 FILLER_110_958 ();
 FILLCELL_X32 FILLER_110_964 ();
 FILLCELL_X32 FILLER_110_996 ();
 FILLCELL_X16 FILLER_110_1028 ();
 FILLCELL_X8 FILLER_110_1044 ();
 FILLCELL_X4 FILLER_110_1052 ();
 FILLCELL_X1 FILLER_110_1056 ();
 FILLCELL_X16 FILLER_110_1061 ();
 FILLCELL_X2 FILLER_110_1077 ();
 FILLCELL_X32 FILLER_110_1089 ();
 FILLCELL_X32 FILLER_110_1121 ();
 FILLCELL_X32 FILLER_110_1153 ();
 FILLCELL_X32 FILLER_110_1185 ();
 FILLCELL_X32 FILLER_110_1217 ();
 FILLCELL_X32 FILLER_110_1249 ();
 FILLCELL_X32 FILLER_110_1281 ();
 FILLCELL_X32 FILLER_110_1313 ();
 FILLCELL_X32 FILLER_110_1345 ();
 FILLCELL_X32 FILLER_110_1377 ();
 FILLCELL_X32 FILLER_110_1409 ();
 FILLCELL_X32 FILLER_110_1441 ();
 FILLCELL_X32 FILLER_110_1473 ();
 FILLCELL_X32 FILLER_110_1505 ();
 FILLCELL_X32 FILLER_110_1537 ();
 FILLCELL_X4 FILLER_110_1569 ();
 FILLCELL_X2 FILLER_110_1573 ();
 FILLCELL_X1 FILLER_110_1575 ();
 FILLCELL_X16 FILLER_110_1584 ();
 FILLCELL_X8 FILLER_110_1600 ();
 FILLCELL_X4 FILLER_110_1608 ();
 FILLCELL_X2 FILLER_110_1612 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X16 FILLER_111_65 ();
 FILLCELL_X8 FILLER_111_81 ();
 FILLCELL_X4 FILLER_111_89 ();
 FILLCELL_X2 FILLER_111_93 ();
 FILLCELL_X1 FILLER_111_95 ();
 FILLCELL_X8 FILLER_111_100 ();
 FILLCELL_X8 FILLER_111_117 ();
 FILLCELL_X4 FILLER_111_125 ();
 FILLCELL_X1 FILLER_111_129 ();
 FILLCELL_X4 FILLER_111_134 ();
 FILLCELL_X2 FILLER_111_138 ();
 FILLCELL_X4 FILLER_111_160 ();
 FILLCELL_X1 FILLER_111_164 ();
 FILLCELL_X4 FILLER_111_174 ();
 FILLCELL_X1 FILLER_111_178 ();
 FILLCELL_X8 FILLER_111_182 ();
 FILLCELL_X4 FILLER_111_190 ();
 FILLCELL_X2 FILLER_111_194 ();
 FILLCELL_X32 FILLER_111_210 ();
 FILLCELL_X32 FILLER_111_242 ();
 FILLCELL_X32 FILLER_111_274 ();
 FILLCELL_X32 FILLER_111_306 ();
 FILLCELL_X32 FILLER_111_338 ();
 FILLCELL_X32 FILLER_111_370 ();
 FILLCELL_X32 FILLER_111_402 ();
 FILLCELL_X32 FILLER_111_434 ();
 FILLCELL_X32 FILLER_111_466 ();
 FILLCELL_X32 FILLER_111_498 ();
 FILLCELL_X32 FILLER_111_530 ();
 FILLCELL_X32 FILLER_111_562 ();
 FILLCELL_X32 FILLER_111_594 ();
 FILLCELL_X32 FILLER_111_626 ();
 FILLCELL_X4 FILLER_111_658 ();
 FILLCELL_X2 FILLER_111_662 ();
 FILLCELL_X2 FILLER_111_667 ();
 FILLCELL_X16 FILLER_111_678 ();
 FILLCELL_X8 FILLER_111_694 ();
 FILLCELL_X2 FILLER_111_702 ();
 FILLCELL_X1 FILLER_111_704 ();
 FILLCELL_X2 FILLER_111_708 ();
 FILLCELL_X2 FILLER_111_726 ();
 FILLCELL_X1 FILLER_111_728 ();
 FILLCELL_X8 FILLER_111_746 ();
 FILLCELL_X4 FILLER_111_754 ();
 FILLCELL_X2 FILLER_111_758 ();
 FILLCELL_X16 FILLER_111_763 ();
 FILLCELL_X4 FILLER_111_779 ();
 FILLCELL_X4 FILLER_111_792 ();
 FILLCELL_X1 FILLER_111_796 ();
 FILLCELL_X4 FILLER_111_806 ();
 FILLCELL_X2 FILLER_111_810 ();
 FILLCELL_X1 FILLER_111_812 ();
 FILLCELL_X8 FILLER_111_822 ();
 FILLCELL_X2 FILLER_111_830 ();
 FILLCELL_X1 FILLER_111_832 ();
 FILLCELL_X2 FILLER_111_844 ();
 FILLCELL_X1 FILLER_111_858 ();
 FILLCELL_X2 FILLER_111_862 ();
 FILLCELL_X2 FILLER_111_867 ();
 FILLCELL_X1 FILLER_111_869 ();
 FILLCELL_X4 FILLER_111_882 ();
 FILLCELL_X2 FILLER_111_886 ();
 FILLCELL_X16 FILLER_111_900 ();
 FILLCELL_X1 FILLER_111_916 ();
 FILLCELL_X2 FILLER_111_927 ();
 FILLCELL_X16 FILLER_111_938 ();
 FILLCELL_X4 FILLER_111_954 ();
 FILLCELL_X1 FILLER_111_958 ();
 FILLCELL_X2 FILLER_111_961 ();
 FILLCELL_X4 FILLER_111_971 ();
 FILLCELL_X2 FILLER_111_977 ();
 FILLCELL_X1 FILLER_111_979 ();
 FILLCELL_X32 FILLER_111_984 ();
 FILLCELL_X32 FILLER_111_1016 ();
 FILLCELL_X32 FILLER_111_1048 ();
 FILLCELL_X32 FILLER_111_1080 ();
 FILLCELL_X32 FILLER_111_1112 ();
 FILLCELL_X32 FILLER_111_1144 ();
 FILLCELL_X32 FILLER_111_1176 ();
 FILLCELL_X32 FILLER_111_1208 ();
 FILLCELL_X16 FILLER_111_1240 ();
 FILLCELL_X4 FILLER_111_1256 ();
 FILLCELL_X2 FILLER_111_1260 ();
 FILLCELL_X1 FILLER_111_1262 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X16 FILLER_111_1584 ();
 FILLCELL_X8 FILLER_111_1600 ();
 FILLCELL_X4 FILLER_111_1608 ();
 FILLCELL_X2 FILLER_111_1612 ();
 FILLCELL_X16 FILLER_112_1 ();
 FILLCELL_X2 FILLER_112_17 ();
 FILLCELL_X32 FILLER_112_27 ();
 FILLCELL_X16 FILLER_112_59 ();
 FILLCELL_X8 FILLER_112_75 ();
 FILLCELL_X4 FILLER_112_83 ();
 FILLCELL_X1 FILLER_112_87 ();
 FILLCELL_X8 FILLER_112_102 ();
 FILLCELL_X8 FILLER_112_117 ();
 FILLCELL_X4 FILLER_112_125 ();
 FILLCELL_X8 FILLER_112_133 ();
 FILLCELL_X4 FILLER_112_150 ();
 FILLCELL_X1 FILLER_112_154 ();
 FILLCELL_X32 FILLER_112_160 ();
 FILLCELL_X32 FILLER_112_192 ();
 FILLCELL_X32 FILLER_112_224 ();
 FILLCELL_X32 FILLER_112_256 ();
 FILLCELL_X32 FILLER_112_288 ();
 FILLCELL_X32 FILLER_112_320 ();
 FILLCELL_X32 FILLER_112_352 ();
 FILLCELL_X32 FILLER_112_384 ();
 FILLCELL_X32 FILLER_112_416 ();
 FILLCELL_X32 FILLER_112_448 ();
 FILLCELL_X32 FILLER_112_480 ();
 FILLCELL_X32 FILLER_112_512 ();
 FILLCELL_X32 FILLER_112_544 ();
 FILLCELL_X32 FILLER_112_576 ();
 FILLCELL_X16 FILLER_112_608 ();
 FILLCELL_X4 FILLER_112_624 ();
 FILLCELL_X2 FILLER_112_628 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X4 FILLER_112_696 ();
 FILLCELL_X16 FILLER_112_707 ();
 FILLCELL_X2 FILLER_112_729 ();
 FILLCELL_X8 FILLER_112_733 ();
 FILLCELL_X4 FILLER_112_741 ();
 FILLCELL_X2 FILLER_112_745 ();
 FILLCELL_X1 FILLER_112_747 ();
 FILLCELL_X2 FILLER_112_752 ();
 FILLCELL_X8 FILLER_112_772 ();
 FILLCELL_X8 FILLER_112_787 ();
 FILLCELL_X4 FILLER_112_795 ();
 FILLCELL_X2 FILLER_112_799 ();
 FILLCELL_X8 FILLER_112_805 ();
 FILLCELL_X2 FILLER_112_813 ();
 FILLCELL_X1 FILLER_112_815 ();
 FILLCELL_X32 FILLER_112_822 ();
 FILLCELL_X8 FILLER_112_854 ();
 FILLCELL_X4 FILLER_112_862 ();
 FILLCELL_X2 FILLER_112_866 ();
 FILLCELL_X4 FILLER_112_874 ();
 FILLCELL_X16 FILLER_112_885 ();
 FILLCELL_X1 FILLER_112_901 ();
 FILLCELL_X2 FILLER_112_939 ();
 FILLCELL_X1 FILLER_112_941 ();
 FILLCELL_X1 FILLER_112_951 ();
 FILLCELL_X2 FILLER_112_963 ();
 FILLCELL_X1 FILLER_112_965 ();
 FILLCELL_X2 FILLER_112_975 ();
 FILLCELL_X1 FILLER_112_981 ();
 FILLCELL_X2 FILLER_112_986 ();
 FILLCELL_X8 FILLER_112_990 ();
 FILLCELL_X4 FILLER_112_998 ();
 FILLCELL_X2 FILLER_112_1002 ();
 FILLCELL_X1 FILLER_112_1004 ();
 FILLCELL_X16 FILLER_112_1011 ();
 FILLCELL_X8 FILLER_112_1027 ();
 FILLCELL_X4 FILLER_112_1035 ();
 FILLCELL_X2 FILLER_112_1039 ();
 FILLCELL_X32 FILLER_112_1051 ();
 FILLCELL_X32 FILLER_112_1083 ();
 FILLCELL_X32 FILLER_112_1115 ();
 FILLCELL_X32 FILLER_112_1147 ();
 FILLCELL_X32 FILLER_112_1179 ();
 FILLCELL_X32 FILLER_112_1211 ();
 FILLCELL_X32 FILLER_112_1243 ();
 FILLCELL_X32 FILLER_112_1275 ();
 FILLCELL_X32 FILLER_112_1307 ();
 FILLCELL_X32 FILLER_112_1339 ();
 FILLCELL_X32 FILLER_112_1371 ();
 FILLCELL_X32 FILLER_112_1403 ();
 FILLCELL_X32 FILLER_112_1435 ();
 FILLCELL_X32 FILLER_112_1467 ();
 FILLCELL_X32 FILLER_112_1499 ();
 FILLCELL_X32 FILLER_112_1531 ();
 FILLCELL_X8 FILLER_112_1563 ();
 FILLCELL_X4 FILLER_112_1571 ();
 FILLCELL_X1 FILLER_112_1575 ();
 FILLCELL_X32 FILLER_112_1579 ();
 FILLCELL_X2 FILLER_112_1611 ();
 FILLCELL_X1 FILLER_112_1613 ();
 FILLCELL_X1 FILLER_113_14 ();
 FILLCELL_X32 FILLER_113_19 ();
 FILLCELL_X32 FILLER_113_51 ();
 FILLCELL_X16 FILLER_113_83 ();
 FILLCELL_X4 FILLER_113_99 ();
 FILLCELL_X2 FILLER_113_103 ();
 FILLCELL_X1 FILLER_113_105 ();
 FILLCELL_X8 FILLER_113_132 ();
 FILLCELL_X1 FILLER_113_140 ();
 FILLCELL_X16 FILLER_113_145 ();
 FILLCELL_X2 FILLER_113_161 ();
 FILLCELL_X16 FILLER_113_176 ();
 FILLCELL_X8 FILLER_113_192 ();
 FILLCELL_X32 FILLER_113_210 ();
 FILLCELL_X32 FILLER_113_242 ();
 FILLCELL_X32 FILLER_113_274 ();
 FILLCELL_X32 FILLER_113_306 ();
 FILLCELL_X32 FILLER_113_338 ();
 FILLCELL_X32 FILLER_113_370 ();
 FILLCELL_X32 FILLER_113_402 ();
 FILLCELL_X32 FILLER_113_434 ();
 FILLCELL_X32 FILLER_113_466 ();
 FILLCELL_X32 FILLER_113_498 ();
 FILLCELL_X32 FILLER_113_530 ();
 FILLCELL_X32 FILLER_113_562 ();
 FILLCELL_X32 FILLER_113_594 ();
 FILLCELL_X32 FILLER_113_626 ();
 FILLCELL_X32 FILLER_113_658 ();
 FILLCELL_X16 FILLER_113_690 ();
 FILLCELL_X8 FILLER_113_706 ();
 FILLCELL_X16 FILLER_113_737 ();
 FILLCELL_X8 FILLER_113_753 ();
 FILLCELL_X4 FILLER_113_761 ();
 FILLCELL_X2 FILLER_113_765 ();
 FILLCELL_X4 FILLER_113_774 ();
 FILLCELL_X2 FILLER_113_778 ();
 FILLCELL_X1 FILLER_113_780 ();
 FILLCELL_X4 FILLER_113_784 ();
 FILLCELL_X2 FILLER_113_788 ();
 FILLCELL_X4 FILLER_113_794 ();
 FILLCELL_X1 FILLER_113_798 ();
 FILLCELL_X8 FILLER_113_806 ();
 FILLCELL_X2 FILLER_113_814 ();
 FILLCELL_X16 FILLER_113_819 ();
 FILLCELL_X8 FILLER_113_835 ();
 FILLCELL_X2 FILLER_113_843 ();
 FILLCELL_X32 FILLER_113_847 ();
 FILLCELL_X4 FILLER_113_879 ();
 FILLCELL_X2 FILLER_113_883 ();
 FILLCELL_X16 FILLER_113_892 ();
 FILLCELL_X4 FILLER_113_908 ();
 FILLCELL_X2 FILLER_113_912 ();
 FILLCELL_X8 FILLER_113_926 ();
 FILLCELL_X2 FILLER_113_934 ();
 FILLCELL_X16 FILLER_113_939 ();
 FILLCELL_X4 FILLER_113_955 ();
 FILLCELL_X1 FILLER_113_959 ();
 FILLCELL_X1 FILLER_113_964 ();
 FILLCELL_X8 FILLER_113_967 ();
 FILLCELL_X2 FILLER_113_975 ();
 FILLCELL_X4 FILLER_113_981 ();
 FILLCELL_X4 FILLER_113_988 ();
 FILLCELL_X2 FILLER_113_992 ();
 FILLCELL_X1 FILLER_113_994 ();
 FILLCELL_X2 FILLER_113_1005 ();
 FILLCELL_X1 FILLER_113_1007 ();
 FILLCELL_X4 FILLER_113_1021 ();
 FILLCELL_X2 FILLER_113_1025 ();
 FILLCELL_X32 FILLER_113_1037 ();
 FILLCELL_X32 FILLER_113_1069 ();
 FILLCELL_X32 FILLER_113_1101 ();
 FILLCELL_X32 FILLER_113_1133 ();
 FILLCELL_X32 FILLER_113_1165 ();
 FILLCELL_X32 FILLER_113_1197 ();
 FILLCELL_X32 FILLER_113_1229 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X16 FILLER_113_1552 ();
 FILLCELL_X8 FILLER_113_1568 ();
 FILLCELL_X4 FILLER_113_1576 ();
 FILLCELL_X2 FILLER_113_1580 ();
 FILLCELL_X1 FILLER_113_1582 ();
 FILLCELL_X16 FILLER_113_1586 ();
 FILLCELL_X8 FILLER_113_1602 ();
 FILLCELL_X4 FILLER_113_1610 ();
 FILLCELL_X2 FILLER_114_1 ();
 FILLCELL_X1 FILLER_114_3 ();
 FILLCELL_X32 FILLER_114_7 ();
 FILLCELL_X32 FILLER_114_39 ();
 FILLCELL_X32 FILLER_114_71 ();
 FILLCELL_X16 FILLER_114_103 ();
 FILLCELL_X4 FILLER_114_119 ();
 FILLCELL_X1 FILLER_114_123 ();
 FILLCELL_X32 FILLER_114_127 ();
 FILLCELL_X32 FILLER_114_159 ();
 FILLCELL_X32 FILLER_114_191 ();
 FILLCELL_X32 FILLER_114_223 ();
 FILLCELL_X32 FILLER_114_255 ();
 FILLCELL_X32 FILLER_114_287 ();
 FILLCELL_X32 FILLER_114_319 ();
 FILLCELL_X32 FILLER_114_351 ();
 FILLCELL_X32 FILLER_114_383 ();
 FILLCELL_X32 FILLER_114_415 ();
 FILLCELL_X32 FILLER_114_447 ();
 FILLCELL_X32 FILLER_114_479 ();
 FILLCELL_X32 FILLER_114_511 ();
 FILLCELL_X32 FILLER_114_543 ();
 FILLCELL_X32 FILLER_114_575 ();
 FILLCELL_X16 FILLER_114_607 ();
 FILLCELL_X8 FILLER_114_623 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X16 FILLER_114_664 ();
 FILLCELL_X8 FILLER_114_680 ();
 FILLCELL_X4 FILLER_114_688 ();
 FILLCELL_X1 FILLER_114_692 ();
 FILLCELL_X32 FILLER_114_698 ();
 FILLCELL_X8 FILLER_114_730 ();
 FILLCELL_X2 FILLER_114_738 ();
 FILLCELL_X1 FILLER_114_740 ();
 FILLCELL_X16 FILLER_114_746 ();
 FILLCELL_X8 FILLER_114_762 ();
 FILLCELL_X4 FILLER_114_770 ();
 FILLCELL_X1 FILLER_114_774 ();
 FILLCELL_X2 FILLER_114_785 ();
 FILLCELL_X8 FILLER_114_796 ();
 FILLCELL_X1 FILLER_114_804 ();
 FILLCELL_X2 FILLER_114_813 ();
 FILLCELL_X32 FILLER_114_826 ();
 FILLCELL_X32 FILLER_114_858 ();
 FILLCELL_X16 FILLER_114_890 ();
 FILLCELL_X4 FILLER_114_906 ();
 FILLCELL_X1 FILLER_114_910 ();
 FILLCELL_X4 FILLER_114_924 ();
 FILLCELL_X2 FILLER_114_928 ();
 FILLCELL_X1 FILLER_114_930 ();
 FILLCELL_X2 FILLER_114_940 ();
 FILLCELL_X16 FILLER_114_958 ();
 FILLCELL_X4 FILLER_114_974 ();
 FILLCELL_X2 FILLER_114_978 ();
 FILLCELL_X1 FILLER_114_980 ();
 FILLCELL_X2 FILLER_114_992 ();
 FILLCELL_X32 FILLER_114_997 ();
 FILLCELL_X32 FILLER_114_1029 ();
 FILLCELL_X32 FILLER_114_1061 ();
 FILLCELL_X32 FILLER_114_1093 ();
 FILLCELL_X32 FILLER_114_1125 ();
 FILLCELL_X32 FILLER_114_1157 ();
 FILLCELL_X32 FILLER_114_1189 ();
 FILLCELL_X32 FILLER_114_1221 ();
 FILLCELL_X32 FILLER_114_1253 ();
 FILLCELL_X32 FILLER_114_1285 ();
 FILLCELL_X32 FILLER_114_1317 ();
 FILLCELL_X32 FILLER_114_1349 ();
 FILLCELL_X32 FILLER_114_1381 ();
 FILLCELL_X32 FILLER_114_1413 ();
 FILLCELL_X32 FILLER_114_1445 ();
 FILLCELL_X32 FILLER_114_1477 ();
 FILLCELL_X32 FILLER_114_1509 ();
 FILLCELL_X32 FILLER_114_1541 ();
 FILLCELL_X2 FILLER_114_1573 ();
 FILLCELL_X32 FILLER_114_1578 ();
 FILLCELL_X4 FILLER_114_1610 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X16 FILLER_115_641 ();
 FILLCELL_X8 FILLER_115_657 ();
 FILLCELL_X4 FILLER_115_665 ();
 FILLCELL_X16 FILLER_115_676 ();
 FILLCELL_X8 FILLER_115_692 ();
 FILLCELL_X4 FILLER_115_700 ();
 FILLCELL_X2 FILLER_115_704 ();
 FILLCELL_X32 FILLER_115_713 ();
 FILLCELL_X8 FILLER_115_745 ();
 FILLCELL_X4 FILLER_115_753 ();
 FILLCELL_X1 FILLER_115_764 ();
 FILLCELL_X16 FILLER_115_770 ();
 FILLCELL_X8 FILLER_115_786 ();
 FILLCELL_X1 FILLER_115_794 ();
 FILLCELL_X32 FILLER_115_816 ();
 FILLCELL_X32 FILLER_115_848 ();
 FILLCELL_X32 FILLER_115_880 ();
 FILLCELL_X8 FILLER_115_912 ();
 FILLCELL_X1 FILLER_115_928 ();
 FILLCELL_X1 FILLER_115_932 ();
 FILLCELL_X16 FILLER_115_937 ();
 FILLCELL_X8 FILLER_115_953 ();
 FILLCELL_X2 FILLER_115_961 ();
 FILLCELL_X1 FILLER_115_963 ();
 FILLCELL_X16 FILLER_115_972 ();
 FILLCELL_X8 FILLER_115_988 ();
 FILLCELL_X4 FILLER_115_996 ();
 FILLCELL_X2 FILLER_115_1004 ();
 FILLCELL_X1 FILLER_115_1006 ();
 FILLCELL_X8 FILLER_115_1011 ();
 FILLCELL_X32 FILLER_115_1026 ();
 FILLCELL_X32 FILLER_115_1058 ();
 FILLCELL_X32 FILLER_115_1090 ();
 FILLCELL_X32 FILLER_115_1122 ();
 FILLCELL_X32 FILLER_115_1154 ();
 FILLCELL_X32 FILLER_115_1186 ();
 FILLCELL_X32 FILLER_115_1218 ();
 FILLCELL_X8 FILLER_115_1250 ();
 FILLCELL_X4 FILLER_115_1258 ();
 FILLCELL_X1 FILLER_115_1262 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X16 FILLER_115_1552 ();
 FILLCELL_X2 FILLER_115_1568 ();
 FILLCELL_X1 FILLER_115_1570 ();
 FILLCELL_X2 FILLER_115_1575 ();
 FILLCELL_X8 FILLER_115_1581 ();
 FILLCELL_X8 FILLER_115_1596 ();
 FILLCELL_X4 FILLER_115_1604 ();
 FILLCELL_X1 FILLER_115_1613 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X8 FILLER_116_728 ();
 FILLCELL_X4 FILLER_116_736 ();
 FILLCELL_X32 FILLER_116_750 ();
 FILLCELL_X32 FILLER_116_782 ();
 FILLCELL_X32 FILLER_116_814 ();
 FILLCELL_X32 FILLER_116_846 ();
 FILLCELL_X32 FILLER_116_878 ();
 FILLCELL_X16 FILLER_116_910 ();
 FILLCELL_X4 FILLER_116_930 ();
 FILLCELL_X32 FILLER_116_947 ();
 FILLCELL_X16 FILLER_116_979 ();
 FILLCELL_X4 FILLER_116_995 ();
 FILLCELL_X2 FILLER_116_999 ();
 FILLCELL_X8 FILLER_116_1004 ();
 FILLCELL_X16 FILLER_116_1021 ();
 FILLCELL_X4 FILLER_116_1037 ();
 FILLCELL_X32 FILLER_116_1051 ();
 FILLCELL_X32 FILLER_116_1083 ();
 FILLCELL_X32 FILLER_116_1115 ();
 FILLCELL_X32 FILLER_116_1147 ();
 FILLCELL_X32 FILLER_116_1179 ();
 FILLCELL_X32 FILLER_116_1211 ();
 FILLCELL_X32 FILLER_116_1243 ();
 FILLCELL_X32 FILLER_116_1275 ();
 FILLCELL_X32 FILLER_116_1307 ();
 FILLCELL_X32 FILLER_116_1339 ();
 FILLCELL_X32 FILLER_116_1371 ();
 FILLCELL_X32 FILLER_116_1403 ();
 FILLCELL_X32 FILLER_116_1435 ();
 FILLCELL_X32 FILLER_116_1467 ();
 FILLCELL_X32 FILLER_116_1499 ();
 FILLCELL_X32 FILLER_116_1531 ();
 FILLCELL_X8 FILLER_116_1563 ();
 FILLCELL_X1 FILLER_116_1571 ();
 FILLCELL_X8 FILLER_116_1579 ();
 FILLCELL_X1 FILLER_116_1587 ();
 FILLCELL_X8 FILLER_116_1592 ();
 FILLCELL_X8 FILLER_116_1604 ();
 FILLCELL_X2 FILLER_116_1612 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X8 FILLER_117_673 ();
 FILLCELL_X2 FILLER_117_681 ();
 FILLCELL_X1 FILLER_117_683 ();
 FILLCELL_X16 FILLER_117_694 ();
 FILLCELL_X2 FILLER_117_710 ();
 FILLCELL_X1 FILLER_117_712 ();
 FILLCELL_X32 FILLER_117_723 ();
 FILLCELL_X1 FILLER_117_755 ();
 FILLCELL_X32 FILLER_117_766 ();
 FILLCELL_X8 FILLER_117_798 ();
 FILLCELL_X4 FILLER_117_806 ();
 FILLCELL_X1 FILLER_117_810 ();
 FILLCELL_X32 FILLER_117_827 ();
 FILLCELL_X32 FILLER_117_859 ();
 FILLCELL_X32 FILLER_117_891 ();
 FILLCELL_X32 FILLER_117_923 ();
 FILLCELL_X32 FILLER_117_955 ();
 FILLCELL_X32 FILLER_117_987 ();
 FILLCELL_X32 FILLER_117_1019 ();
 FILLCELL_X32 FILLER_117_1051 ();
 FILLCELL_X32 FILLER_117_1083 ();
 FILLCELL_X32 FILLER_117_1115 ();
 FILLCELL_X32 FILLER_117_1147 ();
 FILLCELL_X32 FILLER_117_1179 ();
 FILLCELL_X32 FILLER_117_1211 ();
 FILLCELL_X16 FILLER_117_1243 ();
 FILLCELL_X4 FILLER_117_1259 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X8 FILLER_117_1552 ();
 FILLCELL_X4 FILLER_117_1560 ();
 FILLCELL_X2 FILLER_117_1564 ();
 FILLCELL_X1 FILLER_117_1566 ();
 FILLCELL_X1 FILLER_117_1578 ();
 FILLCELL_X8 FILLER_117_1582 ();
 FILLCELL_X4 FILLER_117_1590 ();
 FILLCELL_X1 FILLER_117_1594 ();
 FILLCELL_X2 FILLER_117_1601 ();
 FILLCELL_X1 FILLER_117_1603 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X1 FILLER_118_792 ();
 FILLCELL_X8 FILLER_118_802 ();
 FILLCELL_X4 FILLER_118_810 ();
 FILLCELL_X2 FILLER_118_814 ();
 FILLCELL_X32 FILLER_118_826 ();
 FILLCELL_X32 FILLER_118_858 ();
 FILLCELL_X32 FILLER_118_890 ();
 FILLCELL_X32 FILLER_118_922 ();
 FILLCELL_X32 FILLER_118_954 ();
 FILLCELL_X32 FILLER_118_986 ();
 FILLCELL_X32 FILLER_118_1018 ();
 FILLCELL_X32 FILLER_118_1050 ();
 FILLCELL_X32 FILLER_118_1082 ();
 FILLCELL_X32 FILLER_118_1114 ();
 FILLCELL_X32 FILLER_118_1146 ();
 FILLCELL_X32 FILLER_118_1178 ();
 FILLCELL_X32 FILLER_118_1210 ();
 FILLCELL_X32 FILLER_118_1242 ();
 FILLCELL_X32 FILLER_118_1274 ();
 FILLCELL_X32 FILLER_118_1306 ();
 FILLCELL_X32 FILLER_118_1338 ();
 FILLCELL_X32 FILLER_118_1370 ();
 FILLCELL_X32 FILLER_118_1402 ();
 FILLCELL_X32 FILLER_118_1434 ();
 FILLCELL_X32 FILLER_118_1466 ();
 FILLCELL_X32 FILLER_118_1498 ();
 FILLCELL_X32 FILLER_118_1530 ();
 FILLCELL_X4 FILLER_118_1562 ();
 FILLCELL_X1 FILLER_118_1566 ();
 FILLCELL_X16 FILLER_118_1581 ();
 FILLCELL_X2 FILLER_118_1597 ();
 FILLCELL_X1 FILLER_118_1599 ();
 FILLCELL_X1 FILLER_118_1613 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X16 FILLER_119_769 ();
 FILLCELL_X4 FILLER_119_785 ();
 FILLCELL_X8 FILLER_119_799 ();
 FILLCELL_X2 FILLER_119_807 ();
 FILLCELL_X32 FILLER_119_813 ();
 FILLCELL_X32 FILLER_119_845 ();
 FILLCELL_X32 FILLER_119_877 ();
 FILLCELL_X32 FILLER_119_909 ();
 FILLCELL_X32 FILLER_119_941 ();
 FILLCELL_X32 FILLER_119_973 ();
 FILLCELL_X32 FILLER_119_1005 ();
 FILLCELL_X32 FILLER_119_1037 ();
 FILLCELL_X32 FILLER_119_1069 ();
 FILLCELL_X32 FILLER_119_1101 ();
 FILLCELL_X32 FILLER_119_1133 ();
 FILLCELL_X32 FILLER_119_1165 ();
 FILLCELL_X32 FILLER_119_1197 ();
 FILLCELL_X32 FILLER_119_1229 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X8 FILLER_119_1552 ();
 FILLCELL_X4 FILLER_119_1560 ();
 FILLCELL_X2 FILLER_119_1564 ();
 FILLCELL_X1 FILLER_119_1566 ();
 FILLCELL_X1 FILLER_119_1580 ();
 FILLCELL_X16 FILLER_119_1589 ();
 FILLCELL_X4 FILLER_119_1608 ();
 FILLCELL_X2 FILLER_119_1612 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X8 FILLER_120_792 ();
 FILLCELL_X2 FILLER_120_800 ();
 FILLCELL_X32 FILLER_120_807 ();
 FILLCELL_X32 FILLER_120_839 ();
 FILLCELL_X32 FILLER_120_871 ();
 FILLCELL_X32 FILLER_120_903 ();
 FILLCELL_X32 FILLER_120_935 ();
 FILLCELL_X32 FILLER_120_967 ();
 FILLCELL_X32 FILLER_120_999 ();
 FILLCELL_X32 FILLER_120_1031 ();
 FILLCELL_X32 FILLER_120_1063 ();
 FILLCELL_X32 FILLER_120_1095 ();
 FILLCELL_X32 FILLER_120_1127 ();
 FILLCELL_X32 FILLER_120_1159 ();
 FILLCELL_X32 FILLER_120_1191 ();
 FILLCELL_X32 FILLER_120_1223 ();
 FILLCELL_X32 FILLER_120_1255 ();
 FILLCELL_X32 FILLER_120_1287 ();
 FILLCELL_X32 FILLER_120_1319 ();
 FILLCELL_X32 FILLER_120_1351 ();
 FILLCELL_X32 FILLER_120_1383 ();
 FILLCELL_X32 FILLER_120_1415 ();
 FILLCELL_X32 FILLER_120_1447 ();
 FILLCELL_X32 FILLER_120_1479 ();
 FILLCELL_X32 FILLER_120_1511 ();
 FILLCELL_X32 FILLER_120_1543 ();
 FILLCELL_X8 FILLER_120_1575 ();
 FILLCELL_X4 FILLER_120_1583 ();
 FILLCELL_X2 FILLER_120_1587 ();
 FILLCELL_X1 FILLER_120_1589 ();
 FILLCELL_X4 FILLER_120_1595 ();
 FILLCELL_X2 FILLER_120_1599 ();
 FILLCELL_X4 FILLER_120_1604 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X1 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_812 ();
 FILLCELL_X32 FILLER_121_844 ();
 FILLCELL_X32 FILLER_121_876 ();
 FILLCELL_X32 FILLER_121_908 ();
 FILLCELL_X32 FILLER_121_940 ();
 FILLCELL_X32 FILLER_121_972 ();
 FILLCELL_X32 FILLER_121_1004 ();
 FILLCELL_X32 FILLER_121_1036 ();
 FILLCELL_X32 FILLER_121_1068 ();
 FILLCELL_X32 FILLER_121_1100 ();
 FILLCELL_X32 FILLER_121_1132 ();
 FILLCELL_X32 FILLER_121_1164 ();
 FILLCELL_X32 FILLER_121_1196 ();
 FILLCELL_X32 FILLER_121_1228 ();
 FILLCELL_X2 FILLER_121_1260 ();
 FILLCELL_X1 FILLER_121_1262 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X16 FILLER_121_1552 ();
 FILLCELL_X8 FILLER_121_1568 ();
 FILLCELL_X4 FILLER_121_1576 ();
 FILLCELL_X1 FILLER_121_1584 ();
 FILLCELL_X2 FILLER_121_1611 ();
 FILLCELL_X1 FILLER_121_1613 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X32 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_122_1240 ();
 FILLCELL_X32 FILLER_122_1272 ();
 FILLCELL_X32 FILLER_122_1304 ();
 FILLCELL_X32 FILLER_122_1336 ();
 FILLCELL_X32 FILLER_122_1368 ();
 FILLCELL_X32 FILLER_122_1400 ();
 FILLCELL_X32 FILLER_122_1432 ();
 FILLCELL_X32 FILLER_122_1464 ();
 FILLCELL_X32 FILLER_122_1496 ();
 FILLCELL_X32 FILLER_122_1528 ();
 FILLCELL_X16 FILLER_122_1560 ();
 FILLCELL_X8 FILLER_122_1578 ();
 FILLCELL_X4 FILLER_122_1586 ();
 FILLCELL_X1 FILLER_122_1590 ();
 FILLCELL_X2 FILLER_122_1599 ();
 FILLCELL_X1 FILLER_122_1601 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X32 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1121 ();
 FILLCELL_X32 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X32 FILLER_123_1217 ();
 FILLCELL_X8 FILLER_123_1249 ();
 FILLCELL_X4 FILLER_123_1257 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X16 FILLER_123_1552 ();
 FILLCELL_X8 FILLER_123_1568 ();
 FILLCELL_X4 FILLER_123_1586 ();
 FILLCELL_X2 FILLER_123_1596 ();
 FILLCELL_X4 FILLER_123_1601 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X16 FILLER_124_1592 ();
 FILLCELL_X4 FILLER_124_1608 ();
 FILLCELL_X2 FILLER_124_1612 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X32 FILLER_125_1089 ();
 FILLCELL_X32 FILLER_125_1121 ();
 FILLCELL_X32 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1185 ();
 FILLCELL_X32 FILLER_125_1217 ();
 FILLCELL_X8 FILLER_125_1249 ();
 FILLCELL_X4 FILLER_125_1257 ();
 FILLCELL_X2 FILLER_125_1261 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X16 FILLER_125_1584 ();
 FILLCELL_X8 FILLER_125_1600 ();
 FILLCELL_X4 FILLER_125_1608 ();
 FILLCELL_X2 FILLER_125_1612 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X32 FILLER_126_1112 ();
 FILLCELL_X32 FILLER_126_1144 ();
 FILLCELL_X32 FILLER_126_1176 ();
 FILLCELL_X32 FILLER_126_1208 ();
 FILLCELL_X32 FILLER_126_1240 ();
 FILLCELL_X32 FILLER_126_1272 ();
 FILLCELL_X32 FILLER_126_1304 ();
 FILLCELL_X32 FILLER_126_1336 ();
 FILLCELL_X32 FILLER_126_1368 ();
 FILLCELL_X32 FILLER_126_1400 ();
 FILLCELL_X32 FILLER_126_1432 ();
 FILLCELL_X32 FILLER_126_1464 ();
 FILLCELL_X32 FILLER_126_1496 ();
 FILLCELL_X32 FILLER_126_1528 ();
 FILLCELL_X32 FILLER_126_1560 ();
 FILLCELL_X16 FILLER_126_1592 ();
 FILLCELL_X4 FILLER_126_1608 ();
 FILLCELL_X2 FILLER_126_1612 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X16 FILLER_127_1584 ();
 FILLCELL_X8 FILLER_127_1600 ();
 FILLCELL_X4 FILLER_127_1608 ();
 FILLCELL_X2 FILLER_127_1612 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X32 FILLER_128_1112 ();
 FILLCELL_X32 FILLER_128_1144 ();
 FILLCELL_X32 FILLER_128_1176 ();
 FILLCELL_X32 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_128_1240 ();
 FILLCELL_X32 FILLER_128_1272 ();
 FILLCELL_X32 FILLER_128_1304 ();
 FILLCELL_X32 FILLER_128_1336 ();
 FILLCELL_X32 FILLER_128_1368 ();
 FILLCELL_X32 FILLER_128_1400 ();
 FILLCELL_X32 FILLER_128_1432 ();
 FILLCELL_X32 FILLER_128_1464 ();
 FILLCELL_X32 FILLER_128_1496 ();
 FILLCELL_X32 FILLER_128_1528 ();
 FILLCELL_X32 FILLER_128_1560 ();
 FILLCELL_X16 FILLER_128_1592 ();
 FILLCELL_X4 FILLER_128_1608 ();
 FILLCELL_X2 FILLER_128_1612 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X32 FILLER_129_1089 ();
 FILLCELL_X32 FILLER_129_1121 ();
 FILLCELL_X32 FILLER_129_1153 ();
 FILLCELL_X32 FILLER_129_1185 ();
 FILLCELL_X32 FILLER_129_1217 ();
 FILLCELL_X8 FILLER_129_1249 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X16 FILLER_129_1584 ();
 FILLCELL_X8 FILLER_129_1600 ();
 FILLCELL_X4 FILLER_129_1608 ();
 FILLCELL_X2 FILLER_129_1612 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X32 FILLER_130_1080 ();
 FILLCELL_X32 FILLER_130_1112 ();
 FILLCELL_X32 FILLER_130_1144 ();
 FILLCELL_X32 FILLER_130_1176 ();
 FILLCELL_X32 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_130_1240 ();
 FILLCELL_X32 FILLER_130_1272 ();
 FILLCELL_X32 FILLER_130_1304 ();
 FILLCELL_X32 FILLER_130_1336 ();
 FILLCELL_X32 FILLER_130_1368 ();
 FILLCELL_X32 FILLER_130_1400 ();
 FILLCELL_X32 FILLER_130_1432 ();
 FILLCELL_X32 FILLER_130_1464 ();
 FILLCELL_X32 FILLER_130_1496 ();
 FILLCELL_X32 FILLER_130_1528 ();
 FILLCELL_X32 FILLER_130_1560 ();
 FILLCELL_X16 FILLER_130_1592 ();
 FILLCELL_X4 FILLER_130_1608 ();
 FILLCELL_X2 FILLER_130_1612 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X32 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_1025 ();
 FILLCELL_X32 FILLER_131_1057 ();
 FILLCELL_X32 FILLER_131_1089 ();
 FILLCELL_X32 FILLER_131_1121 ();
 FILLCELL_X32 FILLER_131_1153 ();
 FILLCELL_X32 FILLER_131_1185 ();
 FILLCELL_X32 FILLER_131_1217 ();
 FILLCELL_X8 FILLER_131_1249 ();
 FILLCELL_X4 FILLER_131_1257 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X16 FILLER_131_1584 ();
 FILLCELL_X8 FILLER_131_1600 ();
 FILLCELL_X4 FILLER_131_1608 ();
 FILLCELL_X2 FILLER_131_1612 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X32 FILLER_132_1080 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X32 FILLER_132_1144 ();
 FILLCELL_X32 FILLER_132_1176 ();
 FILLCELL_X32 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_132_1240 ();
 FILLCELL_X32 FILLER_132_1272 ();
 FILLCELL_X32 FILLER_132_1304 ();
 FILLCELL_X32 FILLER_132_1336 ();
 FILLCELL_X32 FILLER_132_1368 ();
 FILLCELL_X32 FILLER_132_1400 ();
 FILLCELL_X32 FILLER_132_1432 ();
 FILLCELL_X32 FILLER_132_1464 ();
 FILLCELL_X32 FILLER_132_1496 ();
 FILLCELL_X32 FILLER_132_1528 ();
 FILLCELL_X32 FILLER_132_1560 ();
 FILLCELL_X16 FILLER_132_1592 ();
 FILLCELL_X4 FILLER_132_1608 ();
 FILLCELL_X2 FILLER_132_1612 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X32 FILLER_133_1121 ();
 FILLCELL_X32 FILLER_133_1153 ();
 FILLCELL_X32 FILLER_133_1185 ();
 FILLCELL_X32 FILLER_133_1217 ();
 FILLCELL_X8 FILLER_133_1249 ();
 FILLCELL_X4 FILLER_133_1257 ();
 FILLCELL_X2 FILLER_133_1261 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X16 FILLER_133_1584 ();
 FILLCELL_X8 FILLER_133_1600 ();
 FILLCELL_X4 FILLER_133_1608 ();
 FILLCELL_X2 FILLER_133_1612 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_134_1048 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X16 FILLER_134_1592 ();
 FILLCELL_X4 FILLER_134_1608 ();
 FILLCELL_X2 FILLER_134_1612 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X32 FILLER_135_993 ();
 FILLCELL_X32 FILLER_135_1025 ();
 FILLCELL_X32 FILLER_135_1057 ();
 FILLCELL_X32 FILLER_135_1089 ();
 FILLCELL_X32 FILLER_135_1121 ();
 FILLCELL_X32 FILLER_135_1153 ();
 FILLCELL_X32 FILLER_135_1185 ();
 FILLCELL_X32 FILLER_135_1217 ();
 FILLCELL_X8 FILLER_135_1249 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X16 FILLER_135_1584 ();
 FILLCELL_X8 FILLER_135_1600 ();
 FILLCELL_X4 FILLER_135_1608 ();
 FILLCELL_X2 FILLER_135_1612 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X32 FILLER_136_1016 ();
 FILLCELL_X32 FILLER_136_1048 ();
 FILLCELL_X32 FILLER_136_1080 ();
 FILLCELL_X32 FILLER_136_1112 ();
 FILLCELL_X32 FILLER_136_1144 ();
 FILLCELL_X32 FILLER_136_1176 ();
 FILLCELL_X32 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_136_1240 ();
 FILLCELL_X32 FILLER_136_1272 ();
 FILLCELL_X32 FILLER_136_1304 ();
 FILLCELL_X32 FILLER_136_1336 ();
 FILLCELL_X32 FILLER_136_1368 ();
 FILLCELL_X32 FILLER_136_1400 ();
 FILLCELL_X32 FILLER_136_1432 ();
 FILLCELL_X32 FILLER_136_1464 ();
 FILLCELL_X32 FILLER_136_1496 ();
 FILLCELL_X32 FILLER_136_1528 ();
 FILLCELL_X32 FILLER_136_1560 ();
 FILLCELL_X16 FILLER_136_1592 ();
 FILLCELL_X4 FILLER_136_1608 ();
 FILLCELL_X2 FILLER_136_1612 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X32 FILLER_137_961 ();
 FILLCELL_X32 FILLER_137_993 ();
 FILLCELL_X32 FILLER_137_1025 ();
 FILLCELL_X32 FILLER_137_1057 ();
 FILLCELL_X32 FILLER_137_1089 ();
 FILLCELL_X32 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1153 ();
 FILLCELL_X32 FILLER_137_1185 ();
 FILLCELL_X32 FILLER_137_1217 ();
 FILLCELL_X8 FILLER_137_1249 ();
 FILLCELL_X4 FILLER_137_1257 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X16 FILLER_137_1584 ();
 FILLCELL_X8 FILLER_137_1600 ();
 FILLCELL_X4 FILLER_137_1608 ();
 FILLCELL_X2 FILLER_137_1612 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X32 FILLER_138_984 ();
 FILLCELL_X32 FILLER_138_1016 ();
 FILLCELL_X32 FILLER_138_1048 ();
 FILLCELL_X32 FILLER_138_1080 ();
 FILLCELL_X32 FILLER_138_1112 ();
 FILLCELL_X32 FILLER_138_1144 ();
 FILLCELL_X32 FILLER_138_1176 ();
 FILLCELL_X32 FILLER_138_1208 ();
 FILLCELL_X32 FILLER_138_1240 ();
 FILLCELL_X32 FILLER_138_1272 ();
 FILLCELL_X32 FILLER_138_1304 ();
 FILLCELL_X32 FILLER_138_1336 ();
 FILLCELL_X32 FILLER_138_1368 ();
 FILLCELL_X32 FILLER_138_1400 ();
 FILLCELL_X32 FILLER_138_1432 ();
 FILLCELL_X32 FILLER_138_1464 ();
 FILLCELL_X32 FILLER_138_1496 ();
 FILLCELL_X32 FILLER_138_1528 ();
 FILLCELL_X32 FILLER_138_1560 ();
 FILLCELL_X16 FILLER_138_1592 ();
 FILLCELL_X4 FILLER_138_1608 ();
 FILLCELL_X2 FILLER_138_1612 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X32 FILLER_139_1057 ();
 FILLCELL_X32 FILLER_139_1089 ();
 FILLCELL_X32 FILLER_139_1121 ();
 FILLCELL_X32 FILLER_139_1153 ();
 FILLCELL_X32 FILLER_139_1185 ();
 FILLCELL_X32 FILLER_139_1217 ();
 FILLCELL_X8 FILLER_139_1249 ();
 FILLCELL_X4 FILLER_139_1257 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X16 FILLER_139_1584 ();
 FILLCELL_X8 FILLER_139_1600 ();
 FILLCELL_X4 FILLER_139_1608 ();
 FILLCELL_X2 FILLER_139_1612 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X16 FILLER_140_1592 ();
 FILLCELL_X4 FILLER_140_1608 ();
 FILLCELL_X2 FILLER_140_1612 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X32 FILLER_141_1121 ();
 FILLCELL_X32 FILLER_141_1153 ();
 FILLCELL_X32 FILLER_141_1185 ();
 FILLCELL_X32 FILLER_141_1217 ();
 FILLCELL_X8 FILLER_141_1249 ();
 FILLCELL_X4 FILLER_141_1257 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X16 FILLER_141_1584 ();
 FILLCELL_X8 FILLER_141_1600 ();
 FILLCELL_X4 FILLER_141_1608 ();
 FILLCELL_X2 FILLER_141_1612 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X16 FILLER_142_1592 ();
 FILLCELL_X4 FILLER_142_1608 ();
 FILLCELL_X2 FILLER_142_1612 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X16 FILLER_143_1584 ();
 FILLCELL_X8 FILLER_143_1600 ();
 FILLCELL_X4 FILLER_143_1608 ();
 FILLCELL_X2 FILLER_143_1612 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X16 FILLER_144_1592 ();
 FILLCELL_X4 FILLER_144_1608 ();
 FILLCELL_X2 FILLER_144_1612 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X16 FILLER_145_1584 ();
 FILLCELL_X8 FILLER_145_1600 ();
 FILLCELL_X4 FILLER_145_1608 ();
 FILLCELL_X2 FILLER_145_1612 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X16 FILLER_146_1592 ();
 FILLCELL_X4 FILLER_146_1608 ();
 FILLCELL_X2 FILLER_146_1612 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X16 FILLER_147_1584 ();
 FILLCELL_X8 FILLER_147_1600 ();
 FILLCELL_X4 FILLER_147_1608 ();
 FILLCELL_X2 FILLER_147_1612 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X16 FILLER_148_1592 ();
 FILLCELL_X4 FILLER_148_1608 ();
 FILLCELL_X2 FILLER_148_1612 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X16 FILLER_149_1584 ();
 FILLCELL_X8 FILLER_149_1600 ();
 FILLCELL_X4 FILLER_149_1608 ();
 FILLCELL_X2 FILLER_149_1612 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X16 FILLER_150_1592 ();
 FILLCELL_X4 FILLER_150_1608 ();
 FILLCELL_X2 FILLER_150_1612 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X16 FILLER_151_1584 ();
 FILLCELL_X8 FILLER_151_1600 ();
 FILLCELL_X4 FILLER_151_1608 ();
 FILLCELL_X2 FILLER_151_1612 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X16 FILLER_152_1592 ();
 FILLCELL_X4 FILLER_152_1608 ();
 FILLCELL_X2 FILLER_152_1612 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X16 FILLER_153_1584 ();
 FILLCELL_X8 FILLER_153_1600 ();
 FILLCELL_X4 FILLER_153_1608 ();
 FILLCELL_X2 FILLER_153_1612 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X16 FILLER_154_1592 ();
 FILLCELL_X4 FILLER_154_1608 ();
 FILLCELL_X2 FILLER_154_1612 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X16 FILLER_155_1584 ();
 FILLCELL_X8 FILLER_155_1600 ();
 FILLCELL_X4 FILLER_155_1608 ();
 FILLCELL_X2 FILLER_155_1612 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X16 FILLER_156_1592 ();
 FILLCELL_X4 FILLER_156_1608 ();
 FILLCELL_X2 FILLER_156_1612 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X16 FILLER_157_1584 ();
 FILLCELL_X8 FILLER_157_1600 ();
 FILLCELL_X4 FILLER_157_1608 ();
 FILLCELL_X2 FILLER_157_1612 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X16 FILLER_158_1592 ();
 FILLCELL_X4 FILLER_158_1608 ();
 FILLCELL_X2 FILLER_158_1612 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X16 FILLER_159_1584 ();
 FILLCELL_X8 FILLER_159_1600 ();
 FILLCELL_X4 FILLER_159_1608 ();
 FILLCELL_X2 FILLER_159_1612 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X16 FILLER_160_1592 ();
 FILLCELL_X4 FILLER_160_1608 ();
 FILLCELL_X2 FILLER_160_1612 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X16 FILLER_161_1584 ();
 FILLCELL_X8 FILLER_161_1600 ();
 FILLCELL_X4 FILLER_161_1608 ();
 FILLCELL_X2 FILLER_161_1612 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1304 ();
 FILLCELL_X32 FILLER_162_1336 ();
 FILLCELL_X32 FILLER_162_1368 ();
 FILLCELL_X32 FILLER_162_1400 ();
 FILLCELL_X32 FILLER_162_1432 ();
 FILLCELL_X32 FILLER_162_1464 ();
 FILLCELL_X32 FILLER_162_1496 ();
 FILLCELL_X32 FILLER_162_1528 ();
 FILLCELL_X32 FILLER_162_1560 ();
 FILLCELL_X16 FILLER_162_1592 ();
 FILLCELL_X4 FILLER_162_1608 ();
 FILLCELL_X2 FILLER_162_1612 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X16 FILLER_163_1584 ();
 FILLCELL_X8 FILLER_163_1600 ();
 FILLCELL_X4 FILLER_163_1608 ();
 FILLCELL_X2 FILLER_163_1612 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X32 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1336 ();
 FILLCELL_X32 FILLER_164_1368 ();
 FILLCELL_X32 FILLER_164_1400 ();
 FILLCELL_X32 FILLER_164_1432 ();
 FILLCELL_X32 FILLER_164_1464 ();
 FILLCELL_X32 FILLER_164_1496 ();
 FILLCELL_X32 FILLER_164_1528 ();
 FILLCELL_X32 FILLER_164_1560 ();
 FILLCELL_X16 FILLER_164_1592 ();
 FILLCELL_X4 FILLER_164_1608 ();
 FILLCELL_X2 FILLER_164_1612 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X16 FILLER_165_1584 ();
 FILLCELL_X8 FILLER_165_1600 ();
 FILLCELL_X4 FILLER_165_1608 ();
 FILLCELL_X2 FILLER_165_1612 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X32 FILLER_166_1112 ();
 FILLCELL_X32 FILLER_166_1144 ();
 FILLCELL_X32 FILLER_166_1176 ();
 FILLCELL_X32 FILLER_166_1208 ();
 FILLCELL_X32 FILLER_166_1240 ();
 FILLCELL_X32 FILLER_166_1272 ();
 FILLCELL_X32 FILLER_166_1304 ();
 FILLCELL_X32 FILLER_166_1336 ();
 FILLCELL_X32 FILLER_166_1368 ();
 FILLCELL_X32 FILLER_166_1400 ();
 FILLCELL_X32 FILLER_166_1432 ();
 FILLCELL_X32 FILLER_166_1464 ();
 FILLCELL_X32 FILLER_166_1496 ();
 FILLCELL_X32 FILLER_166_1528 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X16 FILLER_166_1592 ();
 FILLCELL_X4 FILLER_166_1608 ();
 FILLCELL_X2 FILLER_166_1612 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X16 FILLER_167_1584 ();
 FILLCELL_X8 FILLER_167_1600 ();
 FILLCELL_X4 FILLER_167_1608 ();
 FILLCELL_X2 FILLER_167_1612 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X32 FILLER_168_1304 ();
 FILLCELL_X32 FILLER_168_1336 ();
 FILLCELL_X32 FILLER_168_1368 ();
 FILLCELL_X32 FILLER_168_1400 ();
 FILLCELL_X32 FILLER_168_1432 ();
 FILLCELL_X32 FILLER_168_1464 ();
 FILLCELL_X32 FILLER_168_1496 ();
 FILLCELL_X32 FILLER_168_1528 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X16 FILLER_168_1592 ();
 FILLCELL_X4 FILLER_168_1608 ();
 FILLCELL_X2 FILLER_168_1612 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X32 FILLER_169_1089 ();
 FILLCELL_X32 FILLER_169_1121 ();
 FILLCELL_X32 FILLER_169_1153 ();
 FILLCELL_X32 FILLER_169_1185 ();
 FILLCELL_X32 FILLER_169_1217 ();
 FILLCELL_X8 FILLER_169_1249 ();
 FILLCELL_X4 FILLER_169_1257 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X16 FILLER_169_1584 ();
 FILLCELL_X8 FILLER_169_1600 ();
 FILLCELL_X4 FILLER_169_1608 ();
 FILLCELL_X2 FILLER_169_1612 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X32 FILLER_170_1080 ();
 FILLCELL_X32 FILLER_170_1112 ();
 FILLCELL_X32 FILLER_170_1144 ();
 FILLCELL_X32 FILLER_170_1176 ();
 FILLCELL_X32 FILLER_170_1208 ();
 FILLCELL_X32 FILLER_170_1240 ();
 FILLCELL_X32 FILLER_170_1272 ();
 FILLCELL_X32 FILLER_170_1304 ();
 FILLCELL_X32 FILLER_170_1336 ();
 FILLCELL_X32 FILLER_170_1368 ();
 FILLCELL_X32 FILLER_170_1400 ();
 FILLCELL_X32 FILLER_170_1432 ();
 FILLCELL_X32 FILLER_170_1464 ();
 FILLCELL_X32 FILLER_170_1496 ();
 FILLCELL_X32 FILLER_170_1528 ();
 FILLCELL_X32 FILLER_170_1560 ();
 FILLCELL_X16 FILLER_170_1592 ();
 FILLCELL_X4 FILLER_170_1608 ();
 FILLCELL_X2 FILLER_170_1612 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X32 FILLER_171_1185 ();
 FILLCELL_X32 FILLER_171_1217 ();
 FILLCELL_X8 FILLER_171_1249 ();
 FILLCELL_X4 FILLER_171_1257 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X16 FILLER_171_1584 ();
 FILLCELL_X8 FILLER_171_1600 ();
 FILLCELL_X4 FILLER_171_1608 ();
 FILLCELL_X2 FILLER_171_1612 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X32 FILLER_172_1080 ();
 FILLCELL_X32 FILLER_172_1112 ();
 FILLCELL_X32 FILLER_172_1144 ();
 FILLCELL_X32 FILLER_172_1176 ();
 FILLCELL_X32 FILLER_172_1208 ();
 FILLCELL_X32 FILLER_172_1240 ();
 FILLCELL_X32 FILLER_172_1272 ();
 FILLCELL_X32 FILLER_172_1304 ();
 FILLCELL_X32 FILLER_172_1336 ();
 FILLCELL_X32 FILLER_172_1368 ();
 FILLCELL_X32 FILLER_172_1400 ();
 FILLCELL_X32 FILLER_172_1432 ();
 FILLCELL_X32 FILLER_172_1464 ();
 FILLCELL_X32 FILLER_172_1496 ();
 FILLCELL_X32 FILLER_172_1528 ();
 FILLCELL_X32 FILLER_172_1560 ();
 FILLCELL_X16 FILLER_172_1592 ();
 FILLCELL_X4 FILLER_172_1608 ();
 FILLCELL_X2 FILLER_172_1612 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X16 FILLER_173_1584 ();
 FILLCELL_X8 FILLER_173_1600 ();
 FILLCELL_X4 FILLER_173_1608 ();
 FILLCELL_X2 FILLER_173_1612 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X16 FILLER_174_1592 ();
 FILLCELL_X4 FILLER_174_1608 ();
 FILLCELL_X2 FILLER_174_1612 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X16 FILLER_175_1584 ();
 FILLCELL_X8 FILLER_175_1600 ();
 FILLCELL_X4 FILLER_175_1608 ();
 FILLCELL_X2 FILLER_175_1612 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X32 FILLER_176_1304 ();
 FILLCELL_X32 FILLER_176_1336 ();
 FILLCELL_X32 FILLER_176_1368 ();
 FILLCELL_X32 FILLER_176_1400 ();
 FILLCELL_X32 FILLER_176_1432 ();
 FILLCELL_X32 FILLER_176_1464 ();
 FILLCELL_X32 FILLER_176_1496 ();
 FILLCELL_X32 FILLER_176_1528 ();
 FILLCELL_X32 FILLER_176_1560 ();
 FILLCELL_X16 FILLER_176_1592 ();
 FILLCELL_X4 FILLER_176_1608 ();
 FILLCELL_X2 FILLER_176_1612 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X32 FILLER_177_1121 ();
 FILLCELL_X32 FILLER_177_1153 ();
 FILLCELL_X32 FILLER_177_1185 ();
 FILLCELL_X32 FILLER_177_1217 ();
 FILLCELL_X8 FILLER_177_1249 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X16 FILLER_177_1584 ();
 FILLCELL_X8 FILLER_177_1600 ();
 FILLCELL_X4 FILLER_177_1608 ();
 FILLCELL_X2 FILLER_177_1612 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X16 FILLER_178_1592 ();
 FILLCELL_X4 FILLER_178_1608 ();
 FILLCELL_X2 FILLER_178_1612 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X16 FILLER_179_1584 ();
 FILLCELL_X8 FILLER_179_1600 ();
 FILLCELL_X4 FILLER_179_1608 ();
 FILLCELL_X2 FILLER_179_1612 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X16 FILLER_180_1592 ();
 FILLCELL_X4 FILLER_180_1608 ();
 FILLCELL_X2 FILLER_180_1612 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X16 FILLER_181_1584 ();
 FILLCELL_X8 FILLER_181_1600 ();
 FILLCELL_X4 FILLER_181_1608 ();
 FILLCELL_X2 FILLER_181_1612 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X16 FILLER_182_1592 ();
 FILLCELL_X4 FILLER_182_1608 ();
 FILLCELL_X2 FILLER_182_1612 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X16 FILLER_183_1584 ();
 FILLCELL_X8 FILLER_183_1600 ();
 FILLCELL_X4 FILLER_183_1608 ();
 FILLCELL_X2 FILLER_183_1612 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X16 FILLER_184_1592 ();
 FILLCELL_X4 FILLER_184_1608 ();
 FILLCELL_X2 FILLER_184_1612 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X16 FILLER_185_1584 ();
 FILLCELL_X8 FILLER_185_1600 ();
 FILLCELL_X4 FILLER_185_1608 ();
 FILLCELL_X2 FILLER_185_1612 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X16 FILLER_186_1592 ();
 FILLCELL_X4 FILLER_186_1608 ();
 FILLCELL_X2 FILLER_186_1612 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X16 FILLER_187_1584 ();
 FILLCELL_X8 FILLER_187_1600 ();
 FILLCELL_X4 FILLER_187_1608 ();
 FILLCELL_X2 FILLER_187_1612 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X16 FILLER_188_1592 ();
 FILLCELL_X4 FILLER_188_1608 ();
 FILLCELL_X2 FILLER_188_1612 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X16 FILLER_189_1584 ();
 FILLCELL_X8 FILLER_189_1600 ();
 FILLCELL_X4 FILLER_189_1608 ();
 FILLCELL_X2 FILLER_189_1612 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X16 FILLER_190_1592 ();
 FILLCELL_X4 FILLER_190_1608 ();
 FILLCELL_X2 FILLER_190_1612 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X16 FILLER_191_1584 ();
 FILLCELL_X8 FILLER_191_1600 ();
 FILLCELL_X4 FILLER_191_1608 ();
 FILLCELL_X2 FILLER_191_1612 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X16 FILLER_192_1592 ();
 FILLCELL_X4 FILLER_192_1608 ();
 FILLCELL_X2 FILLER_192_1612 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X16 FILLER_193_1584 ();
 FILLCELL_X8 FILLER_193_1600 ();
 FILLCELL_X4 FILLER_193_1608 ();
 FILLCELL_X2 FILLER_193_1612 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X16 FILLER_194_1592 ();
 FILLCELL_X4 FILLER_194_1608 ();
 FILLCELL_X2 FILLER_194_1612 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X16 FILLER_195_1584 ();
 FILLCELL_X8 FILLER_195_1600 ();
 FILLCELL_X4 FILLER_195_1608 ();
 FILLCELL_X2 FILLER_195_1612 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X16 FILLER_196_1592 ();
 FILLCELL_X4 FILLER_196_1608 ();
 FILLCELL_X2 FILLER_196_1612 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X16 FILLER_197_1584 ();
 FILLCELL_X8 FILLER_197_1600 ();
 FILLCELL_X4 FILLER_197_1608 ();
 FILLCELL_X2 FILLER_197_1612 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X16 FILLER_198_1592 ();
 FILLCELL_X4 FILLER_198_1608 ();
 FILLCELL_X2 FILLER_198_1612 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X16 FILLER_199_1584 ();
 FILLCELL_X8 FILLER_199_1600 ();
 FILLCELL_X4 FILLER_199_1608 ();
 FILLCELL_X2 FILLER_199_1612 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X16 FILLER_200_1592 ();
 FILLCELL_X4 FILLER_200_1608 ();
 FILLCELL_X2 FILLER_200_1612 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X16 FILLER_201_1584 ();
 FILLCELL_X8 FILLER_201_1600 ();
 FILLCELL_X4 FILLER_201_1608 ();
 FILLCELL_X2 FILLER_201_1612 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X16 FILLER_202_1592 ();
 FILLCELL_X4 FILLER_202_1608 ();
 FILLCELL_X2 FILLER_202_1612 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X16 FILLER_203_1584 ();
 FILLCELL_X8 FILLER_203_1600 ();
 FILLCELL_X4 FILLER_203_1608 ();
 FILLCELL_X2 FILLER_203_1612 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X16 FILLER_204_1592 ();
 FILLCELL_X4 FILLER_204_1608 ();
 FILLCELL_X2 FILLER_204_1612 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X16 FILLER_205_1584 ();
 FILLCELL_X8 FILLER_205_1600 ();
 FILLCELL_X4 FILLER_205_1608 ();
 FILLCELL_X2 FILLER_205_1612 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X16 FILLER_206_1592 ();
 FILLCELL_X4 FILLER_206_1608 ();
 FILLCELL_X2 FILLER_206_1612 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X16 FILLER_207_1584 ();
 FILLCELL_X8 FILLER_207_1600 ();
 FILLCELL_X4 FILLER_207_1608 ();
 FILLCELL_X2 FILLER_207_1612 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X16 FILLER_208_1592 ();
 FILLCELL_X4 FILLER_208_1608 ();
 FILLCELL_X2 FILLER_208_1612 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X16 FILLER_209_1584 ();
 FILLCELL_X8 FILLER_209_1600 ();
 FILLCELL_X4 FILLER_209_1608 ();
 FILLCELL_X2 FILLER_209_1612 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X16 FILLER_210_1592 ();
 FILLCELL_X4 FILLER_210_1608 ();
 FILLCELL_X2 FILLER_210_1612 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X16 FILLER_211_1584 ();
 FILLCELL_X8 FILLER_211_1600 ();
 FILLCELL_X4 FILLER_211_1608 ();
 FILLCELL_X2 FILLER_211_1612 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X16 FILLER_212_1592 ();
 FILLCELL_X4 FILLER_212_1608 ();
 FILLCELL_X2 FILLER_212_1612 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X16 FILLER_213_1584 ();
 FILLCELL_X8 FILLER_213_1600 ();
 FILLCELL_X4 FILLER_213_1608 ();
 FILLCELL_X2 FILLER_213_1612 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X16 FILLER_214_1592 ();
 FILLCELL_X4 FILLER_214_1608 ();
 FILLCELL_X2 FILLER_214_1612 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X16 FILLER_215_1584 ();
 FILLCELL_X8 FILLER_215_1600 ();
 FILLCELL_X4 FILLER_215_1608 ();
 FILLCELL_X2 FILLER_215_1612 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X16 FILLER_216_1592 ();
 FILLCELL_X4 FILLER_216_1608 ();
 FILLCELL_X2 FILLER_216_1612 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X16 FILLER_217_769 ();
 FILLCELL_X2 FILLER_217_785 ();
 FILLCELL_X1 FILLER_217_787 ();
 FILLCELL_X8 FILLER_217_792 ();
 FILLCELL_X2 FILLER_217_800 ();
 FILLCELL_X1 FILLER_217_802 ();
 FILLCELL_X32 FILLER_217_807 ();
 FILLCELL_X32 FILLER_217_839 ();
 FILLCELL_X32 FILLER_217_871 ();
 FILLCELL_X32 FILLER_217_903 ();
 FILLCELL_X32 FILLER_217_935 ();
 FILLCELL_X32 FILLER_217_967 ();
 FILLCELL_X32 FILLER_217_999 ();
 FILLCELL_X32 FILLER_217_1031 ();
 FILLCELL_X32 FILLER_217_1063 ();
 FILLCELL_X32 FILLER_217_1095 ();
 FILLCELL_X32 FILLER_217_1127 ();
 FILLCELL_X32 FILLER_217_1159 ();
 FILLCELL_X32 FILLER_217_1191 ();
 FILLCELL_X32 FILLER_217_1223 ();
 FILLCELL_X8 FILLER_217_1255 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X16 FILLER_217_1584 ();
 FILLCELL_X8 FILLER_217_1600 ();
 FILLCELL_X4 FILLER_217_1608 ();
 FILLCELL_X2 FILLER_217_1612 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X16 FILLER_218_664 ();
 FILLCELL_X4 FILLER_218_680 ();
 FILLCELL_X16 FILLER_218_692 ();
 FILLCELL_X4 FILLER_218_708 ();
 FILLCELL_X2 FILLER_218_712 ();
 FILLCELL_X4 FILLER_218_725 ();
 FILLCELL_X2 FILLER_218_729 ();
 FILLCELL_X1 FILLER_218_731 ();
 FILLCELL_X4 FILLER_218_735 ();
 FILLCELL_X2 FILLER_218_743 ();
 FILLCELL_X4 FILLER_218_749 ();
 FILLCELL_X2 FILLER_218_753 ();
 FILLCELL_X1 FILLER_218_755 ();
 FILLCELL_X8 FILLER_218_764 ();
 FILLCELL_X4 FILLER_218_772 ();
 FILLCELL_X8 FILLER_218_779 ();
 FILLCELL_X4 FILLER_218_794 ();
 FILLCELL_X1 FILLER_218_798 ();
 FILLCELL_X32 FILLER_218_806 ();
 FILLCELL_X32 FILLER_218_838 ();
 FILLCELL_X32 FILLER_218_870 ();
 FILLCELL_X32 FILLER_218_902 ();
 FILLCELL_X32 FILLER_218_934 ();
 FILLCELL_X32 FILLER_218_966 ();
 FILLCELL_X32 FILLER_218_998 ();
 FILLCELL_X32 FILLER_218_1030 ();
 FILLCELL_X32 FILLER_218_1062 ();
 FILLCELL_X32 FILLER_218_1094 ();
 FILLCELL_X32 FILLER_218_1126 ();
 FILLCELL_X32 FILLER_218_1158 ();
 FILLCELL_X32 FILLER_218_1190 ();
 FILLCELL_X32 FILLER_218_1222 ();
 FILLCELL_X8 FILLER_218_1254 ();
 FILLCELL_X32 FILLER_218_1263 ();
 FILLCELL_X32 FILLER_218_1295 ();
 FILLCELL_X32 FILLER_218_1327 ();
 FILLCELL_X32 FILLER_218_1359 ();
 FILLCELL_X32 FILLER_218_1391 ();
 FILLCELL_X32 FILLER_218_1423 ();
 FILLCELL_X32 FILLER_218_1455 ();
 FILLCELL_X32 FILLER_218_1487 ();
 FILLCELL_X32 FILLER_218_1519 ();
 FILLCELL_X32 FILLER_218_1551 ();
 FILLCELL_X16 FILLER_218_1583 ();
 FILLCELL_X8 FILLER_218_1599 ();
 FILLCELL_X4 FILLER_218_1607 ();
 FILLCELL_X2 FILLER_218_1611 ();
 FILLCELL_X1 FILLER_218_1613 ();
endmodule
