module alu (clk,
    overflow_flag,
    rst_n,
    zero_flag,
    a,
    b,
    op_code,
    result);
 input clk;
 output overflow_flag;
 input rst_n;
 output zero_flag;
 input [7:0] a;
 input [7:0] b;
 input [2:0] op_code;
 output [7:0] result;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _347_ (.A(net1),
    .ZN(_287_));
 BUF_X2 _348_ (.A(net2),
    .Z(_260_));
 INV_X1 _349_ (.A(_260_),
    .ZN(_282_));
 BUF_X4 _350_ (.A(net3),
    .Z(_261_));
 INV_X1 _351_ (.A(_261_),
    .ZN(_301_));
 BUF_X2 _352_ (.A(net4),
    .Z(_262_));
 INV_X1 _353_ (.A(_262_),
    .ZN(_309_));
 BUF_X2 _354_ (.A(net5),
    .Z(_263_));
 INV_X1 _355_ (.A(_263_),
    .ZN(_317_));
 CLKBUF_X2 _356_ (.A(net6),
    .Z(_264_));
 INV_X1 _357_ (.A(_264_),
    .ZN(_325_));
 CLKBUF_X2 _358_ (.A(net7),
    .Z(_265_));
 INV_X1 _359_ (.A(_265_),
    .ZN(_333_));
 CLKBUF_X2 _360_ (.A(net8),
    .Z(_266_));
 INV_X1 _361_ (.A(_266_),
    .ZN(_341_));
 BUF_X8 _362_ (.A(net9),
    .Z(_267_));
 BUF_X4 _363_ (.A(_267_),
    .Z(_268_));
 INV_X2 _364_ (.A(_268_),
    .ZN(_288_));
 BUF_X2 _365_ (.A(net10),
    .Z(_010_));
 INV_X2 _366_ (.A(_010_),
    .ZN(_011_));
 BUF_X4 _367_ (.A(_011_),
    .Z(_295_));
 INV_X1 _368_ (.A(net11),
    .ZN(_012_));
 BUF_X4 _369_ (.A(_012_),
    .Z(_302_));
 INV_X1 _370_ (.A(net12),
    .ZN(_310_));
 INV_X1 _371_ (.A(net13),
    .ZN(_318_));
 INV_X1 _372_ (.A(net14),
    .ZN(_326_));
 INV_X1 _373_ (.A(net15),
    .ZN(_334_));
 INV_X1 _374_ (.A(net16),
    .ZN(_342_));
 CLKBUF_X2 _375_ (.A(rst_n),
    .Z(_013_));
 BUF_X4 _376_ (.A(op_code[2]),
    .Z(_014_));
 BUF_X4 _377_ (.A(_014_),
    .Z(_015_));
 BUF_X2 _378_ (.A(op_code[1]),
    .Z(_016_));
 BUF_X4 _379_ (.A(_016_),
    .Z(_017_));
 BUF_X2 _380_ (.A(op_code[0]),
    .Z(_018_));
 BUF_X4 _381_ (.A(_018_),
    .Z(_019_));
 NOR3_X4 _382_ (.A1(_015_),
    .A2(_017_),
    .A3(_019_),
    .ZN(_020_));
 NAND2_X1 _383_ (.A1(_345_),
    .A2(_020_),
    .ZN(_021_));
 BUF_X2 _384_ (.A(_344_),
    .Z(_022_));
 CLKBUF_X3 _385_ (.A(_019_),
    .Z(_023_));
 NOR2_X1 _386_ (.A1(_014_),
    .A2(_016_),
    .ZN(_024_));
 AND2_X1 _387_ (.A1(_023_),
    .A2(_024_),
    .ZN(_025_));
 NAND2_X1 _388_ (.A1(_022_),
    .A2(_025_),
    .ZN(_026_));
 INV_X1 _389_ (.A(_337_),
    .ZN(_027_));
 CLKBUF_X3 _390_ (.A(_312_),
    .Z(_028_));
 CLKBUF_X3 _391_ (.A(_320_),
    .Z(_029_));
 BUF_X2 _392_ (.A(_336_),
    .Z(_030_));
 NOR4_X2 _393_ (.A1(_028_),
    .A2(_029_),
    .A3(_328_),
    .A4(_030_),
    .ZN(_031_));
 INV_X1 _394_ (.A(_031_),
    .ZN(_032_));
 BUF_X4 _395_ (.A(_304_),
    .Z(_033_));
 INV_X1 _396_ (.A(_033_),
    .ZN(_034_));
 NOR2_X1 _397_ (.A1(_286_),
    .A2(_283_),
    .ZN(_035_));
 OR2_X1 _398_ (.A1(_297_),
    .A2(_305_),
    .ZN(_036_));
 OAI22_X4 _399_ (.A1(_034_),
    .A2(_305_),
    .B1(_035_),
    .B2(_036_),
    .ZN(_037_));
 OAI21_X1 _400_ (.A(_027_),
    .B1(_032_),
    .B2(_037_),
    .ZN(_038_));
 INV_X1 _401_ (.A(_329_),
    .ZN(_039_));
 INV_X1 _402_ (.A(_029_),
    .ZN(_040_));
 AOI21_X1 _403_ (.A(_321_),
    .B1(_040_),
    .B2(_313_),
    .ZN(_041_));
 CLKBUF_X3 _404_ (.A(_328_),
    .Z(_042_));
 OAI21_X1 _405_ (.A(_039_),
    .B1(_041_),
    .B2(_042_),
    .ZN(_043_));
 INV_X1 _406_ (.A(_030_),
    .ZN(_044_));
 AOI21_X2 _407_ (.A(_038_),
    .B1(_043_),
    .B2(_044_),
    .ZN(_045_));
 XNOR2_X1 _408_ (.A(_341_),
    .B(_045_),
    .ZN(_046_));
 CLKBUF_X2 _409_ (.A(_339_),
    .Z(_047_));
 INV_X1 _410_ (.A(_331_),
    .ZN(_048_));
 NAND3_X1 _411_ (.A1(_280_),
    .A2(_033_),
    .A3(_028_),
    .ZN(_049_));
 CLKBUF_X2 _412_ (.A(_307_),
    .Z(_050_));
 AOI21_X1 _413_ (.A(_315_),
    .B1(_028_),
    .B2(_050_),
    .ZN(_051_));
 AOI21_X1 _414_ (.A(_040_),
    .B1(_049_),
    .B2(_051_),
    .ZN(_052_));
 OAI21_X1 _415_ (.A(_042_),
    .B1(_052_),
    .B2(_323_),
    .ZN(_053_));
 NAND2_X1 _416_ (.A1(_048_),
    .A2(_053_),
    .ZN(_054_));
 AOI21_X1 _417_ (.A(_047_),
    .B1(_054_),
    .B2(_030_),
    .ZN(_055_));
 NAND2_X1 _418_ (.A1(_022_),
    .A2(_020_),
    .ZN(_056_));
 OAI221_X1 _419_ (.A(_021_),
    .B1(_026_),
    .B2(_046_),
    .C1(_055_),
    .C2(_056_),
    .ZN(_057_));
 AND2_X1 _420_ (.A1(_013_),
    .A2(_057_),
    .ZN(_000_));
 CLKBUF_X2 _421_ (.A(_290_),
    .Z(_058_));
 NOR4_X1 _422_ (.A1(_058_),
    .A2(_033_),
    .A3(_286_),
    .A4(_022_),
    .ZN(_059_));
 NAND2_X1 _423_ (.A1(_031_),
    .A2(_059_),
    .ZN(_060_));
 CLKBUF_X3 _424_ (.A(_017_),
    .Z(_061_));
 NAND2_X1 _425_ (.A1(_061_),
    .A2(_023_),
    .ZN(_062_));
 OAI21_X1 _426_ (.A(_015_),
    .B1(_060_),
    .B2(_062_),
    .ZN(_063_));
 NOR2_X1 _427_ (.A1(_019_),
    .A2(_279_),
    .ZN(_064_));
 AOI21_X1 _428_ (.A(_064_),
    .B1(_289_),
    .B2(_023_),
    .ZN(_065_));
 MUX2_X1 _429_ (.A(_058_),
    .B(_065_),
    .S(_061_),
    .Z(_066_));
 OAI21_X1 _430_ (.A(_063_),
    .B1(_066_),
    .B2(_015_),
    .ZN(_067_));
 INV_X4 _431_ (.A(_018_),
    .ZN(_068_));
 NAND3_X2 _432_ (.A1(_014_),
    .A2(_017_),
    .A3(_068_),
    .ZN(_069_));
 CLKBUF_X3 _433_ (.A(net11),
    .Z(_070_));
 MUX2_X1 _434_ (.A(_261_),
    .B(_262_),
    .S(_268_),
    .Z(_071_));
 NOR2_X1 _435_ (.A1(_295_),
    .A2(_071_),
    .ZN(_072_));
 MUX2_X1 _436_ (.A(net1),
    .B(_260_),
    .S(_268_),
    .Z(_073_));
 NOR2_X1 _437_ (.A1(_010_),
    .A2(_073_),
    .ZN(_074_));
 NOR3_X1 _438_ (.A1(_070_),
    .A2(_072_),
    .A3(_074_),
    .ZN(_075_));
 MUX2_X1 _439_ (.A(_265_),
    .B(_266_),
    .S(_267_),
    .Z(_076_));
 MUX2_X1 _440_ (.A(_263_),
    .B(_264_),
    .S(_267_),
    .Z(_077_));
 MUX2_X1 _441_ (.A(_076_),
    .B(_077_),
    .S(_295_),
    .Z(_078_));
 AOI21_X1 _442_ (.A(_075_),
    .B1(_078_),
    .B2(_070_),
    .ZN(_079_));
 OR2_X1 _443_ (.A1(_010_),
    .A2(_070_),
    .ZN(_080_));
 NAND2_X2 _444_ (.A1(_014_),
    .A2(_018_),
    .ZN(_081_));
 NOR2_X1 _445_ (.A1(_080_),
    .A2(_081_),
    .ZN(_082_));
 AOI22_X1 _446_ (.A1(_068_),
    .A2(_058_),
    .B1(_292_),
    .B2(_082_),
    .ZN(_083_));
 OAI221_X1 _447_ (.A(_067_),
    .B1(_069_),
    .B2(_079_),
    .C1(_083_),
    .C2(_061_),
    .ZN(_084_));
 AND2_X1 _448_ (.A1(_013_),
    .A2(_084_),
    .ZN(_001_));
 INV_X2 _449_ (.A(_013_),
    .ZN(_085_));
 NOR2_X2 _450_ (.A1(_010_),
    .A2(_070_),
    .ZN(_086_));
 NOR2_X4 _451_ (.A1(_016_),
    .A2(_081_),
    .ZN(_087_));
 MUX2_X1 _452_ (.A(_260_),
    .B(net1),
    .S(_267_),
    .Z(_088_));
 NAND3_X1 _453_ (.A1(_086_),
    .A2(_087_),
    .A3(_088_),
    .ZN(_089_));
 AOI21_X1 _454_ (.A(_015_),
    .B1(_023_),
    .B2(_285_),
    .ZN(_090_));
 AOI21_X1 _455_ (.A(_090_),
    .B1(_286_),
    .B2(_068_),
    .ZN(_091_));
 INV_X1 _456_ (.A(_014_),
    .ZN(_092_));
 NAND2_X1 _457_ (.A1(_092_),
    .A2(_017_),
    .ZN(_093_));
 NAND2_X1 _458_ (.A1(_023_),
    .A2(_296_),
    .ZN(_094_));
 OAI21_X1 _459_ (.A(_094_),
    .B1(_299_),
    .B2(_023_),
    .ZN(_095_));
 OAI221_X1 _460_ (.A(_089_),
    .B1(_091_),
    .B2(_061_),
    .C1(_093_),
    .C2(_095_),
    .ZN(_096_));
 NOR2_X1 _461_ (.A1(_268_),
    .A2(_341_),
    .ZN(_097_));
 MUX2_X1 _462_ (.A(_264_),
    .B(_265_),
    .S(_268_),
    .Z(_098_));
 MUX2_X1 _463_ (.A(_097_),
    .B(_098_),
    .S(_295_),
    .Z(_099_));
 MUX2_X1 _464_ (.A(_262_),
    .B(_263_),
    .S(_268_),
    .Z(_100_));
 MUX2_X1 _465_ (.A(_260_),
    .B(_261_),
    .S(_268_),
    .Z(_101_));
 MUX2_X1 _466_ (.A(_100_),
    .B(_101_),
    .S(_295_),
    .Z(_102_));
 MUX2_X1 _467_ (.A(_099_),
    .B(_102_),
    .S(_302_),
    .Z(_103_));
 INV_X1 _468_ (.A(_069_),
    .ZN(_104_));
 AOI21_X1 _469_ (.A(_096_),
    .B1(_103_),
    .B2(_104_),
    .ZN(_105_));
 NAND2_X1 _470_ (.A1(_068_),
    .A2(_024_),
    .ZN(_106_));
 NOR2_X1 _471_ (.A1(_281_),
    .A2(_106_),
    .ZN(_107_));
 NOR3_X1 _472_ (.A1(_085_),
    .A2(_105_),
    .A3(_107_),
    .ZN(_002_));
 AND3_X1 _473_ (.A1(_295_),
    .A2(_070_),
    .A3(_076_),
    .ZN(_108_));
 NOR2_X1 _474_ (.A1(_295_),
    .A2(_070_),
    .ZN(_109_));
 AOI221_X2 _475_ (.A(_108_),
    .B1(_109_),
    .B2(_077_),
    .C1(_071_),
    .C2(_086_),
    .ZN(_110_));
 NOR2_X1 _476_ (.A1(_069_),
    .A2(_110_),
    .ZN(_111_));
 AOI21_X1 _477_ (.A(_023_),
    .B1(_034_),
    .B2(_015_),
    .ZN(_112_));
 NOR2_X1 _478_ (.A1(_070_),
    .A2(_081_),
    .ZN(_113_));
 MUX2_X1 _479_ (.A(_261_),
    .B(_260_),
    .S(_267_),
    .Z(_114_));
 MUX2_X1 _480_ (.A(_292_),
    .B(_114_),
    .S(_011_),
    .Z(_115_));
 AOI21_X1 _481_ (.A(_112_),
    .B1(_113_),
    .B2(_115_),
    .ZN(_116_));
 NOR2_X1 _482_ (.A1(_019_),
    .A2(_050_),
    .ZN(_117_));
 AOI21_X1 _483_ (.A(_117_),
    .B1(_303_),
    .B2(_023_),
    .ZN(_118_));
 XOR2_X2 _484_ (.A(_033_),
    .B(_284_),
    .Z(_119_));
 NOR2_X1 _485_ (.A1(_061_),
    .A2(_068_),
    .ZN(_120_));
 AOI22_X1 _486_ (.A1(_061_),
    .A2(_118_),
    .B1(_119_),
    .B2(_120_),
    .ZN(_121_));
 OAI22_X1 _487_ (.A1(_061_),
    .A2(_116_),
    .B1(_121_),
    .B2(_015_),
    .ZN(_122_));
 XOR2_X2 _488_ (.A(_280_),
    .B(_033_),
    .Z(_123_));
 OAI221_X1 _489_ (.A(_013_),
    .B1(_111_),
    .B2(_122_),
    .C1(_123_),
    .C2(_106_),
    .ZN(_124_));
 INV_X1 _490_ (.A(_124_),
    .ZN(_003_));
 NAND2_X1 _491_ (.A1(_019_),
    .A2(_024_),
    .ZN(_125_));
 XNOR2_X1 _492_ (.A(_028_),
    .B(_037_),
    .ZN(_126_));
 NOR2_X1 _493_ (.A1(_125_),
    .A2(_126_),
    .ZN(_127_));
 MUX2_X1 _494_ (.A(_262_),
    .B(_261_),
    .S(_267_),
    .Z(_128_));
 MUX2_X1 _495_ (.A(_088_),
    .B(_128_),
    .S(_011_),
    .Z(_129_));
 NAND3_X1 _496_ (.A1(_302_),
    .A2(_087_),
    .A3(_129_),
    .ZN(_130_));
 NAND3_X2 _497_ (.A1(_092_),
    .A2(_017_),
    .A3(_019_),
    .ZN(_131_));
 INV_X1 _498_ (.A(_315_),
    .ZN(_132_));
 AOI21_X1 _499_ (.A(_015_),
    .B1(_017_),
    .B2(_132_),
    .ZN(_133_));
 INV_X2 _500_ (.A(_016_),
    .ZN(_134_));
 AOI21_X1 _501_ (.A(_133_),
    .B1(_028_),
    .B2(_134_),
    .ZN(_135_));
 OAI221_X1 _502_ (.A(_130_),
    .B1(_131_),
    .B2(_311_),
    .C1(_023_),
    .C2(_135_),
    .ZN(_136_));
 NOR2_X1 _503_ (.A1(_127_),
    .A2(_136_),
    .ZN(_137_));
 NAND3_X1 _504_ (.A1(_070_),
    .A2(_288_),
    .A3(_266_),
    .ZN(_138_));
 NAND2_X1 _505_ (.A1(_302_),
    .A2(_100_),
    .ZN(_139_));
 AOI21_X1 _506_ (.A(_010_),
    .B1(_138_),
    .B2(_139_),
    .ZN(_140_));
 AOI21_X1 _507_ (.A(_140_),
    .B1(_109_),
    .B2(_098_),
    .ZN(_141_));
 OR2_X1 _508_ (.A1(_069_),
    .A2(_141_),
    .ZN(_142_));
 INV_X1 _509_ (.A(_050_),
    .ZN(_143_));
 AOI21_X2 _510_ (.A(_299_),
    .B1(_279_),
    .B2(_286_),
    .ZN(_144_));
 OAI21_X1 _511_ (.A(_143_),
    .B1(_144_),
    .B2(_034_),
    .ZN(_145_));
 XNOR2_X1 _512_ (.A(_028_),
    .B(_145_),
    .ZN(_146_));
 AOI221_X1 _513_ (.A(_085_),
    .B1(_137_),
    .B2(_142_),
    .C1(_146_),
    .C2(_020_),
    .ZN(_004_));
 INV_X1 _514_ (.A(_305_),
    .ZN(_147_));
 OR2_X1 _515_ (.A1(_033_),
    .A2(_284_),
    .ZN(_148_));
 AOI21_X1 _516_ (.A(_028_),
    .B1(_147_),
    .B2(_148_),
    .ZN(_149_));
 NOR2_X1 _517_ (.A1(_313_),
    .A2(_149_),
    .ZN(_150_));
 XNOR2_X1 _518_ (.A(_029_),
    .B(_150_),
    .ZN(_151_));
 OR2_X1 _519_ (.A1(_125_),
    .A2(_151_),
    .ZN(_152_));
 INV_X1 _520_ (.A(_323_),
    .ZN(_153_));
 AOI21_X1 _521_ (.A(_014_),
    .B1(_017_),
    .B2(_153_),
    .ZN(_154_));
 AOI21_X1 _522_ (.A(_154_),
    .B1(_029_),
    .B2(_134_),
    .ZN(_155_));
 OAI22_X2 _523_ (.A1(_319_),
    .A2(_131_),
    .B1(_155_),
    .B2(_019_),
    .ZN(_156_));
 NOR2_X1 _524_ (.A1(_070_),
    .A2(_069_),
    .ZN(_157_));
 AOI21_X1 _525_ (.A(_011_),
    .B1(_302_),
    .B2(_114_),
    .ZN(_158_));
 MUX2_X1 _526_ (.A(_263_),
    .B(_262_),
    .S(_267_),
    .Z(_159_));
 OAI22_X1 _527_ (.A1(_292_),
    .A2(_302_),
    .B1(_080_),
    .B2(_159_),
    .ZN(_160_));
 NOR2_X1 _528_ (.A1(_158_),
    .A2(_160_),
    .ZN(_161_));
 AOI221_X2 _529_ (.A(_156_),
    .B1(_157_),
    .B2(_078_),
    .C1(_087_),
    .C2(_161_),
    .ZN(_162_));
 AND3_X1 _530_ (.A1(_040_),
    .A2(_049_),
    .A3(_051_),
    .ZN(_163_));
 OR2_X1 _531_ (.A1(_052_),
    .A2(_163_),
    .ZN(_164_));
 AOI221_X1 _532_ (.A(_085_),
    .B1(_152_),
    .B2(_162_),
    .C1(_164_),
    .C2(_020_),
    .ZN(_005_));
 AOI21_X1 _533_ (.A(_323_),
    .B1(_029_),
    .B2(_315_),
    .ZN(_165_));
 NAND3_X1 _534_ (.A1(_033_),
    .A2(_028_),
    .A3(_029_),
    .ZN(_166_));
 NAND2_X1 _535_ (.A1(_050_),
    .A2(_028_),
    .ZN(_167_));
 OAI221_X2 _536_ (.A(_165_),
    .B1(_166_),
    .B2(_144_),
    .C1(_167_),
    .C2(_040_),
    .ZN(_168_));
 XOR2_X1 _537_ (.A(_042_),
    .B(_168_),
    .Z(_169_));
 OAI21_X1 _538_ (.A(_013_),
    .B1(_106_),
    .B2(_169_),
    .ZN(_170_));
 NAND2_X1 _539_ (.A1(_099_),
    .A2(_157_),
    .ZN(_171_));
 AOI21_X1 _540_ (.A(_014_),
    .B1(_017_),
    .B2(_048_),
    .ZN(_172_));
 AOI21_X1 _541_ (.A(_172_),
    .B1(_042_),
    .B2(_134_),
    .ZN(_173_));
 OAI221_X2 _542_ (.A(_171_),
    .B1(_131_),
    .B2(_327_),
    .C1(_023_),
    .C2(_173_),
    .ZN(_174_));
 INV_X1 _543_ (.A(_313_),
    .ZN(_175_));
 OAI21_X1 _544_ (.A(_175_),
    .B1(_037_),
    .B2(_028_),
    .ZN(_176_));
 AOI21_X2 _545_ (.A(_321_),
    .B1(_176_),
    .B2(_040_),
    .ZN(_177_));
 XOR2_X2 _546_ (.A(_042_),
    .B(_177_),
    .Z(_178_));
 AND2_X1 _547_ (.A1(_012_),
    .A2(_128_),
    .ZN(_179_));
 MUX2_X1 _548_ (.A(_264_),
    .B(_263_),
    .S(_267_),
    .Z(_180_));
 MUX2_X1 _549_ (.A(_088_),
    .B(_180_),
    .S(_012_),
    .Z(_181_));
 MUX2_X1 _550_ (.A(_179_),
    .B(_181_),
    .S(_011_),
    .Z(_182_));
 AOI221_X2 _551_ (.A(_174_),
    .B1(_178_),
    .B2(_025_),
    .C1(_087_),
    .C2(_182_),
    .ZN(_183_));
 NOR2_X1 _552_ (.A1(_170_),
    .A2(_183_),
    .ZN(_006_));
 NOR2_X1 _553_ (.A1(_019_),
    .A2(_080_),
    .ZN(_184_));
 NAND3_X1 _554_ (.A1(_015_),
    .A2(_076_),
    .A3(_184_),
    .ZN(_185_));
 NAND2_X1 _555_ (.A1(_092_),
    .A2(_019_),
    .ZN(_186_));
 OAI21_X1 _556_ (.A(_185_),
    .B1(_186_),
    .B2(_335_),
    .ZN(_187_));
 OAI21_X1 _557_ (.A(_092_),
    .B1(_134_),
    .B2(_047_),
    .ZN(_188_));
 OAI21_X1 _558_ (.A(_188_),
    .B1(_044_),
    .B2(_017_),
    .ZN(_189_));
 MUX2_X1 _559_ (.A(_265_),
    .B(_264_),
    .S(_267_),
    .Z(_190_));
 MUX2_X1 _560_ (.A(_159_),
    .B(_190_),
    .S(_011_),
    .Z(_191_));
 MUX2_X1 _561_ (.A(_115_),
    .B(_191_),
    .S(_302_),
    .Z(_192_));
 AOI222_X2 _562_ (.A1(_061_),
    .A2(_187_),
    .B1(_189_),
    .B2(_068_),
    .C1(_192_),
    .C2(_087_),
    .ZN(_193_));
 NOR2_X1 _563_ (.A1(_305_),
    .A2(_313_),
    .ZN(_194_));
 AOI221_X2 _564_ (.A(_029_),
    .B1(_148_),
    .B2(_194_),
    .C1(_175_),
    .C2(_312_),
    .ZN(_195_));
 NOR2_X1 _565_ (.A1(_321_),
    .A2(_195_),
    .ZN(_196_));
 OAI21_X1 _566_ (.A(_039_),
    .B1(_196_),
    .B2(_042_),
    .ZN(_197_));
 XNOR2_X1 _567_ (.A(_044_),
    .B(_197_),
    .ZN(_198_));
 OR2_X1 _568_ (.A1(_125_),
    .A2(_198_),
    .ZN(_199_));
 XNOR2_X1 _569_ (.A(_030_),
    .B(_054_),
    .ZN(_200_));
 AOI221_X1 _570_ (.A(_085_),
    .B1(_193_),
    .B2(_199_),
    .C1(_200_),
    .C2(_020_),
    .ZN(_007_));
 NAND3_X1 _571_ (.A1(_042_),
    .A2(_030_),
    .A3(_168_),
    .ZN(_201_));
 AOI21_X2 _572_ (.A(_047_),
    .B1(_030_),
    .B2(_331_),
    .ZN(_202_));
 NAND2_X1 _573_ (.A1(_201_),
    .A2(_202_),
    .ZN(_203_));
 XNOR2_X1 _574_ (.A(_022_),
    .B(_203_),
    .ZN(_204_));
 NAND3_X1 _575_ (.A1(_015_),
    .A2(_097_),
    .A3(_184_),
    .ZN(_205_));
 OAI21_X1 _576_ (.A(_205_),
    .B1(_186_),
    .B2(_343_),
    .ZN(_206_));
 OAI21_X1 _577_ (.A(_092_),
    .B1(_134_),
    .B2(_345_),
    .ZN(_207_));
 INV_X1 _578_ (.A(_022_),
    .ZN(_208_));
 OAI21_X1 _579_ (.A(_207_),
    .B1(_208_),
    .B2(_061_),
    .ZN(_209_));
 MUX2_X1 _580_ (.A(_266_),
    .B(_265_),
    .S(_267_),
    .Z(_210_));
 MUX2_X1 _581_ (.A(_180_),
    .B(_210_),
    .S(_011_),
    .Z(_211_));
 MUX2_X1 _582_ (.A(_129_),
    .B(_211_),
    .S(_302_),
    .Z(_212_));
 AOI222_X2 _583_ (.A1(_061_),
    .A2(_206_),
    .B1(_209_),
    .B2(_068_),
    .C1(_212_),
    .C2(_087_),
    .ZN(_213_));
 XNOR2_X1 _584_ (.A(_022_),
    .B(_045_),
    .ZN(_214_));
 OR2_X1 _585_ (.A1(_125_),
    .A2(_214_),
    .ZN(_215_));
 AOI221_X2 _586_ (.A(_085_),
    .B1(_020_),
    .B2(_204_),
    .C1(_213_),
    .C2(_215_),
    .ZN(_008_));
 NOR2_X1 _587_ (.A1(_030_),
    .A2(_047_),
    .ZN(_216_));
 XNOR2_X1 _588_ (.A(_208_),
    .B(_216_),
    .ZN(_217_));
 NAND3_X1 _589_ (.A1(_042_),
    .A2(_168_),
    .A3(_217_),
    .ZN(_218_));
 XNOR2_X1 _590_ (.A(_022_),
    .B(_202_),
    .ZN(_219_));
 OR2_X1 _591_ (.A1(_168_),
    .A2(_219_),
    .ZN(_220_));
 OAI21_X1 _592_ (.A(_218_),
    .B1(_220_),
    .B2(_042_),
    .ZN(_221_));
 NOR3_X1 _593_ (.A1(_058_),
    .A2(_085_),
    .A3(_123_),
    .ZN(_222_));
 AND3_X1 _594_ (.A1(_107_),
    .A2(_164_),
    .A3(_222_),
    .ZN(_223_));
 AND4_X1 _595_ (.A1(_146_),
    .A2(_200_),
    .A3(_221_),
    .A4(_223_),
    .ZN(_224_));
 MUX2_X1 _596_ (.A(_261_),
    .B(_263_),
    .S(_268_),
    .Z(_225_));
 NOR4_X1 _597_ (.A1(_295_),
    .A2(_070_),
    .A3(_262_),
    .A4(_225_),
    .ZN(_226_));
 AOI21_X1 _598_ (.A(_080_),
    .B1(_288_),
    .B2(net1),
    .ZN(_227_));
 AOI21_X1 _599_ (.A(_260_),
    .B1(_268_),
    .B2(_261_),
    .ZN(_228_));
 AOI21_X1 _600_ (.A(_226_),
    .B1(_227_),
    .B2(_228_),
    .ZN(_229_));
 NOR2_X1 _601_ (.A1(_295_),
    .A2(_098_),
    .ZN(_230_));
 AOI21_X1 _602_ (.A(_266_),
    .B1(_265_),
    .B2(_288_),
    .ZN(_231_));
 AOI21_X1 _603_ (.A(_230_),
    .B1(_231_),
    .B2(_295_),
    .ZN(_232_));
 OAI21_X1 _604_ (.A(_302_),
    .B1(_229_),
    .B2(_232_),
    .ZN(_233_));
 MUX2_X1 _605_ (.A(_263_),
    .B(_265_),
    .S(_268_),
    .Z(_234_));
 NOR3_X1 _606_ (.A1(_010_),
    .A2(_264_),
    .A3(_234_),
    .ZN(_235_));
 AOI21_X1 _607_ (.A(_235_),
    .B1(_231_),
    .B2(_010_),
    .ZN(_236_));
 NOR3_X1 _608_ (.A1(_069_),
    .A2(_140_),
    .A3(_236_),
    .ZN(_237_));
 NAND3_X1 _609_ (.A1(_110_),
    .A2(_233_),
    .A3(_237_),
    .ZN(_238_));
 NAND4_X1 _610_ (.A1(_319_),
    .A2(_327_),
    .A3(_335_),
    .A4(_343_),
    .ZN(_239_));
 NAND4_X1 _611_ (.A1(_289_),
    .A2(_296_),
    .A3(_303_),
    .A4(_311_),
    .ZN(_240_));
 OR3_X1 _612_ (.A1(_068_),
    .A2(_239_),
    .A3(_240_),
    .ZN(_241_));
 NOR4_X1 _613_ (.A1(_323_),
    .A2(_331_),
    .A3(_345_),
    .A4(_047_),
    .ZN(_242_));
 NOR4_X1 _614_ (.A1(_299_),
    .A2(_050_),
    .A3(_279_),
    .A4(_315_),
    .ZN(_243_));
 NAND3_X1 _615_ (.A1(_068_),
    .A2(_242_),
    .A3(_243_),
    .ZN(_244_));
 AOI21_X1 _616_ (.A(_093_),
    .B1(_241_),
    .B2(_244_),
    .ZN(_245_));
 NOR2_X1 _617_ (.A1(_161_),
    .A2(_182_),
    .ZN(_246_));
 NOR2_X1 _618_ (.A1(_115_),
    .A2(_129_),
    .ZN(_247_));
 OAI21_X1 _619_ (.A(_086_),
    .B1(_088_),
    .B2(_292_),
    .ZN(_248_));
 OAI21_X1 _620_ (.A(_302_),
    .B1(_191_),
    .B2(_211_),
    .ZN(_249_));
 AND4_X1 _621_ (.A1(_087_),
    .A2(_247_),
    .A3(_248_),
    .A4(_249_),
    .ZN(_250_));
 NAND3_X1 _622_ (.A1(_017_),
    .A2(_019_),
    .A3(_060_),
    .ZN(_251_));
 NAND2_X1 _623_ (.A1(_134_),
    .A2(_068_),
    .ZN(_252_));
 OAI21_X1 _624_ (.A(_251_),
    .B1(_252_),
    .B2(_060_),
    .ZN(_253_));
 AOI221_X2 _625_ (.A(_245_),
    .B1(_246_),
    .B2(_250_),
    .C1(_015_),
    .C2(_253_),
    .ZN(_254_));
 AOI21_X1 _626_ (.A(_085_),
    .B1(_238_),
    .B2(_254_),
    .ZN(_255_));
 XNOR2_X1 _627_ (.A(_042_),
    .B(_177_),
    .ZN(_256_));
 NOR4_X1 _628_ (.A1(_058_),
    .A2(_085_),
    .A3(_125_),
    .A4(_119_),
    .ZN(_257_));
 AND4_X1 _629_ (.A1(_285_),
    .A2(_126_),
    .A3(_151_),
    .A4(_257_),
    .ZN(_258_));
 AND4_X1 _630_ (.A1(_256_),
    .A2(_198_),
    .A3(_214_),
    .A4(_258_),
    .ZN(_259_));
 OR3_X1 _631_ (.A1(_224_),
    .A2(_255_),
    .A3(_259_),
    .ZN(_009_));
 FA_X1 _632_ (.A(net2),
    .B(net10),
    .CI(_279_),
    .CO(_280_),
    .S(_281_));
 FA_X1 _633_ (.A(_282_),
    .B(net10),
    .CI(_283_),
    .CO(_284_),
    .S(_285_));
 HA_X1 _634_ (.A(_287_),
    .B(_288_),
    .CO(_289_),
    .S(_290_));
 HA_X1 _635_ (.A(_287_),
    .B(net9),
    .CO(_283_),
    .S(_291_));
 HA_X1 _636_ (.A(net1),
    .B(_288_),
    .CO(_292_),
    .S(_293_));
 HA_X1 _637_ (.A(net1),
    .B(net9),
    .CO(_279_),
    .S(_294_));
 HA_X1 _638_ (.A(_282_),
    .B(_295_),
    .CO(_296_),
    .S(_286_));
 HA_X1 _639_ (.A(net2),
    .B(_295_),
    .CO(_297_),
    .S(_298_));
 HA_X1 _640_ (.A(net2),
    .B(net10),
    .CO(_299_),
    .S(_300_));
 HA_X1 _641_ (.A(_301_),
    .B(_302_),
    .CO(_303_),
    .S(_304_));
 HA_X1 _642_ (.A(net3),
    .B(_302_),
    .CO(_305_),
    .S(_306_));
 HA_X1 _643_ (.A(net3),
    .B(net11),
    .CO(_307_),
    .S(_308_));
 HA_X1 _644_ (.A(_309_),
    .B(_310_),
    .CO(_311_),
    .S(_312_));
 HA_X1 _645_ (.A(net4),
    .B(_310_),
    .CO(_313_),
    .S(_314_));
 HA_X1 _646_ (.A(net4),
    .B(net12),
    .CO(_315_),
    .S(_316_));
 HA_X1 _647_ (.A(_317_),
    .B(_318_),
    .CO(_319_),
    .S(_320_));
 HA_X1 _648_ (.A(net5),
    .B(_318_),
    .CO(_321_),
    .S(_322_));
 HA_X1 _649_ (.A(net5),
    .B(net13),
    .CO(_323_),
    .S(_324_));
 HA_X1 _650_ (.A(_325_),
    .B(_326_),
    .CO(_327_),
    .S(_328_));
 HA_X1 _651_ (.A(net6),
    .B(_326_),
    .CO(_329_),
    .S(_330_));
 HA_X1 _652_ (.A(net6),
    .B(net14),
    .CO(_331_),
    .S(_332_));
 HA_X1 _653_ (.A(_333_),
    .B(_334_),
    .CO(_335_),
    .S(_336_));
 HA_X1 _654_ (.A(net7),
    .B(_334_),
    .CO(_337_),
    .S(_338_));
 HA_X1 _655_ (.A(net7),
    .B(net15),
    .CO(_339_),
    .S(_340_));
 HA_X1 _656_ (.A(_341_),
    .B(_342_),
    .CO(_343_),
    .S(_344_));
 HA_X1 _657_ (.A(net8),
    .B(net16),
    .CO(_345_),
    .S(_346_));
 DFF_X1 \overflow_flag$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net17),
    .QN(_278_));
 DFF_X1 \result[0]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_277_));
 DFF_X1 \result[1]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_276_));
 DFF_X1 \result[2]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_275_));
 DFF_X1 \result[3]$_SDFF_PN0_  (.D(_004_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net21),
    .QN(_274_));
 DFF_X1 \result[4]$_SDFF_PN0_  (.D(_005_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net22),
    .QN(_273_));
 DFF_X1 \result[5]$_SDFF_PN0_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net23),
    .QN(_272_));
 DFF_X1 \result[6]$_SDFF_PN0_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net24),
    .QN(_271_));
 DFF_X1 \result[7]$_SDFF_PN0_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net25),
    .QN(_270_));
 DFF_X1 \zero_flag$_SDFF_PN0_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net26),
    .QN(_269_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_83 ();
 BUF_X2 input1 (.A(a[0]),
    .Z(net1));
 BUF_X2 input2 (.A(a[1]),
    .Z(net2));
 CLKBUF_X2 input3 (.A(a[2]),
    .Z(net3));
 BUF_X1 input4 (.A(a[3]),
    .Z(net4));
 BUF_X1 input5 (.A(a[4]),
    .Z(net5));
 BUF_X1 input6 (.A(a[5]),
    .Z(net6));
 BUF_X1 input7 (.A(a[6]),
    .Z(net7));
 BUF_X1 input8 (.A(a[7]),
    .Z(net8));
 BUF_X2 input9 (.A(b[0]),
    .Z(net9));
 BUF_X2 input10 (.A(b[1]),
    .Z(net10));
 BUF_X1 input11 (.A(b[2]),
    .Z(net11));
 BUF_X1 input12 (.A(b[3]),
    .Z(net12));
 BUF_X1 input13 (.A(b[4]),
    .Z(net13));
 BUF_X1 input14 (.A(b[5]),
    .Z(net14));
 BUF_X1 input15 (.A(b[6]),
    .Z(net15));
 BUF_X1 input16 (.A(b[7]),
    .Z(net16));
 BUF_X1 output17 (.A(net17),
    .Z(overflow_flag));
 BUF_X1 output18 (.A(net18),
    .Z(result[0]));
 BUF_X1 output19 (.A(net19),
    .Z(result[1]));
 BUF_X1 output20 (.A(net20),
    .Z(result[2]));
 BUF_X1 output21 (.A(net21),
    .Z(result[3]));
 BUF_X1 output22 (.A(net22),
    .Z(result[4]));
 BUF_X1 output23 (.A(net23),
    .Z(result[5]));
 BUF_X1 output24 (.A(net24),
    .Z(result[6]));
 BUF_X1 output25 (.A(net25),
    .Z(result[7]));
 BUF_X1 output26 (.A(net26),
    .Z(zero_flag));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_97 ();
 FILLCELL_X16 FILLER_0_104 ();
 FILLCELL_X8 FILLER_0_120 ();
 FILLCELL_X4 FILLER_0_128 ();
 FILLCELL_X2 FILLER_0_132 ();
 FILLCELL_X2 FILLER_0_137 ();
 FILLCELL_X1 FILLER_0_139 ();
 FILLCELL_X2 FILLER_0_143 ();
 FILLCELL_X1 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_149 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X32 FILLER_0_160 ();
 FILLCELL_X32 FILLER_0_192 ();
 FILLCELL_X32 FILLER_0_224 ();
 FILLCELL_X32 FILLER_0_256 ();
 FILLCELL_X16 FILLER_0_288 ();
 FILLCELL_X8 FILLER_0_304 ();
 FILLCELL_X2 FILLER_0_312 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X16 FILLER_1_289 ();
 FILLCELL_X8 FILLER_1_305 ();
 FILLCELL_X1 FILLER_1_313 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X16 FILLER_2_289 ();
 FILLCELL_X8 FILLER_2_305 ();
 FILLCELL_X1 FILLER_2_313 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X16 FILLER_3_289 ();
 FILLCELL_X8 FILLER_3_305 ();
 FILLCELL_X1 FILLER_3_313 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X16 FILLER_4_289 ();
 FILLCELL_X8 FILLER_4_305 ();
 FILLCELL_X1 FILLER_4_313 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X1 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_174 ();
 FILLCELL_X32 FILLER_5_206 ();
 FILLCELL_X32 FILLER_5_238 ();
 FILLCELL_X32 FILLER_5_270 ();
 FILLCELL_X8 FILLER_5_302 ();
 FILLCELL_X4 FILLER_5_310 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X1 FILLER_6_175 ();
 FILLCELL_X32 FILLER_6_180 ();
 FILLCELL_X32 FILLER_6_212 ();
 FILLCELL_X32 FILLER_6_244 ();
 FILLCELL_X32 FILLER_6_276 ();
 FILLCELL_X4 FILLER_6_308 ();
 FILLCELL_X2 FILLER_6_312 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X8 FILLER_7_161 ();
 FILLCELL_X1 FILLER_7_169 ();
 FILLCELL_X2 FILLER_7_182 ();
 FILLCELL_X32 FILLER_7_186 ();
 FILLCELL_X32 FILLER_7_218 ();
 FILLCELL_X32 FILLER_7_250 ();
 FILLCELL_X32 FILLER_7_282 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X16 FILLER_8_129 ();
 FILLCELL_X4 FILLER_8_145 ();
 FILLCELL_X2 FILLER_8_151 ();
 FILLCELL_X4 FILLER_8_163 ();
 FILLCELL_X2 FILLER_8_167 ();
 FILLCELL_X2 FILLER_8_171 ();
 FILLCELL_X32 FILLER_8_177 ();
 FILLCELL_X32 FILLER_8_209 ();
 FILLCELL_X32 FILLER_8_241 ();
 FILLCELL_X32 FILLER_8_273 ();
 FILLCELL_X8 FILLER_8_305 ();
 FILLCELL_X1 FILLER_8_313 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X16 FILLER_9_129 ();
 FILLCELL_X1 FILLER_9_145 ();
 FILLCELL_X8 FILLER_9_160 ();
 FILLCELL_X32 FILLER_9_182 ();
 FILLCELL_X32 FILLER_9_217 ();
 FILLCELL_X32 FILLER_9_249 ();
 FILLCELL_X32 FILLER_9_281 ();
 FILLCELL_X1 FILLER_9_313 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X8 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_163 ();
 FILLCELL_X2 FILLER_10_167 ();
 FILLCELL_X16 FILLER_10_183 ();
 FILLCELL_X8 FILLER_10_199 ();
 FILLCELL_X2 FILLER_10_214 ();
 FILLCELL_X2 FILLER_10_228 ();
 FILLCELL_X2 FILLER_10_239 ();
 FILLCELL_X32 FILLER_10_249 ();
 FILLCELL_X32 FILLER_10_281 ();
 FILLCELL_X1 FILLER_10_313 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_125 ();
 FILLCELL_X4 FILLER_11_157 ();
 FILLCELL_X2 FILLER_11_161 ();
 FILLCELL_X1 FILLER_11_163 ();
 FILLCELL_X8 FILLER_11_166 ();
 FILLCELL_X2 FILLER_11_174 ();
 FILLCELL_X2 FILLER_11_181 ();
 FILLCELL_X1 FILLER_11_183 ();
 FILLCELL_X16 FILLER_11_189 ();
 FILLCELL_X1 FILLER_11_205 ();
 FILLCELL_X4 FILLER_11_208 ();
 FILLCELL_X2 FILLER_11_212 ();
 FILLCELL_X1 FILLER_11_214 ();
 FILLCELL_X4 FILLER_11_218 ();
 FILLCELL_X2 FILLER_11_222 ();
 FILLCELL_X4 FILLER_11_227 ();
 FILLCELL_X4 FILLER_11_237 ();
 FILLCELL_X2 FILLER_11_241 ();
 FILLCELL_X32 FILLER_11_247 ();
 FILLCELL_X32 FILLER_11_279 ();
 FILLCELL_X2 FILLER_11_311 ();
 FILLCELL_X1 FILLER_11_313 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X8 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_105 ();
 FILLCELL_X1 FILLER_12_109 ();
 FILLCELL_X1 FILLER_12_114 ();
 FILLCELL_X32 FILLER_12_122 ();
 FILLCELL_X16 FILLER_12_154 ();
 FILLCELL_X4 FILLER_12_170 ();
 FILLCELL_X4 FILLER_12_183 ();
 FILLCELL_X2 FILLER_12_187 ();
 FILLCELL_X1 FILLER_12_189 ();
 FILLCELL_X4 FILLER_12_196 ();
 FILLCELL_X2 FILLER_12_200 ();
 FILLCELL_X1 FILLER_12_202 ();
 FILLCELL_X2 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_210 ();
 FILLCELL_X8 FILLER_12_227 ();
 FILLCELL_X4 FILLER_12_235 ();
 FILLCELL_X2 FILLER_12_239 ();
 FILLCELL_X16 FILLER_12_252 ();
 FILLCELL_X4 FILLER_12_268 ();
 FILLCELL_X2 FILLER_12_272 ();
 FILLCELL_X16 FILLER_12_294 ();
 FILLCELL_X1 FILLER_12_310 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_136 ();
 FILLCELL_X4 FILLER_13_168 ();
 FILLCELL_X1 FILLER_13_180 ();
 FILLCELL_X2 FILLER_13_187 ();
 FILLCELL_X4 FILLER_13_202 ();
 FILLCELL_X2 FILLER_13_210 ();
 FILLCELL_X1 FILLER_13_212 ();
 FILLCELL_X4 FILLER_13_220 ();
 FILLCELL_X1 FILLER_13_224 ();
 FILLCELL_X8 FILLER_13_231 ();
 FILLCELL_X2 FILLER_13_239 ();
 FILLCELL_X1 FILLER_13_241 ();
 FILLCELL_X16 FILLER_13_256 ();
 FILLCELL_X4 FILLER_13_272 ();
 FILLCELL_X16 FILLER_13_293 ();
 FILLCELL_X4 FILLER_13_309 ();
 FILLCELL_X1 FILLER_13_313 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X1 FILLER_14_113 ();
 FILLCELL_X4 FILLER_14_128 ();
 FILLCELL_X4 FILLER_14_134 ();
 FILLCELL_X1 FILLER_14_138 ();
 FILLCELL_X2 FILLER_14_145 ();
 FILLCELL_X16 FILLER_14_160 ();
 FILLCELL_X4 FILLER_14_176 ();
 FILLCELL_X16 FILLER_14_184 ();
 FILLCELL_X2 FILLER_14_200 ();
 FILLCELL_X1 FILLER_14_202 ();
 FILLCELL_X4 FILLER_14_211 ();
 FILLCELL_X2 FILLER_14_219 ();
 FILLCELL_X1 FILLER_14_221 ();
 FILLCELL_X4 FILLER_14_227 ();
 FILLCELL_X2 FILLER_14_231 ();
 FILLCELL_X4 FILLER_14_239 ();
 FILLCELL_X2 FILLER_14_249 ();
 FILLCELL_X16 FILLER_14_255 ();
 FILLCELL_X8 FILLER_14_271 ();
 FILLCELL_X4 FILLER_14_279 ();
 FILLCELL_X4 FILLER_14_308 ();
 FILLCELL_X2 FILLER_14_312 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X4 FILLER_15_25 ();
 FILLCELL_X2 FILLER_15_29 ();
 FILLCELL_X32 FILLER_15_37 ();
 FILLCELL_X16 FILLER_15_69 ();
 FILLCELL_X4 FILLER_15_85 ();
 FILLCELL_X2 FILLER_15_89 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X2 FILLER_15_117 ();
 FILLCELL_X4 FILLER_15_124 ();
 FILLCELL_X2 FILLER_15_128 ();
 FILLCELL_X2 FILLER_15_134 ();
 FILLCELL_X1 FILLER_15_136 ();
 FILLCELL_X4 FILLER_15_140 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X16 FILLER_15_169 ();
 FILLCELL_X4 FILLER_15_185 ();
 FILLCELL_X4 FILLER_15_200 ();
 FILLCELL_X8 FILLER_15_208 ();
 FILLCELL_X2 FILLER_15_216 ();
 FILLCELL_X1 FILLER_15_218 ();
 FILLCELL_X8 FILLER_15_228 ();
 FILLCELL_X4 FILLER_15_236 ();
 FILLCELL_X2 FILLER_15_240 ();
 FILLCELL_X1 FILLER_15_242 ();
 FILLCELL_X1 FILLER_15_249 ();
 FILLCELL_X16 FILLER_15_261 ();
 FILLCELL_X1 FILLER_15_277 ();
 FILLCELL_X2 FILLER_15_295 ();
 FILLCELL_X1 FILLER_15_297 ();
 FILLCELL_X8 FILLER_15_301 ();
 FILLCELL_X4 FILLER_15_309 ();
 FILLCELL_X1 FILLER_15_313 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_97 ();
 FILLCELL_X4 FILLER_16_105 ();
 FILLCELL_X1 FILLER_16_109 ();
 FILLCELL_X8 FILLER_16_126 ();
 FILLCELL_X4 FILLER_16_134 ();
 FILLCELL_X2 FILLER_16_138 ();
 FILLCELL_X2 FILLER_16_150 ();
 FILLCELL_X2 FILLER_16_159 ();
 FILLCELL_X8 FILLER_16_165 ();
 FILLCELL_X4 FILLER_16_173 ();
 FILLCELL_X1 FILLER_16_177 ();
 FILLCELL_X16 FILLER_16_227 ();
 FILLCELL_X2 FILLER_16_243 ();
 FILLCELL_X32 FILLER_16_249 ();
 FILLCELL_X32 FILLER_16_281 ();
 FILLCELL_X1 FILLER_16_313 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X16 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_113 ();
 FILLCELL_X4 FILLER_17_121 ();
 FILLCELL_X2 FILLER_17_125 ();
 FILLCELL_X32 FILLER_17_131 ();
 FILLCELL_X4 FILLER_17_165 ();
 FILLCELL_X1 FILLER_17_169 ();
 FILLCELL_X16 FILLER_17_175 ();
 FILLCELL_X4 FILLER_17_211 ();
 FILLCELL_X2 FILLER_17_215 ();
 FILLCELL_X4 FILLER_17_232 ();
 FILLCELL_X4 FILLER_17_239 ();
 FILLCELL_X32 FILLER_17_246 ();
 FILLCELL_X8 FILLER_17_278 ();
 FILLCELL_X4 FILLER_17_286 ();
 FILLCELL_X4 FILLER_17_310 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_165 ();
 FILLCELL_X2 FILLER_18_173 ();
 FILLCELL_X1 FILLER_18_175 ();
 FILLCELL_X4 FILLER_18_190 ();
 FILLCELL_X2 FILLER_18_194 ();
 FILLCELL_X1 FILLER_18_196 ();
 FILLCELL_X16 FILLER_18_204 ();
 FILLCELL_X2 FILLER_18_220 ();
 FILLCELL_X4 FILLER_18_225 ();
 FILLCELL_X1 FILLER_18_229 ();
 FILLCELL_X2 FILLER_18_233 ();
 FILLCELL_X1 FILLER_18_235 ();
 FILLCELL_X32 FILLER_18_242 ();
 FILLCELL_X32 FILLER_18_274 ();
 FILLCELL_X8 FILLER_18_306 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X8 FILLER_19_113 ();
 FILLCELL_X4 FILLER_19_121 ();
 FILLCELL_X16 FILLER_19_151 ();
 FILLCELL_X8 FILLER_19_167 ();
 FILLCELL_X4 FILLER_19_175 ();
 FILLCELL_X2 FILLER_19_179 ();
 FILLCELL_X4 FILLER_19_183 ();
 FILLCELL_X1 FILLER_19_195 ();
 FILLCELL_X8 FILLER_19_202 ();
 FILLCELL_X2 FILLER_19_210 ();
 FILLCELL_X8 FILLER_19_226 ();
 FILLCELL_X1 FILLER_19_234 ();
 FILLCELL_X16 FILLER_19_254 ();
 FILLCELL_X4 FILLER_19_270 ();
 FILLCELL_X1 FILLER_19_274 ();
 FILLCELL_X8 FILLER_19_300 ();
 FILLCELL_X4 FILLER_19_308 ();
 FILLCELL_X2 FILLER_19_312 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X2 FILLER_20_113 ();
 FILLCELL_X16 FILLER_20_142 ();
 FILLCELL_X2 FILLER_20_165 ();
 FILLCELL_X1 FILLER_20_167 ();
 FILLCELL_X2 FILLER_20_173 ();
 FILLCELL_X2 FILLER_20_187 ();
 FILLCELL_X1 FILLER_20_189 ();
 FILLCELL_X2 FILLER_20_194 ();
 FILLCELL_X16 FILLER_20_199 ();
 FILLCELL_X8 FILLER_20_215 ();
 FILLCELL_X2 FILLER_20_223 ();
 FILLCELL_X8 FILLER_20_228 ();
 FILLCELL_X4 FILLER_20_236 ();
 FILLCELL_X16 FILLER_20_256 ();
 FILLCELL_X8 FILLER_20_272 ();
 FILLCELL_X4 FILLER_20_280 ();
 FILLCELL_X1 FILLER_20_284 ();
 FILLCELL_X8 FILLER_20_302 ();
 FILLCELL_X1 FILLER_20_313 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_97 ();
 FILLCELL_X2 FILLER_21_105 ();
 FILLCELL_X1 FILLER_21_123 ();
 FILLCELL_X4 FILLER_21_142 ();
 FILLCELL_X4 FILLER_21_156 ();
 FILLCELL_X2 FILLER_21_160 ();
 FILLCELL_X1 FILLER_21_170 ();
 FILLCELL_X8 FILLER_21_175 ();
 FILLCELL_X1 FILLER_21_183 ();
 FILLCELL_X16 FILLER_21_197 ();
 FILLCELL_X8 FILLER_21_213 ();
 FILLCELL_X8 FILLER_21_229 ();
 FILLCELL_X4 FILLER_21_237 ();
 FILLCELL_X32 FILLER_21_247 ();
 FILLCELL_X32 FILLER_21_279 ();
 FILLCELL_X2 FILLER_21_311 ();
 FILLCELL_X1 FILLER_21_313 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_13 ();
 FILLCELL_X32 FILLER_22_45 ();
 FILLCELL_X32 FILLER_22_77 ();
 FILLCELL_X8 FILLER_22_109 ();
 FILLCELL_X2 FILLER_22_117 ();
 FILLCELL_X4 FILLER_22_126 ();
 FILLCELL_X16 FILLER_22_134 ();
 FILLCELL_X8 FILLER_22_150 ();
 FILLCELL_X16 FILLER_22_170 ();
 FILLCELL_X8 FILLER_22_186 ();
 FILLCELL_X4 FILLER_22_204 ();
 FILLCELL_X2 FILLER_22_208 ();
 FILLCELL_X1 FILLER_22_210 ();
 FILLCELL_X2 FILLER_22_237 ();
 FILLCELL_X32 FILLER_22_251 ();
 FILLCELL_X4 FILLER_22_283 ();
 FILLCELL_X1 FILLER_22_287 ();
 FILLCELL_X8 FILLER_22_305 ();
 FILLCELL_X1 FILLER_22_313 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_117 ();
 FILLCELL_X32 FILLER_23_128 ();
 FILLCELL_X4 FILLER_23_160 ();
 FILLCELL_X2 FILLER_23_164 ();
 FILLCELL_X16 FILLER_23_177 ();
 FILLCELL_X1 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_211 ();
 FILLCELL_X4 FILLER_23_215 ();
 FILLCELL_X1 FILLER_23_219 ();
 FILLCELL_X8 FILLER_23_232 ();
 FILLCELL_X16 FILLER_23_246 ();
 FILLCELL_X8 FILLER_23_262 ();
 FILLCELL_X4 FILLER_23_270 ();
 FILLCELL_X8 FILLER_23_276 ();
 FILLCELL_X1 FILLER_23_284 ();
 FILLCELL_X4 FILLER_23_308 ();
 FILLCELL_X2 FILLER_23_312 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X16 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_113 ();
 FILLCELL_X32 FILLER_24_124 ();
 FILLCELL_X16 FILLER_24_156 ();
 FILLCELL_X2 FILLER_24_175 ();
 FILLCELL_X2 FILLER_24_184 ();
 FILLCELL_X1 FILLER_24_204 ();
 FILLCELL_X4 FILLER_24_230 ();
 FILLCELL_X2 FILLER_24_234 ();
 FILLCELL_X1 FILLER_24_236 ();
 FILLCELL_X32 FILLER_24_241 ();
 FILLCELL_X16 FILLER_24_273 ();
 FILLCELL_X4 FILLER_24_289 ();
 FILLCELL_X1 FILLER_24_293 ();
 FILLCELL_X8 FILLER_24_299 ();
 FILLCELL_X4 FILLER_24_307 ();
 FILLCELL_X2 FILLER_24_311 ();
 FILLCELL_X1 FILLER_24_313 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_17 ();
 FILLCELL_X1 FILLER_25_19 ();
 FILLCELL_X32 FILLER_25_24 ();
 FILLCELL_X32 FILLER_25_56 ();
 FILLCELL_X16 FILLER_25_88 ();
 FILLCELL_X4 FILLER_25_104 ();
 FILLCELL_X2 FILLER_25_108 ();
 FILLCELL_X4 FILLER_25_122 ();
 FILLCELL_X2 FILLER_25_126 ();
 FILLCELL_X2 FILLER_25_140 ();
 FILLCELL_X4 FILLER_25_149 ();
 FILLCELL_X2 FILLER_25_153 ();
 FILLCELL_X1 FILLER_25_155 ();
 FILLCELL_X2 FILLER_25_166 ();
 FILLCELL_X1 FILLER_25_168 ();
 FILLCELL_X16 FILLER_25_173 ();
 FILLCELL_X2 FILLER_25_189 ();
 FILLCELL_X1 FILLER_25_191 ();
 FILLCELL_X4 FILLER_25_195 ();
 FILLCELL_X1 FILLER_25_199 ();
 FILLCELL_X2 FILLER_25_207 ();
 FILLCELL_X2 FILLER_25_223 ();
 FILLCELL_X1 FILLER_25_225 ();
 FILLCELL_X4 FILLER_25_240 ();
 FILLCELL_X2 FILLER_25_251 ();
 FILLCELL_X1 FILLER_25_253 ();
 FILLCELL_X16 FILLER_25_258 ();
 FILLCELL_X8 FILLER_25_274 ();
 FILLCELL_X4 FILLER_25_286 ();
 FILLCELL_X2 FILLER_25_307 ();
 FILLCELL_X1 FILLER_25_309 ();
 FILLCELL_X1 FILLER_25_313 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_17 ();
 FILLCELL_X1 FILLER_26_19 ();
 FILLCELL_X32 FILLER_26_24 ();
 FILLCELL_X32 FILLER_26_56 ();
 FILLCELL_X16 FILLER_26_88 ();
 FILLCELL_X4 FILLER_26_104 ();
 FILLCELL_X1 FILLER_26_108 ();
 FILLCELL_X4 FILLER_26_119 ();
 FILLCELL_X1 FILLER_26_123 ();
 FILLCELL_X4 FILLER_26_128 ();
 FILLCELL_X1 FILLER_26_132 ();
 FILLCELL_X1 FILLER_26_144 ();
 FILLCELL_X4 FILLER_26_152 ();
 FILLCELL_X1 FILLER_26_163 ();
 FILLCELL_X16 FILLER_26_171 ();
 FILLCELL_X8 FILLER_26_187 ();
 FILLCELL_X2 FILLER_26_195 ();
 FILLCELL_X1 FILLER_26_197 ();
 FILLCELL_X4 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_206 ();
 FILLCELL_X1 FILLER_26_208 ();
 FILLCELL_X4 FILLER_26_212 ();
 FILLCELL_X8 FILLER_26_219 ();
 FILLCELL_X2 FILLER_26_227 ();
 FILLCELL_X1 FILLER_26_229 ();
 FILLCELL_X4 FILLER_26_235 ();
 FILLCELL_X2 FILLER_26_239 ();
 FILLCELL_X1 FILLER_26_241 ();
 FILLCELL_X32 FILLER_26_246 ();
 FILLCELL_X32 FILLER_26_278 ();
 FILLCELL_X4 FILLER_26_310 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X16 FILLER_27_97 ();
 FILLCELL_X2 FILLER_27_113 ();
 FILLCELL_X4 FILLER_27_122 ();
 FILLCELL_X2 FILLER_27_126 ();
 FILLCELL_X1 FILLER_27_128 ();
 FILLCELL_X2 FILLER_27_136 ();
 FILLCELL_X1 FILLER_27_138 ();
 FILLCELL_X1 FILLER_27_142 ();
 FILLCELL_X8 FILLER_27_147 ();
 FILLCELL_X2 FILLER_27_155 ();
 FILLCELL_X1 FILLER_27_157 ();
 FILLCELL_X2 FILLER_27_162 ();
 FILLCELL_X1 FILLER_27_164 ();
 FILLCELL_X2 FILLER_27_180 ();
 FILLCELL_X8 FILLER_27_189 ();
 FILLCELL_X8 FILLER_27_201 ();
 FILLCELL_X2 FILLER_27_209 ();
 FILLCELL_X32 FILLER_27_215 ();
 FILLCELL_X32 FILLER_27_247 ();
 FILLCELL_X32 FILLER_27_279 ();
 FILLCELL_X2 FILLER_27_311 ();
 FILLCELL_X1 FILLER_27_313 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X16 FILLER_28_97 ();
 FILLCELL_X8 FILLER_28_113 ();
 FILLCELL_X4 FILLER_28_121 ();
 FILLCELL_X2 FILLER_28_125 ();
 FILLCELL_X1 FILLER_28_127 ();
 FILLCELL_X4 FILLER_28_140 ();
 FILLCELL_X1 FILLER_28_144 ();
 FILLCELL_X1 FILLER_28_148 ();
 FILLCELL_X4 FILLER_28_153 ();
 FILLCELL_X2 FILLER_28_190 ();
 FILLCELL_X32 FILLER_28_209 ();
 FILLCELL_X32 FILLER_28_241 ();
 FILLCELL_X32 FILLER_28_273 ();
 FILLCELL_X8 FILLER_28_305 ();
 FILLCELL_X1 FILLER_28_313 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X4 FILLER_29_129 ();
 FILLCELL_X1 FILLER_29_133 ();
 FILLCELL_X8 FILLER_29_146 ();
 FILLCELL_X2 FILLER_29_154 ();
 FILLCELL_X8 FILLER_29_164 ();
 FILLCELL_X2 FILLER_29_172 ();
 FILLCELL_X1 FILLER_29_174 ();
 FILLCELL_X2 FILLER_29_178 ();
 FILLCELL_X1 FILLER_29_180 ();
 FILLCELL_X16 FILLER_29_184 ();
 FILLCELL_X1 FILLER_29_200 ();
 FILLCELL_X32 FILLER_29_208 ();
 FILLCELL_X32 FILLER_29_240 ();
 FILLCELL_X32 FILLER_29_272 ();
 FILLCELL_X8 FILLER_29_304 ();
 FILLCELL_X2 FILLER_29_312 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X8 FILLER_30_97 ();
 FILLCELL_X2 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_107 ();
 FILLCELL_X4 FILLER_30_121 ();
 FILLCELL_X2 FILLER_30_125 ();
 FILLCELL_X1 FILLER_30_134 ();
 FILLCELL_X2 FILLER_30_143 ();
 FILLCELL_X2 FILLER_30_152 ();
 FILLCELL_X4 FILLER_30_161 ();
 FILLCELL_X1 FILLER_30_165 ();
 FILLCELL_X4 FILLER_30_173 ();
 FILLCELL_X2 FILLER_30_177 ();
 FILLCELL_X1 FILLER_30_179 ();
 FILLCELL_X4 FILLER_30_187 ();
 FILLCELL_X1 FILLER_30_203 ();
 FILLCELL_X1 FILLER_30_208 ();
 FILLCELL_X32 FILLER_30_212 ();
 FILLCELL_X32 FILLER_30_244 ();
 FILLCELL_X32 FILLER_30_276 ();
 FILLCELL_X4 FILLER_30_308 ();
 FILLCELL_X2 FILLER_30_312 ();
 FILLCELL_X16 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_17 ();
 FILLCELL_X4 FILLER_31_21 ();
 FILLCELL_X2 FILLER_31_25 ();
 FILLCELL_X1 FILLER_31_27 ();
 FILLCELL_X32 FILLER_31_32 ();
 FILLCELL_X32 FILLER_31_64 ();
 FILLCELL_X16 FILLER_31_96 ();
 FILLCELL_X4 FILLER_31_142 ();
 FILLCELL_X4 FILLER_31_156 ();
 FILLCELL_X1 FILLER_31_160 ();
 FILLCELL_X1 FILLER_31_168 ();
 FILLCELL_X2 FILLER_31_176 ();
 FILLCELL_X4 FILLER_31_199 ();
 FILLCELL_X32 FILLER_31_214 ();
 FILLCELL_X32 FILLER_31_246 ();
 FILLCELL_X32 FILLER_31_278 ();
 FILLCELL_X4 FILLER_31_310 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X8 FILLER_32_129 ();
 FILLCELL_X4 FILLER_32_137 ();
 FILLCELL_X1 FILLER_32_141 ();
 FILLCELL_X8 FILLER_32_149 ();
 FILLCELL_X2 FILLER_32_157 ();
 FILLCELL_X4 FILLER_32_173 ();
 FILLCELL_X4 FILLER_32_184 ();
 FILLCELL_X32 FILLER_32_199 ();
 FILLCELL_X32 FILLER_32_231 ();
 FILLCELL_X32 FILLER_32_263 ();
 FILLCELL_X16 FILLER_32_295 ();
 FILLCELL_X2 FILLER_32_311 ();
 FILLCELL_X1 FILLER_32_313 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X16 FILLER_33_289 ();
 FILLCELL_X8 FILLER_33_305 ();
 FILLCELL_X1 FILLER_33_313 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X16 FILLER_34_289 ();
 FILLCELL_X8 FILLER_34_305 ();
 FILLCELL_X1 FILLER_34_313 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X16 FILLER_35_289 ();
 FILLCELL_X8 FILLER_35_305 ();
 FILLCELL_X1 FILLER_35_313 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X16 FILLER_36_289 ();
 FILLCELL_X8 FILLER_36_305 ();
 FILLCELL_X1 FILLER_36_313 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X16 FILLER_37_289 ();
 FILLCELL_X8 FILLER_37_305 ();
 FILLCELL_X1 FILLER_37_313 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X16 FILLER_38_289 ();
 FILLCELL_X8 FILLER_38_305 ();
 FILLCELL_X1 FILLER_38_313 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X16 FILLER_39_289 ();
 FILLCELL_X8 FILLER_39_305 ();
 FILLCELL_X1 FILLER_39_313 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X16 FILLER_40_289 ();
 FILLCELL_X8 FILLER_40_305 ();
 FILLCELL_X1 FILLER_40_313 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X8 FILLER_41_97 ();
 FILLCELL_X4 FILLER_41_105 ();
 FILLCELL_X32 FILLER_41_113 ();
 FILLCELL_X32 FILLER_41_145 ();
 FILLCELL_X32 FILLER_41_177 ();
 FILLCELL_X4 FILLER_41_209 ();
 FILLCELL_X2 FILLER_41_213 ();
 FILLCELL_X32 FILLER_41_222 ();
 FILLCELL_X32 FILLER_41_254 ();
 FILLCELL_X16 FILLER_41_286 ();
 FILLCELL_X8 FILLER_41_302 ();
 FILLCELL_X4 FILLER_41_310 ();
endmodule
