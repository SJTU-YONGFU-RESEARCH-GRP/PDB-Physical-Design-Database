module wishbone_master (clk,
    read_done,
    read_err,
    read_req,
    rst_n,
    wb_ack_i,
    wb_cyc_o,
    wb_err_i,
    wb_rty_i,
    wb_stb_o,
    wb_tgd_i,
    wb_tgd_o,
    wb_we_o,
    write_done,
    write_err,
    write_req,
    read_addr,
    read_data,
    read_sel,
    wb_adr_o,
    wb_dat_i,
    wb_dat_o,
    wb_sel_o,
    write_addr,
    write_data,
    write_sel);
 input clk;
 output read_done;
 output read_err;
 input read_req;
 input rst_n;
 input wb_ack_i;
 output wb_cyc_o;
 input wb_err_i;
 input wb_rty_i;
 output wb_stb_o;
 input wb_tgd_i;
 output wb_tgd_o;
 output wb_we_o;
 output write_done;
 output write_err;
 input write_req;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [3:0] read_sel;
 output [31:0] wb_adr_o;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 output [3:0] wb_sel_o;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_sel;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire clknet_0_clk;
 wire \retry_count[0] ;
 wire \retry_count[1] ;
 wire \retry_count[2] ;
 wire \retry_count[3] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X4 _464_ (.A(\state[1] ),
    .Z(_116_));
 BUF_X4 _465_ (.A(\state[2] ),
    .Z(_117_));
 OR2_X1 _466_ (.A1(_116_),
    .A2(_117_),
    .ZN(_118_));
 BUF_X4 _467_ (.A(_118_),
    .Z(_119_));
 BUF_X2 _468_ (.A(wb_ack_i),
    .Z(_120_));
 OAI21_X1 _469_ (.A(_119_),
    .B1(net69),
    .B2(_120_),
    .ZN(_121_));
 BUF_X2 _470_ (.A(rst_n),
    .Z(_122_));
 INV_X4 _471_ (.A(_122_),
    .ZN(_123_));
 BUF_X2 _472_ (.A(\state[3] ),
    .Z(_124_));
 AOI21_X1 _473_ (.A(_123_),
    .B1(_124_),
    .B2(\retry_count[3] ),
    .ZN(_125_));
 CLKBUF_X3 _474_ (.A(\state[0] ),
    .Z(_126_));
 BUF_X2 _475_ (.A(read_req),
    .Z(_127_));
 BUF_X4 _476_ (.A(write_req),
    .Z(_128_));
 NOR2_X2 _477_ (.A1(_127_),
    .A2(_128_),
    .ZN(_129_));
 NAND2_X1 _478_ (.A1(_126_),
    .A2(_129_),
    .ZN(_130_));
 NAND3_X1 _479_ (.A1(_121_),
    .A2(_125_),
    .A3(_130_),
    .ZN(_001_));
 CLKBUF_X3 _480_ (.A(_122_),
    .Z(_131_));
 CLKBUF_X2 _481_ (.A(_131_),
    .Z(_132_));
 INV_X1 _482_ (.A(_128_),
    .ZN(_133_));
 NAND3_X1 _483_ (.A1(_127_),
    .A2(_133_),
    .A3(_126_),
    .ZN(_134_));
 INV_X1 _484_ (.A(\retry_count[3] ),
    .ZN(_135_));
 NAND2_X1 _485_ (.A1(_135_),
    .A2(_124_),
    .ZN(_136_));
 OR3_X1 _486_ (.A1(_120_),
    .A2(net69),
    .A3(net70),
    .ZN(_137_));
 INV_X1 _487_ (.A(_116_),
    .ZN(_138_));
 OAI221_X1 _488_ (.A(_134_),
    .B1(_136_),
    .B2(net243),
    .C1(_137_),
    .C2(_138_),
    .ZN(_139_));
 AND2_X1 _489_ (.A1(_132_),
    .A2(_139_),
    .ZN(_002_));
 NAND2_X2 _490_ (.A1(_128_),
    .A2(_126_),
    .ZN(_140_));
 CLKBUF_X3 _491_ (.A(_140_),
    .Z(_141_));
 INV_X1 _492_ (.A(net243),
    .ZN(_142_));
 INV_X1 _493_ (.A(_117_),
    .ZN(_143_));
 OAI221_X1 _494_ (.A(_141_),
    .B1(_136_),
    .B2(_142_),
    .C1(_143_),
    .C2(_137_),
    .ZN(_144_));
 AND2_X1 _495_ (.A1(_132_),
    .A2(_144_),
    .ZN(_003_));
 NOR2_X2 _496_ (.A1(_120_),
    .A2(net69),
    .ZN(_145_));
 NAND3_X2 _497_ (.A1(net70),
    .A2(_119_),
    .A3(_145_),
    .ZN(_146_));
 NOR2_X1 _498_ (.A1(_123_),
    .A2(_146_),
    .ZN(_000_));
 NAND2_X2 _499_ (.A1(_120_),
    .A2(_116_),
    .ZN(_147_));
 CLKBUF_X3 _500_ (.A(_147_),
    .Z(_148_));
 MUX2_X1 _501_ (.A(net37),
    .B(net139),
    .S(_148_),
    .Z(_149_));
 AND2_X1 _502_ (.A1(_132_),
    .A2(_149_),
    .ZN(_006_));
 MUX2_X1 _503_ (.A(net38),
    .B(net140),
    .S(_148_),
    .Z(_150_));
 AND2_X1 _504_ (.A1(_132_),
    .A2(_150_),
    .ZN(_007_));
 MUX2_X1 _505_ (.A(net39),
    .B(net141),
    .S(_148_),
    .Z(_151_));
 AND2_X1 _506_ (.A1(_132_),
    .A2(_151_),
    .ZN(_008_));
 MUX2_X1 _507_ (.A(net40),
    .B(net142),
    .S(_148_),
    .Z(_152_));
 AND2_X1 _508_ (.A1(_132_),
    .A2(_152_),
    .ZN(_009_));
 MUX2_X1 _509_ (.A(net41),
    .B(net143),
    .S(_148_),
    .Z(_153_));
 AND2_X1 _510_ (.A1(_132_),
    .A2(_153_),
    .ZN(_010_));
 MUX2_X1 _511_ (.A(net42),
    .B(net144),
    .S(_148_),
    .Z(_154_));
 AND2_X1 _512_ (.A1(_132_),
    .A2(_154_),
    .ZN(_011_));
 MUX2_X1 _513_ (.A(net43),
    .B(net145),
    .S(_148_),
    .Z(_155_));
 AND2_X1 _514_ (.A1(_132_),
    .A2(_155_),
    .ZN(_012_));
 MUX2_X1 _515_ (.A(net44),
    .B(net146),
    .S(_148_),
    .Z(_156_));
 AND2_X1 _516_ (.A1(_132_),
    .A2(_156_),
    .ZN(_013_));
 CLKBUF_X2 _517_ (.A(_131_),
    .Z(_157_));
 MUX2_X1 _518_ (.A(net45),
    .B(net147),
    .S(_148_),
    .Z(_158_));
 AND2_X1 _519_ (.A1(_157_),
    .A2(_158_),
    .ZN(_014_));
 CLKBUF_X3 _520_ (.A(_147_),
    .Z(_159_));
 MUX2_X1 _521_ (.A(net46),
    .B(net148),
    .S(_159_),
    .Z(_160_));
 AND2_X1 _522_ (.A1(_157_),
    .A2(_160_),
    .ZN(_015_));
 MUX2_X1 _523_ (.A(net47),
    .B(net149),
    .S(_159_),
    .Z(_161_));
 AND2_X1 _524_ (.A1(_157_),
    .A2(_161_),
    .ZN(_016_));
 MUX2_X1 _525_ (.A(net48),
    .B(net150),
    .S(_159_),
    .Z(_162_));
 AND2_X1 _526_ (.A1(_157_),
    .A2(_162_),
    .ZN(_017_));
 MUX2_X1 _527_ (.A(net49),
    .B(net151),
    .S(_159_),
    .Z(_163_));
 AND2_X1 _528_ (.A1(_157_),
    .A2(_163_),
    .ZN(_018_));
 MUX2_X1 _529_ (.A(net50),
    .B(net152),
    .S(_159_),
    .Z(_164_));
 AND2_X1 _530_ (.A1(_157_),
    .A2(_164_),
    .ZN(_019_));
 MUX2_X1 _531_ (.A(net51),
    .B(net153),
    .S(_159_),
    .Z(_165_));
 AND2_X1 _532_ (.A1(_157_),
    .A2(_165_),
    .ZN(_020_));
 MUX2_X1 _533_ (.A(net52),
    .B(net154),
    .S(_159_),
    .Z(_166_));
 AND2_X1 _534_ (.A1(_157_),
    .A2(_166_),
    .ZN(_021_));
 MUX2_X1 _535_ (.A(net53),
    .B(net155),
    .S(_159_),
    .Z(_167_));
 AND2_X1 _536_ (.A1(_157_),
    .A2(_167_),
    .ZN(_022_));
 MUX2_X1 _537_ (.A(net54),
    .B(net156),
    .S(_159_),
    .Z(_168_));
 AND2_X1 _538_ (.A1(_157_),
    .A2(_168_),
    .ZN(_023_));
 BUF_X2 _539_ (.A(_131_),
    .Z(_169_));
 MUX2_X1 _540_ (.A(net55),
    .B(net157),
    .S(_159_),
    .Z(_170_));
 AND2_X1 _541_ (.A1(_169_),
    .A2(_170_),
    .ZN(_024_));
 CLKBUF_X3 _542_ (.A(_147_),
    .Z(_171_));
 MUX2_X1 _543_ (.A(net56),
    .B(net158),
    .S(_171_),
    .Z(_172_));
 AND2_X1 _544_ (.A1(_169_),
    .A2(_172_),
    .ZN(_025_));
 MUX2_X1 _545_ (.A(net57),
    .B(net159),
    .S(_171_),
    .Z(_173_));
 AND2_X1 _546_ (.A1(_169_),
    .A2(_173_),
    .ZN(_026_));
 MUX2_X1 _547_ (.A(net58),
    .B(net160),
    .S(_171_),
    .Z(_174_));
 AND2_X1 _548_ (.A1(_169_),
    .A2(_174_),
    .ZN(_027_));
 MUX2_X1 _549_ (.A(net59),
    .B(net161),
    .S(_171_),
    .Z(_175_));
 AND2_X1 _550_ (.A1(_169_),
    .A2(_175_),
    .ZN(_028_));
 MUX2_X1 _551_ (.A(net60),
    .B(net162),
    .S(_171_),
    .Z(_176_));
 AND2_X1 _552_ (.A1(_169_),
    .A2(_176_),
    .ZN(_029_));
 MUX2_X1 _553_ (.A(net61),
    .B(net163),
    .S(_171_),
    .Z(_177_));
 AND2_X1 _554_ (.A1(_169_),
    .A2(_177_),
    .ZN(_030_));
 MUX2_X1 _555_ (.A(net62),
    .B(net164),
    .S(_171_),
    .Z(_178_));
 AND2_X1 _556_ (.A1(_169_),
    .A2(_178_),
    .ZN(_031_));
 MUX2_X1 _557_ (.A(net63),
    .B(net165),
    .S(_171_),
    .Z(_179_));
 AND2_X1 _558_ (.A1(_169_),
    .A2(_179_),
    .ZN(_032_));
 MUX2_X1 _559_ (.A(net64),
    .B(net166),
    .S(_171_),
    .Z(_180_));
 AND2_X1 _560_ (.A1(_169_),
    .A2(_180_),
    .ZN(_033_));
 BUF_X2 _561_ (.A(_131_),
    .Z(_181_));
 MUX2_X1 _562_ (.A(net65),
    .B(net167),
    .S(_171_),
    .Z(_182_));
 AND2_X1 _563_ (.A1(_181_),
    .A2(_182_),
    .ZN(_034_));
 MUX2_X1 _564_ (.A(net66),
    .B(net168),
    .S(_147_),
    .Z(_183_));
 AND2_X1 _565_ (.A1(_181_),
    .A2(_183_),
    .ZN(_035_));
 MUX2_X1 _566_ (.A(net67),
    .B(net169),
    .S(_147_),
    .Z(_184_));
 AND2_X1 _567_ (.A1(_181_),
    .A2(_184_),
    .ZN(_036_));
 MUX2_X1 _568_ (.A(net68),
    .B(net170),
    .S(_147_),
    .Z(_185_));
 AND2_X1 _569_ (.A1(_181_),
    .A2(_185_),
    .ZN(_037_));
 INV_X1 _570_ (.A(net171),
    .ZN(_186_));
 INV_X1 _571_ (.A(_127_),
    .ZN(_187_));
 BUF_X4 _572_ (.A(_128_),
    .Z(_188_));
 NOR2_X1 _573_ (.A1(_187_),
    .A2(_188_),
    .ZN(_189_));
 MUX2_X1 _574_ (.A(_186_),
    .B(_138_),
    .S(_189_),
    .Z(_190_));
 AOI221_X1 _575_ (.A(_123_),
    .B1(_186_),
    .B2(_148_),
    .C1(_190_),
    .C2(_126_),
    .ZN(_038_));
 INV_X1 _576_ (.A(_126_),
    .ZN(_191_));
 AOI21_X1 _577_ (.A(_191_),
    .B1(_133_),
    .B2(_127_),
    .ZN(_192_));
 INV_X1 _578_ (.A(_004_),
    .ZN(_193_));
 NOR2_X1 _579_ (.A1(_126_),
    .A2(_193_),
    .ZN(_194_));
 NOR4_X2 _580_ (.A1(_124_),
    .A2(_116_),
    .A3(_192_),
    .A4(_194_),
    .ZN(_195_));
 OAI21_X1 _581_ (.A(_124_),
    .B1(net243),
    .B2(_135_),
    .ZN(_196_));
 AOI21_X1 _582_ (.A(_116_),
    .B1(_004_),
    .B2(_191_),
    .ZN(_197_));
 INV_X1 _583_ (.A(net69),
    .ZN(_198_));
 NOR3_X1 _584_ (.A1(_120_),
    .A2(_138_),
    .A3(_198_),
    .ZN(_199_));
 OAI221_X2 _585_ (.A(_196_),
    .B1(_197_),
    .B2(_199_),
    .C1(_189_),
    .C2(_191_),
    .ZN(_200_));
 INV_X1 _586_ (.A(net172),
    .ZN(_201_));
 AOI211_X2 _587_ (.A(_123_),
    .B(_195_),
    .C1(_200_),
    .C2(_201_),
    .ZN(_039_));
 BUF_X2 _588_ (.A(_005_),
    .Z(_202_));
 OR3_X1 _589_ (.A1(_116_),
    .A2(_117_),
    .A3(_202_),
    .ZN(_203_));
 NAND2_X1 _590_ (.A1(\retry_count[0] ),
    .A2(_203_),
    .ZN(_204_));
 MUX2_X1 _591_ (.A(\retry_count[0] ),
    .B(_204_),
    .S(_146_),
    .Z(_205_));
 NOR2_X1 _592_ (.A1(_123_),
    .A2(_205_),
    .ZN(_040_));
 NAND4_X1 _593_ (.A1(net70),
    .A2(_462_),
    .A3(_119_),
    .A4(_145_),
    .ZN(_206_));
 NAND3_X1 _594_ (.A1(\retry_count[1] ),
    .A2(_146_),
    .A3(_203_),
    .ZN(_207_));
 AOI21_X1 _595_ (.A(_123_),
    .B1(_206_),
    .B2(_207_),
    .ZN(_041_));
 INV_X1 _596_ (.A(_461_),
    .ZN(_208_));
 OAI221_X1 _597_ (.A(\retry_count[2] ),
    .B1(_208_),
    .B2(_146_),
    .C1(_119_),
    .C2(_202_),
    .ZN(_209_));
 OR3_X1 _598_ (.A1(\retry_count[2] ),
    .A2(_208_),
    .A3(_146_),
    .ZN(_210_));
 AOI21_X1 _599_ (.A(_123_),
    .B1(_209_),
    .B2(_210_),
    .ZN(_042_));
 NAND3_X1 _600_ (.A1(\retry_count[0] ),
    .A2(\retry_count[2] ),
    .A3(\retry_count[1] ),
    .ZN(_211_));
 OAI221_X1 _601_ (.A(\retry_count[3] ),
    .B1(_202_),
    .B2(_119_),
    .C1(_146_),
    .C2(_211_),
    .ZN(_212_));
 OR3_X1 _602_ (.A1(\retry_count[3] ),
    .A2(_146_),
    .A3(_211_),
    .ZN(_213_));
 AOI21_X1 _603_ (.A(_123_),
    .B1(_212_),
    .B2(_213_),
    .ZN(_043_));
 BUF_X4 _604_ (.A(_128_),
    .Z(_214_));
 MUX2_X1 _605_ (.A(net1),
    .B(net71),
    .S(_214_),
    .Z(_215_));
 NOR2_X4 _606_ (.A1(_202_),
    .A2(_129_),
    .ZN(_216_));
 BUF_X8 _607_ (.A(_216_),
    .Z(_217_));
 MUX2_X1 _608_ (.A(net173),
    .B(_215_),
    .S(_217_),
    .Z(_218_));
 AND2_X1 _609_ (.A1(_181_),
    .A2(_218_),
    .ZN(_044_));
 MUX2_X1 _610_ (.A(net2),
    .B(net72),
    .S(_214_),
    .Z(_219_));
 MUX2_X1 _611_ (.A(net174),
    .B(_219_),
    .S(_217_),
    .Z(_220_));
 AND2_X1 _612_ (.A1(_181_),
    .A2(_220_),
    .ZN(_045_));
 MUX2_X1 _613_ (.A(net3),
    .B(net73),
    .S(_214_),
    .Z(_221_));
 MUX2_X1 _614_ (.A(net175),
    .B(_221_),
    .S(_217_),
    .Z(_222_));
 AND2_X1 _615_ (.A1(_181_),
    .A2(_222_),
    .ZN(_046_));
 MUX2_X1 _616_ (.A(net4),
    .B(net74),
    .S(_214_),
    .Z(_223_));
 MUX2_X1 _617_ (.A(net176),
    .B(_223_),
    .S(_217_),
    .Z(_224_));
 AND2_X1 _618_ (.A1(_181_),
    .A2(_224_),
    .ZN(_047_));
 MUX2_X1 _619_ (.A(net5),
    .B(net75),
    .S(_214_),
    .Z(_225_));
 MUX2_X1 _620_ (.A(net177),
    .B(_225_),
    .S(_217_),
    .Z(_226_));
 AND2_X1 _621_ (.A1(_181_),
    .A2(_226_),
    .ZN(_048_));
 MUX2_X1 _622_ (.A(net6),
    .B(net76),
    .S(_214_),
    .Z(_227_));
 MUX2_X1 _623_ (.A(net178),
    .B(_227_),
    .S(_217_),
    .Z(_228_));
 AND2_X1 _624_ (.A1(_181_),
    .A2(_228_),
    .ZN(_049_));
 BUF_X2 _625_ (.A(_131_),
    .Z(_229_));
 MUX2_X1 _626_ (.A(net7),
    .B(net77),
    .S(_214_),
    .Z(_230_));
 MUX2_X1 _627_ (.A(net179),
    .B(_230_),
    .S(_217_),
    .Z(_231_));
 AND2_X1 _628_ (.A1(_229_),
    .A2(_231_),
    .ZN(_050_));
 CLKBUF_X3 _629_ (.A(_128_),
    .Z(_232_));
 MUX2_X1 _630_ (.A(net8),
    .B(net78),
    .S(_232_),
    .Z(_233_));
 MUX2_X1 _631_ (.A(net180),
    .B(_233_),
    .S(_217_),
    .Z(_234_));
 AND2_X1 _632_ (.A1(_229_),
    .A2(_234_),
    .ZN(_051_));
 MUX2_X1 _633_ (.A(net9),
    .B(net79),
    .S(_232_),
    .Z(_235_));
 MUX2_X1 _634_ (.A(net181),
    .B(_235_),
    .S(_217_),
    .Z(_236_));
 AND2_X1 _635_ (.A1(_229_),
    .A2(_236_),
    .ZN(_052_));
 MUX2_X1 _636_ (.A(net10),
    .B(net80),
    .S(_232_),
    .Z(_237_));
 MUX2_X1 _637_ (.A(net182),
    .B(_237_),
    .S(_217_),
    .Z(_238_));
 AND2_X1 _638_ (.A1(_229_),
    .A2(_238_),
    .ZN(_053_));
 MUX2_X1 _639_ (.A(net11),
    .B(net81),
    .S(_232_),
    .Z(_239_));
 BUF_X8 _640_ (.A(_216_),
    .Z(_240_));
 MUX2_X1 _641_ (.A(net183),
    .B(_239_),
    .S(_240_),
    .Z(_241_));
 AND2_X1 _642_ (.A1(_229_),
    .A2(_241_),
    .ZN(_054_));
 MUX2_X1 _643_ (.A(net12),
    .B(net82),
    .S(_232_),
    .Z(_242_));
 MUX2_X1 _644_ (.A(net184),
    .B(_242_),
    .S(_240_),
    .Z(_243_));
 AND2_X1 _645_ (.A1(_229_),
    .A2(_243_),
    .ZN(_055_));
 MUX2_X1 _646_ (.A(net13),
    .B(net83),
    .S(_232_),
    .Z(_244_));
 MUX2_X1 _647_ (.A(net185),
    .B(_244_),
    .S(_240_),
    .Z(_245_));
 AND2_X1 _648_ (.A1(_229_),
    .A2(_245_),
    .ZN(_056_));
 MUX2_X1 _649_ (.A(net14),
    .B(net84),
    .S(_232_),
    .Z(_246_));
 MUX2_X1 _650_ (.A(net186),
    .B(_246_),
    .S(_240_),
    .Z(_247_));
 AND2_X1 _651_ (.A1(_229_),
    .A2(_247_),
    .ZN(_057_));
 MUX2_X1 _652_ (.A(net15),
    .B(net85),
    .S(_232_),
    .Z(_248_));
 MUX2_X1 _653_ (.A(net187),
    .B(_248_),
    .S(_240_),
    .Z(_249_));
 AND2_X1 _654_ (.A1(_229_),
    .A2(_249_),
    .ZN(_058_));
 MUX2_X1 _655_ (.A(net16),
    .B(net86),
    .S(_232_),
    .Z(_250_));
 MUX2_X1 _656_ (.A(net188),
    .B(_250_),
    .S(_240_),
    .Z(_251_));
 AND2_X1 _657_ (.A1(_229_),
    .A2(_251_),
    .ZN(_059_));
 BUF_X2 _658_ (.A(_131_),
    .Z(_252_));
 MUX2_X1 _659_ (.A(net17),
    .B(net87),
    .S(_232_),
    .Z(_253_));
 MUX2_X1 _660_ (.A(net189),
    .B(_253_),
    .S(_240_),
    .Z(_254_));
 AND2_X1 _661_ (.A1(_252_),
    .A2(_254_),
    .ZN(_060_));
 CLKBUF_X3 _662_ (.A(_128_),
    .Z(_255_));
 MUX2_X1 _663_ (.A(net18),
    .B(net88),
    .S(_255_),
    .Z(_256_));
 MUX2_X1 _664_ (.A(net190),
    .B(_256_),
    .S(_240_),
    .Z(_257_));
 AND2_X1 _665_ (.A1(_252_),
    .A2(_257_),
    .ZN(_061_));
 MUX2_X1 _666_ (.A(net19),
    .B(net89),
    .S(_255_),
    .Z(_258_));
 MUX2_X1 _667_ (.A(net191),
    .B(_258_),
    .S(_240_),
    .Z(_259_));
 AND2_X1 _668_ (.A1(_252_),
    .A2(_259_),
    .ZN(_062_));
 MUX2_X1 _669_ (.A(net20),
    .B(net90),
    .S(_255_),
    .Z(_260_));
 MUX2_X1 _670_ (.A(net192),
    .B(_260_),
    .S(_240_),
    .Z(_261_));
 AND2_X1 _671_ (.A1(_252_),
    .A2(_261_),
    .ZN(_063_));
 MUX2_X1 _672_ (.A(net21),
    .B(net91),
    .S(_255_),
    .Z(_262_));
 BUF_X8 _673_ (.A(_216_),
    .Z(_263_));
 MUX2_X1 _674_ (.A(net193),
    .B(_262_),
    .S(_263_),
    .Z(_264_));
 AND2_X1 _675_ (.A1(_252_),
    .A2(_264_),
    .ZN(_064_));
 MUX2_X1 _676_ (.A(net22),
    .B(net92),
    .S(_255_),
    .Z(_265_));
 MUX2_X1 _677_ (.A(net194),
    .B(_265_),
    .S(_263_),
    .Z(_266_));
 AND2_X1 _678_ (.A1(_252_),
    .A2(_266_),
    .ZN(_065_));
 MUX2_X1 _679_ (.A(net23),
    .B(net93),
    .S(_255_),
    .Z(_267_));
 MUX2_X1 _680_ (.A(net195),
    .B(_267_),
    .S(_263_),
    .Z(_268_));
 AND2_X1 _681_ (.A1(_252_),
    .A2(_268_),
    .ZN(_066_));
 MUX2_X1 _682_ (.A(net24),
    .B(net94),
    .S(_255_),
    .Z(_269_));
 MUX2_X1 _683_ (.A(net196),
    .B(_269_),
    .S(_263_),
    .Z(_270_));
 AND2_X1 _684_ (.A1(_252_),
    .A2(_270_),
    .ZN(_067_));
 MUX2_X1 _685_ (.A(net25),
    .B(net95),
    .S(_255_),
    .Z(_271_));
 MUX2_X1 _686_ (.A(net197),
    .B(_271_),
    .S(_263_),
    .Z(_272_));
 AND2_X1 _687_ (.A1(_252_),
    .A2(_272_),
    .ZN(_068_));
 MUX2_X1 _688_ (.A(net26),
    .B(net96),
    .S(_255_),
    .Z(_273_));
 MUX2_X1 _689_ (.A(net198),
    .B(_273_),
    .S(_263_),
    .Z(_274_));
 AND2_X1 _690_ (.A1(_252_),
    .A2(_274_),
    .ZN(_069_));
 BUF_X2 _691_ (.A(_122_),
    .Z(_275_));
 MUX2_X1 _692_ (.A(net27),
    .B(net97),
    .S(_255_),
    .Z(_276_));
 MUX2_X1 _693_ (.A(net199),
    .B(_276_),
    .S(_263_),
    .Z(_277_));
 AND2_X1 _694_ (.A1(_275_),
    .A2(_277_),
    .ZN(_070_));
 MUX2_X1 _695_ (.A(net28),
    .B(net98),
    .S(_188_),
    .Z(_278_));
 MUX2_X1 _696_ (.A(net200),
    .B(_278_),
    .S(_263_),
    .Z(_279_));
 AND2_X1 _697_ (.A1(_275_),
    .A2(_279_),
    .ZN(_071_));
 MUX2_X1 _698_ (.A(net29),
    .B(net99),
    .S(_188_),
    .Z(_280_));
 MUX2_X1 _699_ (.A(net201),
    .B(_280_),
    .S(_263_),
    .Z(_281_));
 AND2_X1 _700_ (.A1(_275_),
    .A2(_281_),
    .ZN(_072_));
 MUX2_X1 _701_ (.A(net30),
    .B(net100),
    .S(_188_),
    .Z(_282_));
 MUX2_X1 _702_ (.A(net202),
    .B(_282_),
    .S(_263_),
    .Z(_283_));
 AND2_X1 _703_ (.A1(_275_),
    .A2(_283_),
    .ZN(_073_));
 MUX2_X1 _704_ (.A(net31),
    .B(net101),
    .S(_188_),
    .Z(_284_));
 MUX2_X1 _705_ (.A(net203),
    .B(_284_),
    .S(_216_),
    .Z(_285_));
 AND2_X1 _706_ (.A1(_275_),
    .A2(_285_),
    .ZN(_074_));
 MUX2_X1 _707_ (.A(net32),
    .B(net102),
    .S(_188_),
    .Z(_286_));
 MUX2_X1 _708_ (.A(net204),
    .B(_286_),
    .S(_216_),
    .Z(_287_));
 AND2_X1 _709_ (.A1(_275_),
    .A2(_287_),
    .ZN(_075_));
 NOR3_X1 _710_ (.A1(_127_),
    .A2(_214_),
    .A3(_119_),
    .ZN(_288_));
 MUX2_X1 _711_ (.A(_193_),
    .B(_137_),
    .S(_119_),
    .Z(_289_));
 AOI221_X2 _712_ (.A(_123_),
    .B1(_004_),
    .B2(_288_),
    .C1(_289_),
    .C2(_136_),
    .ZN(_076_));
 MUX2_X1 _713_ (.A(net103),
    .B(net206),
    .S(_141_),
    .Z(_290_));
 AND2_X1 _714_ (.A1(_275_),
    .A2(_290_),
    .ZN(_077_));
 MUX2_X1 _715_ (.A(net104),
    .B(net207),
    .S(_141_),
    .Z(_291_));
 AND2_X1 _716_ (.A1(_275_),
    .A2(_291_),
    .ZN(_078_));
 MUX2_X1 _717_ (.A(net105),
    .B(net208),
    .S(_141_),
    .Z(_292_));
 AND2_X1 _718_ (.A1(_275_),
    .A2(_292_),
    .ZN(_079_));
 MUX2_X1 _719_ (.A(net106),
    .B(net209),
    .S(_141_),
    .Z(_293_));
 AND2_X1 _720_ (.A1(_275_),
    .A2(_293_),
    .ZN(_080_));
 CLKBUF_X2 _721_ (.A(_122_),
    .Z(_294_));
 MUX2_X1 _722_ (.A(net107),
    .B(net210),
    .S(_141_),
    .Z(_295_));
 AND2_X1 _723_ (.A1(_294_),
    .A2(_295_),
    .ZN(_081_));
 MUX2_X1 _724_ (.A(net108),
    .B(net211),
    .S(_141_),
    .Z(_296_));
 AND2_X1 _725_ (.A1(_294_),
    .A2(_296_),
    .ZN(_082_));
 MUX2_X1 _726_ (.A(net109),
    .B(net212),
    .S(_141_),
    .Z(_297_));
 AND2_X1 _727_ (.A1(_294_),
    .A2(_297_),
    .ZN(_083_));
 MUX2_X1 _728_ (.A(net110),
    .B(net213),
    .S(_141_),
    .Z(_298_));
 AND2_X1 _729_ (.A1(_294_),
    .A2(_298_),
    .ZN(_084_));
 MUX2_X1 _730_ (.A(net111),
    .B(net214),
    .S(_141_),
    .Z(_299_));
 AND2_X1 _731_ (.A1(_294_),
    .A2(_299_),
    .ZN(_085_));
 CLKBUF_X3 _732_ (.A(_140_),
    .Z(_300_));
 MUX2_X1 _733_ (.A(net112),
    .B(net215),
    .S(_300_),
    .Z(_301_));
 AND2_X1 _734_ (.A1(_294_),
    .A2(_301_),
    .ZN(_086_));
 MUX2_X1 _735_ (.A(net113),
    .B(net216),
    .S(_300_),
    .Z(_302_));
 AND2_X1 _736_ (.A1(_294_),
    .A2(_302_),
    .ZN(_087_));
 MUX2_X1 _737_ (.A(net114),
    .B(net217),
    .S(_300_),
    .Z(_303_));
 AND2_X1 _738_ (.A1(_294_),
    .A2(_303_),
    .ZN(_088_));
 MUX2_X1 _739_ (.A(net115),
    .B(net218),
    .S(_300_),
    .Z(_304_));
 AND2_X1 _740_ (.A1(_294_),
    .A2(_304_),
    .ZN(_089_));
 MUX2_X1 _741_ (.A(net116),
    .B(net219),
    .S(_300_),
    .Z(_305_));
 AND2_X1 _742_ (.A1(_294_),
    .A2(_305_),
    .ZN(_090_));
 CLKBUF_X2 _743_ (.A(_122_),
    .Z(_306_));
 MUX2_X1 _744_ (.A(net117),
    .B(net220),
    .S(_300_),
    .Z(_307_));
 AND2_X1 _745_ (.A1(_306_),
    .A2(_307_),
    .ZN(_091_));
 MUX2_X1 _746_ (.A(net118),
    .B(net221),
    .S(_300_),
    .Z(_308_));
 AND2_X1 _747_ (.A1(_306_),
    .A2(_308_),
    .ZN(_092_));
 MUX2_X1 _748_ (.A(net119),
    .B(net222),
    .S(_300_),
    .Z(_309_));
 AND2_X1 _749_ (.A1(_306_),
    .A2(_309_),
    .ZN(_093_));
 MUX2_X1 _750_ (.A(net120),
    .B(net223),
    .S(_300_),
    .Z(_310_));
 AND2_X1 _751_ (.A1(_306_),
    .A2(_310_),
    .ZN(_094_));
 MUX2_X1 _752_ (.A(net121),
    .B(net224),
    .S(_300_),
    .Z(_311_));
 AND2_X1 _753_ (.A1(_306_),
    .A2(_311_),
    .ZN(_095_));
 CLKBUF_X3 _754_ (.A(_140_),
    .Z(_312_));
 MUX2_X1 _755_ (.A(net122),
    .B(net225),
    .S(_312_),
    .Z(_313_));
 AND2_X1 _756_ (.A1(_306_),
    .A2(_313_),
    .ZN(_096_));
 MUX2_X1 _757_ (.A(net123),
    .B(net226),
    .S(_312_),
    .Z(_314_));
 AND2_X1 _758_ (.A1(_306_),
    .A2(_314_),
    .ZN(_097_));
 MUX2_X1 _759_ (.A(net124),
    .B(net227),
    .S(_312_),
    .Z(_315_));
 AND2_X1 _760_ (.A1(_306_),
    .A2(_315_),
    .ZN(_098_));
 MUX2_X1 _761_ (.A(net125),
    .B(net228),
    .S(_312_),
    .Z(_316_));
 AND2_X1 _762_ (.A1(_306_),
    .A2(_316_),
    .ZN(_099_));
 MUX2_X1 _763_ (.A(net126),
    .B(net229),
    .S(_312_),
    .Z(_317_));
 AND2_X1 _764_ (.A1(_306_),
    .A2(_317_),
    .ZN(_100_));
 BUF_X2 _765_ (.A(_122_),
    .Z(_318_));
 MUX2_X1 _766_ (.A(net127),
    .B(net230),
    .S(_312_),
    .Z(_319_));
 AND2_X1 _767_ (.A1(_318_),
    .A2(_319_),
    .ZN(_101_));
 MUX2_X1 _768_ (.A(net128),
    .B(net231),
    .S(_312_),
    .Z(_320_));
 AND2_X1 _769_ (.A1(_318_),
    .A2(_320_),
    .ZN(_102_));
 MUX2_X1 _770_ (.A(net129),
    .B(net232),
    .S(_312_),
    .Z(_321_));
 AND2_X1 _771_ (.A1(_318_),
    .A2(_321_),
    .ZN(_103_));
 MUX2_X1 _772_ (.A(net130),
    .B(net233),
    .S(_312_),
    .Z(_322_));
 AND2_X1 _773_ (.A1(_318_),
    .A2(_322_),
    .ZN(_104_));
 MUX2_X1 _774_ (.A(net131),
    .B(net234),
    .S(_312_),
    .Z(_323_));
 AND2_X1 _775_ (.A1(_318_),
    .A2(_323_),
    .ZN(_105_));
 MUX2_X1 _776_ (.A(net132),
    .B(net235),
    .S(_140_),
    .Z(_324_));
 AND2_X1 _777_ (.A1(_318_),
    .A2(_324_),
    .ZN(_106_));
 MUX2_X1 _778_ (.A(net133),
    .B(net236),
    .S(_140_),
    .Z(_325_));
 AND2_X1 _779_ (.A1(_318_),
    .A2(_325_),
    .ZN(_107_));
 MUX2_X1 _780_ (.A(net134),
    .B(net237),
    .S(_140_),
    .Z(_326_));
 AND2_X1 _781_ (.A1(_318_),
    .A2(_326_),
    .ZN(_108_));
 MUX2_X1 _782_ (.A(net33),
    .B(net135),
    .S(_188_),
    .Z(_327_));
 MUX2_X1 _783_ (.A(net238),
    .B(_327_),
    .S(_216_),
    .Z(_328_));
 AND2_X1 _784_ (.A1(_318_),
    .A2(_328_),
    .ZN(_109_));
 MUX2_X1 _785_ (.A(net34),
    .B(net136),
    .S(_188_),
    .Z(_329_));
 MUX2_X1 _786_ (.A(net239),
    .B(_329_),
    .S(_216_),
    .Z(_330_));
 AND2_X1 _787_ (.A1(_318_),
    .A2(_330_),
    .ZN(_110_));
 MUX2_X1 _788_ (.A(net35),
    .B(net137),
    .S(_188_),
    .Z(_331_));
 MUX2_X1 _789_ (.A(net240),
    .B(_331_),
    .S(_216_),
    .Z(_332_));
 AND2_X1 _790_ (.A1(_131_),
    .A2(_332_),
    .ZN(_111_));
 MUX2_X1 _791_ (.A(net36),
    .B(net138),
    .S(_188_),
    .Z(_333_));
 MUX2_X1 _792_ (.A(net241),
    .B(_333_),
    .S(_216_),
    .Z(_334_));
 AND2_X1 _793_ (.A1(_131_),
    .A2(_334_),
    .ZN(_112_));
 OAI21_X1 _794_ (.A(net243),
    .B1(_202_),
    .B2(_187_),
    .ZN(_335_));
 OAI21_X1 _795_ (.A(_335_),
    .B1(_202_),
    .B2(_133_),
    .ZN(_336_));
 AND2_X1 _796_ (.A1(_131_),
    .A2(_336_),
    .ZN(_113_));
 AND2_X1 _797_ (.A1(_120_),
    .A2(_117_),
    .ZN(_337_));
 OAI21_X1 _798_ (.A(_131_),
    .B1(net244),
    .B2(_337_),
    .ZN(_338_));
 NAND2_X1 _799_ (.A1(_214_),
    .A2(_143_),
    .ZN(_339_));
 OAI21_X1 _800_ (.A(_339_),
    .B1(net244),
    .B2(_214_),
    .ZN(_340_));
 AOI21_X1 _801_ (.A(_338_),
    .B1(_340_),
    .B2(_126_),
    .ZN(_114_));
 INV_X1 _802_ (.A(net245),
    .ZN(_341_));
 AOI21_X1 _803_ (.A(_337_),
    .B1(_126_),
    .B2(_133_),
    .ZN(_342_));
 OAI21_X1 _804_ (.A(_124_),
    .B1(_142_),
    .B2(_135_),
    .ZN(_343_));
 NAND2_X1 _805_ (.A1(_117_),
    .A2(_145_),
    .ZN(_344_));
 NAND3_X1 _806_ (.A1(_191_),
    .A2(_143_),
    .A3(_004_),
    .ZN(_345_));
 NAND4_X1 _807_ (.A1(_342_),
    .A2(_343_),
    .A3(_344_),
    .A4(_345_),
    .ZN(_346_));
 AOI21_X1 _808_ (.A(_117_),
    .B1(_126_),
    .B2(_133_),
    .ZN(_347_));
 NOR2_X1 _809_ (.A1(_124_),
    .A2(_194_),
    .ZN(_348_));
 AOI221_X1 _810_ (.A(_123_),
    .B1(_341_),
    .B2(_346_),
    .C1(_347_),
    .C2(_348_),
    .ZN(_115_));
 HA_X1 _811_ (.A(\retry_count[0] ),
    .B(\retry_count[1] ),
    .CO(_461_),
    .S(_462_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _813_ (.A(net205),
    .Z(net242));
 BUF_X1 _814_ (.A(net246),
    .Z(wb_tgd_o));
 DFF_X1 \read_data[0]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_4_10_0_clk),
    .Q(net139),
    .QN(_457_));
 DFF_X1 \read_data[10]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_4_10_0_clk),
    .Q(net140),
    .QN(_456_));
 DFF_X1 \read_data[11]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_4_8_0_clk),
    .Q(net141),
    .QN(_455_));
 DFF_X1 \read_data[12]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_4_8_0_clk),
    .Q(net142),
    .QN(_454_));
 DFF_X1 \read_data[13]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_4_10_0_clk),
    .Q(net143),
    .QN(_453_));
 DFF_X1 \read_data[14]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_4_8_0_clk),
    .Q(net144),
    .QN(_452_));
 DFF_X1 \read_data[15]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_4_8_0_clk),
    .Q(net145),
    .QN(_451_));
 DFF_X1 \read_data[16]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_4_10_0_clk),
    .Q(net146),
    .QN(_450_));
 DFF_X1 \read_data[17]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_4_10_0_clk),
    .Q(net147),
    .QN(_449_));
 DFF_X1 \read_data[18]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_4_9_0_clk),
    .Q(net148),
    .QN(_448_));
 DFF_X1 \read_data[19]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_4_10_0_clk),
    .Q(net149),
    .QN(_447_));
 DFF_X1 \read_data[1]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_4_9_0_clk),
    .Q(net150),
    .QN(_446_));
 DFF_X1 \read_data[20]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_4_11_0_clk),
    .Q(net151),
    .QN(_445_));
 DFF_X1 \read_data[21]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_4_11_0_clk),
    .Q(net152),
    .QN(_444_));
 DFF_X1 \read_data[22]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_4_11_0_clk),
    .Q(net153),
    .QN(_443_));
 DFF_X1 \read_data[23]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_4_11_0_clk),
    .Q(net154),
    .QN(_442_));
 DFF_X1 \read_data[24]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_4_11_0_clk),
    .Q(net155),
    .QN(_441_));
 DFF_X1 \read_data[25]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_4_10_0_clk),
    .Q(net156),
    .QN(_440_));
 DFF_X1 \read_data[26]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_4_14_0_clk),
    .Q(net157),
    .QN(_439_));
 DFF_X1 \read_data[27]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_4_15_0_clk),
    .Q(net158),
    .QN(_438_));
 DFF_X1 \read_data[28]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_4_15_0_clk),
    .Q(net159),
    .QN(_437_));
 DFF_X1 \read_data[29]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_4_15_0_clk),
    .Q(net160),
    .QN(_436_));
 DFF_X1 \read_data[2]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_4_15_0_clk),
    .Q(net161),
    .QN(_435_));
 DFF_X1 \read_data[30]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_4_14_0_clk),
    .Q(net162),
    .QN(_434_));
 DFF_X1 \read_data[31]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_4_15_0_clk),
    .Q(net163),
    .QN(_433_));
 DFF_X1 \read_data[3]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_4_15_0_clk),
    .Q(net164),
    .QN(_432_));
 DFF_X1 \read_data[4]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_4_14_0_clk),
    .Q(net165),
    .QN(_431_));
 DFF_X1 \read_data[5]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_4_15_0_clk),
    .Q(net166),
    .QN(_430_));
 DFF_X1 \read_data[6]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_4_14_0_clk),
    .Q(net167),
    .QN(_429_));
 DFF_X1 \read_data[7]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_4_14_0_clk),
    .Q(net168),
    .QN(_428_));
 DFF_X1 \read_data[8]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_4_11_0_clk),
    .Q(net169),
    .QN(_427_));
 DFF_X1 \read_data[9]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_4_14_0_clk),
    .Q(net170),
    .QN(_426_));
 DFF_X1 \read_done$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_4_9_0_clk),
    .Q(net171),
    .QN(_425_));
 DFF_X1 \read_err$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_4_12_0_clk),
    .Q(net172),
    .QN(_424_));
 DFF_X1 \retry_count[0]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_4_3_0_clk),
    .Q(\retry_count[0] ),
    .QN(_423_));
 DFF_X1 \retry_count[1]$_SDFFE_PN0P_  (.D(_041_),
    .CK(clknet_4_3_0_clk),
    .Q(\retry_count[1] ),
    .QN(_422_));
 DFF_X1 \retry_count[2]$_SDFFE_PN0P_  (.D(_042_),
    .CK(clknet_4_3_0_clk),
    .Q(\retry_count[2] ),
    .QN(_421_));
 DFF_X1 \retry_count[3]$_SDFFE_PN0P_  (.D(_043_),
    .CK(clknet_4_3_0_clk),
    .Q(\retry_count[3] ),
    .QN(_458_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_4_3_0_clk),
    .Q(\state[0] ),
    .QN(_005_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_002_),
    .CK(clknet_4_9_0_clk),
    .Q(\state[1] ),
    .QN(_459_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_003_),
    .CK(clknet_4_8_0_clk),
    .Q(\state[2] ),
    .QN(_460_));
 DFF_X2 \state[3]$_DFF_P_  (.D(_000_),
    .CK(clknet_4_3_0_clk),
    .Q(\state[3] ),
    .QN(_004_));
 DFF_X1 \wb_adr_o[0]$_SDFFE_PN0P_  (.D(_044_),
    .CK(clknet_4_15_0_clk),
    .Q(net173),
    .QN(_420_));
 DFF_X1 \wb_adr_o[10]$_SDFFE_PN0P_  (.D(_045_),
    .CK(clknet_4_12_0_clk),
    .Q(net174),
    .QN(_419_));
 DFF_X1 \wb_adr_o[11]$_SDFFE_PN0P_  (.D(_046_),
    .CK(clknet_4_12_0_clk),
    .Q(net175),
    .QN(_418_));
 DFF_X1 \wb_adr_o[12]$_SDFFE_PN0P_  (.D(_047_),
    .CK(clknet_4_14_0_clk),
    .Q(net176),
    .QN(_417_));
 DFF_X1 \wb_adr_o[13]$_SDFFE_PN0P_  (.D(_048_),
    .CK(clknet_4_14_0_clk),
    .Q(net177),
    .QN(_416_));
 DFF_X1 \wb_adr_o[14]$_SDFFE_PN0P_  (.D(_049_),
    .CK(clknet_4_13_0_clk),
    .Q(net178),
    .QN(_415_));
 DFF_X1 \wb_adr_o[15]$_SDFFE_PN0P_  (.D(_050_),
    .CK(clknet_4_15_0_clk),
    .Q(net179),
    .QN(_414_));
 DFF_X1 \wb_adr_o[16]$_SDFFE_PN0P_  (.D(_051_),
    .CK(clknet_4_13_0_clk),
    .Q(net180),
    .QN(_413_));
 DFF_X1 \wb_adr_o[17]$_SDFFE_PN0P_  (.D(_052_),
    .CK(clknet_4_13_0_clk),
    .Q(net181),
    .QN(_412_));
 DFF_X1 \wb_adr_o[18]$_SDFFE_PN0P_  (.D(_053_),
    .CK(clknet_4_15_0_clk),
    .Q(net182),
    .QN(_411_));
 DFF_X1 \wb_adr_o[19]$_SDFFE_PN0P_  (.D(_054_),
    .CK(clknet_4_7_0_clk),
    .Q(net183),
    .QN(_410_));
 DFF_X1 \wb_adr_o[1]$_SDFFE_PN0P_  (.D(_055_),
    .CK(clknet_4_13_0_clk),
    .Q(net184),
    .QN(_409_));
 DFF_X1 \wb_adr_o[20]$_SDFFE_PN0P_  (.D(_056_),
    .CK(clknet_4_12_0_clk),
    .Q(net185),
    .QN(_408_));
 DFF_X1 \wb_adr_o[21]$_SDFFE_PN0P_  (.D(_057_),
    .CK(clknet_4_13_0_clk),
    .Q(net186),
    .QN(_407_));
 DFF_X1 \wb_adr_o[22]$_SDFFE_PN0P_  (.D(_058_),
    .CK(clknet_4_13_0_clk),
    .Q(net187),
    .QN(_406_));
 DFF_X1 \wb_adr_o[23]$_SDFFE_PN0P_  (.D(_059_),
    .CK(clknet_4_13_0_clk),
    .Q(net188),
    .QN(_405_));
 DFF_X1 \wb_adr_o[24]$_SDFFE_PN0P_  (.D(_060_),
    .CK(clknet_4_7_0_clk),
    .Q(net189),
    .QN(_404_));
 DFF_X1 \wb_adr_o[25]$_SDFFE_PN0P_  (.D(_061_),
    .CK(clknet_4_7_0_clk),
    .Q(net190),
    .QN(_403_));
 DFF_X1 \wb_adr_o[26]$_SDFFE_PN0P_  (.D(_062_),
    .CK(clknet_4_6_0_clk),
    .Q(net191),
    .QN(_402_));
 DFF_X1 \wb_adr_o[27]$_SDFFE_PN0P_  (.D(_063_),
    .CK(clknet_4_7_0_clk),
    .Q(net192),
    .QN(_401_));
 DFF_X1 \wb_adr_o[28]$_SDFFE_PN0P_  (.D(_064_),
    .CK(clknet_4_5_0_clk),
    .Q(net193),
    .QN(_400_));
 DFF_X1 \wb_adr_o[29]$_SDFFE_PN0P_  (.D(_065_),
    .CK(clknet_4_6_0_clk),
    .Q(net194),
    .QN(_399_));
 DFF_X1 \wb_adr_o[2]$_SDFFE_PN0P_  (.D(_066_),
    .CK(clknet_4_5_0_clk),
    .Q(net195),
    .QN(_398_));
 DFF_X1 \wb_adr_o[30]$_SDFFE_PN0P_  (.D(_067_),
    .CK(clknet_4_5_0_clk),
    .Q(net196),
    .QN(_397_));
 DFF_X1 \wb_adr_o[31]$_SDFFE_PN0P_  (.D(_068_),
    .CK(clknet_4_5_0_clk),
    .Q(net197),
    .QN(_396_));
 DFF_X1 \wb_adr_o[3]$_SDFFE_PN0P_  (.D(_069_),
    .CK(clknet_4_5_0_clk),
    .Q(net198),
    .QN(_395_));
 DFF_X1 \wb_adr_o[4]$_SDFFE_PN0P_  (.D(_070_),
    .CK(clknet_4_5_0_clk),
    .Q(net199),
    .QN(_394_));
 DFF_X1 \wb_adr_o[5]$_SDFFE_PN0P_  (.D(_071_),
    .CK(clknet_4_5_0_clk),
    .Q(net200),
    .QN(_393_));
 DFF_X1 \wb_adr_o[6]$_SDFFE_PN0P_  (.D(_072_),
    .CK(clknet_4_6_0_clk),
    .Q(net201),
    .QN(_392_));
 DFF_X1 \wb_adr_o[7]$_SDFFE_PN0P_  (.D(_073_),
    .CK(clknet_4_5_0_clk),
    .Q(net202),
    .QN(_391_));
 DFF_X1 \wb_adr_o[8]$_SDFFE_PN0P_  (.D(_074_),
    .CK(clknet_4_4_0_clk),
    .Q(net203),
    .QN(_390_));
 DFF_X1 \wb_adr_o[9]$_SDFFE_PN0P_  (.D(_075_),
    .CK(clknet_4_6_0_clk),
    .Q(net204),
    .QN(_389_));
 DFF_X1 \wb_cyc_o$_SDFF_PN0_  (.D(_076_),
    .CK(clknet_4_12_0_clk),
    .Q(net205),
    .QN(_388_));
 DFF_X1 \wb_dat_o[0]$_SDFFE_PN0P_  (.D(_077_),
    .CK(clknet_4_5_0_clk),
    .Q(net206),
    .QN(_387_));
 DFF_X1 \wb_dat_o[10]$_SDFFE_PN0P_  (.D(_078_),
    .CK(clknet_4_5_0_clk),
    .Q(net207),
    .QN(_386_));
 DFF_X1 \wb_dat_o[11]$_SDFFE_PN0P_  (.D(_079_),
    .CK(clknet_4_4_0_clk),
    .Q(net208),
    .QN(_385_));
 DFF_X1 \wb_dat_o[12]$_SDFFE_PN0P_  (.D(_080_),
    .CK(clknet_4_4_0_clk),
    .Q(net209),
    .QN(_384_));
 DFF_X1 \wb_dat_o[13]$_SDFFE_PN0P_  (.D(_081_),
    .CK(clknet_4_1_0_clk),
    .Q(net210),
    .QN(_383_));
 DFF_X1 \wb_dat_o[14]$_SDFFE_PN0P_  (.D(_082_),
    .CK(clknet_4_4_0_clk),
    .Q(net211),
    .QN(_382_));
 DFF_X1 \wb_dat_o[15]$_SDFFE_PN0P_  (.D(_083_),
    .CK(clknet_4_1_0_clk),
    .Q(net212),
    .QN(_381_));
 DFF_X1 \wb_dat_o[16]$_SDFFE_PN0P_  (.D(_084_),
    .CK(clknet_4_1_0_clk),
    .Q(net213),
    .QN(_380_));
 DFF_X1 \wb_dat_o[17]$_SDFFE_PN0P_  (.D(_085_),
    .CK(clknet_4_4_0_clk),
    .Q(net214),
    .QN(_379_));
 DFF_X1 \wb_dat_o[18]$_SDFFE_PN0P_  (.D(_086_),
    .CK(clknet_4_0_0_clk),
    .Q(net215),
    .QN(_378_));
 DFF_X1 \wb_dat_o[19]$_SDFFE_PN0P_  (.D(_087_),
    .CK(clknet_4_1_0_clk),
    .Q(net216),
    .QN(_377_));
 DFF_X1 \wb_dat_o[1]$_SDFFE_PN0P_  (.D(_088_),
    .CK(clknet_4_1_0_clk),
    .Q(net217),
    .QN(_376_));
 DFF_X1 \wb_dat_o[20]$_SDFFE_PN0P_  (.D(_089_),
    .CK(clknet_4_1_0_clk),
    .Q(net218),
    .QN(_375_));
 DFF_X1 \wb_dat_o[21]$_SDFFE_PN0P_  (.D(_090_),
    .CK(clknet_4_1_0_clk),
    .Q(net219),
    .QN(_374_));
 DFF_X1 \wb_dat_o[22]$_SDFFE_PN0P_  (.D(_091_),
    .CK(clknet_4_2_0_clk),
    .Q(net220),
    .QN(_373_));
 DFF_X1 \wb_dat_o[23]$_SDFFE_PN0P_  (.D(_092_),
    .CK(clknet_4_0_0_clk),
    .Q(net221),
    .QN(_372_));
 DFF_X1 \wb_dat_o[24]$_SDFFE_PN0P_  (.D(_093_),
    .CK(clknet_4_0_0_clk),
    .Q(net222),
    .QN(_371_));
 DFF_X1 \wb_dat_o[25]$_SDFFE_PN0P_  (.D(_094_),
    .CK(clknet_4_0_0_clk),
    .Q(net223),
    .QN(_370_));
 DFF_X1 \wb_dat_o[26]$_SDFFE_PN0P_  (.D(_095_),
    .CK(clknet_4_1_0_clk),
    .Q(net224),
    .QN(_369_));
 DFF_X1 \wb_dat_o[27]$_SDFFE_PN0P_  (.D(_096_),
    .CK(clknet_4_0_0_clk),
    .Q(net225),
    .QN(_368_));
 DFF_X1 \wb_dat_o[28]$_SDFFE_PN0P_  (.D(_097_),
    .CK(clknet_4_0_0_clk),
    .Q(net226),
    .QN(_367_));
 DFF_X1 \wb_dat_o[29]$_SDFFE_PN0P_  (.D(_098_),
    .CK(clknet_4_0_0_clk),
    .Q(net227),
    .QN(_366_));
 DFF_X1 \wb_dat_o[2]$_SDFFE_PN0P_  (.D(_099_),
    .CK(clknet_4_0_0_clk),
    .Q(net228),
    .QN(_365_));
 DFF_X1 \wb_dat_o[30]$_SDFFE_PN0P_  (.D(_100_),
    .CK(clknet_4_0_0_clk),
    .Q(net229),
    .QN(_364_));
 DFF_X1 \wb_dat_o[31]$_SDFFE_PN0P_  (.D(_101_),
    .CK(clknet_4_2_0_clk),
    .Q(net230),
    .QN(_363_));
 DFF_X1 \wb_dat_o[3]$_SDFFE_PN0P_  (.D(_102_),
    .CK(clknet_4_2_0_clk),
    .Q(net231),
    .QN(_362_));
 DFF_X1 \wb_dat_o[4]$_SDFFE_PN0P_  (.D(_103_),
    .CK(clknet_4_2_0_clk),
    .Q(net232),
    .QN(_361_));
 DFF_X1 \wb_dat_o[5]$_SDFFE_PN0P_  (.D(_104_),
    .CK(clknet_4_2_0_clk),
    .Q(net233),
    .QN(_360_));
 DFF_X1 \wb_dat_o[6]$_SDFFE_PN0P_  (.D(_105_),
    .CK(clknet_4_2_0_clk),
    .Q(net234),
    .QN(_359_));
 DFF_X1 \wb_dat_o[7]$_SDFFE_PN0P_  (.D(_106_),
    .CK(clknet_4_2_0_clk),
    .Q(net235),
    .QN(_358_));
 DFF_X1 \wb_dat_o[8]$_SDFFE_PN0P_  (.D(_107_),
    .CK(clknet_4_1_0_clk),
    .Q(net236),
    .QN(_357_));
 DFF_X1 \wb_dat_o[9]$_SDFFE_PN0P_  (.D(_108_),
    .CK(clknet_4_2_0_clk),
    .Q(net237),
    .QN(_356_));
 DFF_X1 \wb_sel_o[0]$_SDFFE_PN0P_  (.D(_109_),
    .CK(clknet_4_4_0_clk),
    .Q(net238),
    .QN(_355_));
 DFF_X1 \wb_sel_o[1]$_SDFFE_PN0P_  (.D(_110_),
    .CK(clknet_4_4_0_clk),
    .Q(net239),
    .QN(_354_));
 DFF_X1 \wb_sel_o[2]$_SDFFE_PN0P_  (.D(_111_),
    .CK(clknet_4_7_0_clk),
    .Q(net240),
    .QN(_353_));
 DFF_X1 \wb_sel_o[3]$_SDFFE_PN0P_  (.D(_112_),
    .CK(clknet_4_7_0_clk),
    .Q(net241),
    .QN(_352_));
 DFF_X2 \wb_we_o$_SDFFE_PN0P_  (.D(_113_),
    .CK(clknet_4_12_0_clk),
    .Q(net243),
    .QN(_351_));
 DFF_X1 \write_done$_SDFFE_PN0P_  (.D(_114_),
    .CK(clknet_4_11_0_clk),
    .Q(net244),
    .QN(_350_));
 DFF_X1 \write_err$_SDFFE_PN0P_  (.D(_115_),
    .CK(clknet_4_8_0_clk),
    .Q(net245),
    .QN(_349_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_63 ();
 BUF_X1 input1 (.A(read_addr[0]),
    .Z(net1));
 BUF_X1 input2 (.A(read_addr[10]),
    .Z(net2));
 BUF_X1 input3 (.A(read_addr[11]),
    .Z(net3));
 BUF_X1 input4 (.A(read_addr[12]),
    .Z(net4));
 BUF_X1 input5 (.A(read_addr[13]),
    .Z(net5));
 BUF_X1 input6 (.A(read_addr[14]),
    .Z(net6));
 BUF_X1 input7 (.A(read_addr[15]),
    .Z(net7));
 BUF_X1 input8 (.A(read_addr[16]),
    .Z(net8));
 BUF_X1 input9 (.A(read_addr[17]),
    .Z(net9));
 BUF_X1 input10 (.A(read_addr[18]),
    .Z(net10));
 BUF_X1 input11 (.A(read_addr[19]),
    .Z(net11));
 BUF_X1 input12 (.A(read_addr[1]),
    .Z(net12));
 BUF_X1 input13 (.A(read_addr[20]),
    .Z(net13));
 BUF_X1 input14 (.A(read_addr[21]),
    .Z(net14));
 BUF_X1 input15 (.A(read_addr[22]),
    .Z(net15));
 BUF_X1 input16 (.A(read_addr[23]),
    .Z(net16));
 BUF_X1 input17 (.A(read_addr[24]),
    .Z(net17));
 BUF_X1 input18 (.A(read_addr[25]),
    .Z(net18));
 BUF_X1 input19 (.A(read_addr[26]),
    .Z(net19));
 BUF_X1 input20 (.A(read_addr[27]),
    .Z(net20));
 BUF_X1 input21 (.A(read_addr[28]),
    .Z(net21));
 BUF_X1 input22 (.A(read_addr[29]),
    .Z(net22));
 BUF_X1 input23 (.A(read_addr[2]),
    .Z(net23));
 BUF_X1 input24 (.A(read_addr[30]),
    .Z(net24));
 BUF_X1 input25 (.A(read_addr[31]),
    .Z(net25));
 BUF_X1 input26 (.A(read_addr[3]),
    .Z(net26));
 BUF_X1 input27 (.A(read_addr[4]),
    .Z(net27));
 BUF_X1 input28 (.A(read_addr[5]),
    .Z(net28));
 BUF_X1 input29 (.A(read_addr[6]),
    .Z(net29));
 BUF_X1 input30 (.A(read_addr[7]),
    .Z(net30));
 BUF_X1 input31 (.A(read_addr[8]),
    .Z(net31));
 BUF_X1 input32 (.A(read_addr[9]),
    .Z(net32));
 BUF_X1 input33 (.A(read_sel[0]),
    .Z(net33));
 BUF_X1 input34 (.A(read_sel[1]),
    .Z(net34));
 BUF_X1 input35 (.A(read_sel[2]),
    .Z(net35));
 BUF_X1 input36 (.A(read_sel[3]),
    .Z(net36));
 BUF_X1 input37 (.A(wb_dat_i[0]),
    .Z(net37));
 BUF_X1 input38 (.A(wb_dat_i[10]),
    .Z(net38));
 BUF_X1 input39 (.A(wb_dat_i[11]),
    .Z(net39));
 BUF_X1 input40 (.A(wb_dat_i[12]),
    .Z(net40));
 BUF_X1 input41 (.A(wb_dat_i[13]),
    .Z(net41));
 BUF_X1 input42 (.A(wb_dat_i[14]),
    .Z(net42));
 BUF_X1 input43 (.A(wb_dat_i[15]),
    .Z(net43));
 BUF_X1 input44 (.A(wb_dat_i[16]),
    .Z(net44));
 BUF_X1 input45 (.A(wb_dat_i[17]),
    .Z(net45));
 BUF_X1 input46 (.A(wb_dat_i[18]),
    .Z(net46));
 BUF_X1 input47 (.A(wb_dat_i[19]),
    .Z(net47));
 BUF_X1 input48 (.A(wb_dat_i[1]),
    .Z(net48));
 BUF_X1 input49 (.A(wb_dat_i[20]),
    .Z(net49));
 BUF_X1 input50 (.A(wb_dat_i[21]),
    .Z(net50));
 BUF_X1 input51 (.A(wb_dat_i[22]),
    .Z(net51));
 BUF_X1 input52 (.A(wb_dat_i[23]),
    .Z(net52));
 BUF_X1 input53 (.A(wb_dat_i[24]),
    .Z(net53));
 BUF_X1 input54 (.A(wb_dat_i[25]),
    .Z(net54));
 BUF_X1 input55 (.A(wb_dat_i[26]),
    .Z(net55));
 BUF_X1 input56 (.A(wb_dat_i[27]),
    .Z(net56));
 BUF_X1 input57 (.A(wb_dat_i[28]),
    .Z(net57));
 BUF_X1 input58 (.A(wb_dat_i[29]),
    .Z(net58));
 BUF_X1 input59 (.A(wb_dat_i[2]),
    .Z(net59));
 BUF_X1 input60 (.A(wb_dat_i[30]),
    .Z(net60));
 BUF_X1 input61 (.A(wb_dat_i[31]),
    .Z(net61));
 BUF_X1 input62 (.A(wb_dat_i[3]),
    .Z(net62));
 BUF_X1 input63 (.A(wb_dat_i[4]),
    .Z(net63));
 BUF_X1 input64 (.A(wb_dat_i[5]),
    .Z(net64));
 BUF_X1 input65 (.A(wb_dat_i[6]),
    .Z(net65));
 BUF_X1 input66 (.A(wb_dat_i[7]),
    .Z(net66));
 BUF_X1 input67 (.A(wb_dat_i[8]),
    .Z(net67));
 BUF_X1 input68 (.A(wb_dat_i[9]),
    .Z(net68));
 BUF_X1 input69 (.A(wb_err_i),
    .Z(net69));
 BUF_X1 input70 (.A(wb_rty_i),
    .Z(net70));
 BUF_X1 input71 (.A(write_addr[0]),
    .Z(net71));
 BUF_X1 input72 (.A(write_addr[10]),
    .Z(net72));
 BUF_X1 input73 (.A(write_addr[11]),
    .Z(net73));
 BUF_X1 input74 (.A(write_addr[12]),
    .Z(net74));
 BUF_X1 input75 (.A(write_addr[13]),
    .Z(net75));
 BUF_X1 input76 (.A(write_addr[14]),
    .Z(net76));
 BUF_X1 input77 (.A(write_addr[15]),
    .Z(net77));
 BUF_X1 input78 (.A(write_addr[16]),
    .Z(net78));
 BUF_X1 input79 (.A(write_addr[17]),
    .Z(net79));
 BUF_X1 input80 (.A(write_addr[18]),
    .Z(net80));
 BUF_X1 input81 (.A(write_addr[19]),
    .Z(net81));
 BUF_X1 input82 (.A(write_addr[1]),
    .Z(net82));
 BUF_X1 input83 (.A(write_addr[20]),
    .Z(net83));
 BUF_X1 input84 (.A(write_addr[21]),
    .Z(net84));
 BUF_X1 input85 (.A(write_addr[22]),
    .Z(net85));
 BUF_X1 input86 (.A(write_addr[23]),
    .Z(net86));
 BUF_X1 input87 (.A(write_addr[24]),
    .Z(net87));
 BUF_X1 input88 (.A(write_addr[25]),
    .Z(net88));
 BUF_X1 input89 (.A(write_addr[26]),
    .Z(net89));
 BUF_X1 input90 (.A(write_addr[27]),
    .Z(net90));
 BUF_X1 input91 (.A(write_addr[28]),
    .Z(net91));
 BUF_X1 input92 (.A(write_addr[29]),
    .Z(net92));
 BUF_X1 input93 (.A(write_addr[2]),
    .Z(net93));
 BUF_X1 input94 (.A(write_addr[30]),
    .Z(net94));
 BUF_X1 input95 (.A(write_addr[31]),
    .Z(net95));
 BUF_X1 input96 (.A(write_addr[3]),
    .Z(net96));
 BUF_X1 input97 (.A(write_addr[4]),
    .Z(net97));
 BUF_X1 input98 (.A(write_addr[5]),
    .Z(net98));
 BUF_X1 input99 (.A(write_addr[6]),
    .Z(net99));
 BUF_X1 input100 (.A(write_addr[7]),
    .Z(net100));
 BUF_X1 input101 (.A(write_addr[8]),
    .Z(net101));
 BUF_X1 input102 (.A(write_addr[9]),
    .Z(net102));
 BUF_X1 input103 (.A(write_data[0]),
    .Z(net103));
 BUF_X1 input104 (.A(write_data[10]),
    .Z(net104));
 BUF_X1 input105 (.A(write_data[11]),
    .Z(net105));
 BUF_X1 input106 (.A(write_data[12]),
    .Z(net106));
 BUF_X1 input107 (.A(write_data[13]),
    .Z(net107));
 BUF_X1 input108 (.A(write_data[14]),
    .Z(net108));
 BUF_X1 input109 (.A(write_data[15]),
    .Z(net109));
 BUF_X1 input110 (.A(write_data[16]),
    .Z(net110));
 BUF_X1 input111 (.A(write_data[17]),
    .Z(net111));
 BUF_X1 input112 (.A(write_data[18]),
    .Z(net112));
 BUF_X1 input113 (.A(write_data[19]),
    .Z(net113));
 BUF_X1 input114 (.A(write_data[1]),
    .Z(net114));
 BUF_X1 input115 (.A(write_data[20]),
    .Z(net115));
 BUF_X1 input116 (.A(write_data[21]),
    .Z(net116));
 BUF_X1 input117 (.A(write_data[22]),
    .Z(net117));
 BUF_X1 input118 (.A(write_data[23]),
    .Z(net118));
 BUF_X1 input119 (.A(write_data[24]),
    .Z(net119));
 BUF_X1 input120 (.A(write_data[25]),
    .Z(net120));
 BUF_X1 input121 (.A(write_data[26]),
    .Z(net121));
 BUF_X1 input122 (.A(write_data[27]),
    .Z(net122));
 BUF_X1 input123 (.A(write_data[28]),
    .Z(net123));
 BUF_X1 input124 (.A(write_data[29]),
    .Z(net124));
 BUF_X1 input125 (.A(write_data[2]),
    .Z(net125));
 BUF_X1 input126 (.A(write_data[30]),
    .Z(net126));
 BUF_X1 input127 (.A(write_data[31]),
    .Z(net127));
 BUF_X1 input128 (.A(write_data[3]),
    .Z(net128));
 BUF_X1 input129 (.A(write_data[4]),
    .Z(net129));
 BUF_X1 input130 (.A(write_data[5]),
    .Z(net130));
 BUF_X1 input131 (.A(write_data[6]),
    .Z(net131));
 BUF_X1 input132 (.A(write_data[7]),
    .Z(net132));
 BUF_X1 input133 (.A(write_data[8]),
    .Z(net133));
 BUF_X1 input134 (.A(write_data[9]),
    .Z(net134));
 BUF_X1 input135 (.A(write_sel[0]),
    .Z(net135));
 BUF_X1 input136 (.A(write_sel[1]),
    .Z(net136));
 BUF_X1 input137 (.A(write_sel[2]),
    .Z(net137));
 BUF_X1 input138 (.A(write_sel[3]),
    .Z(net138));
 BUF_X1 output139 (.A(net139),
    .Z(read_data[0]));
 BUF_X1 output140 (.A(net140),
    .Z(read_data[10]));
 BUF_X1 output141 (.A(net141),
    .Z(read_data[11]));
 BUF_X1 output142 (.A(net142),
    .Z(read_data[12]));
 BUF_X1 output143 (.A(net143),
    .Z(read_data[13]));
 BUF_X1 output144 (.A(net144),
    .Z(read_data[14]));
 BUF_X1 output145 (.A(net145),
    .Z(read_data[15]));
 BUF_X1 output146 (.A(net146),
    .Z(read_data[16]));
 BUF_X1 output147 (.A(net147),
    .Z(read_data[17]));
 BUF_X1 output148 (.A(net148),
    .Z(read_data[18]));
 BUF_X1 output149 (.A(net149),
    .Z(read_data[19]));
 BUF_X1 output150 (.A(net150),
    .Z(read_data[1]));
 BUF_X1 output151 (.A(net151),
    .Z(read_data[20]));
 BUF_X1 output152 (.A(net152),
    .Z(read_data[21]));
 BUF_X1 output153 (.A(net153),
    .Z(read_data[22]));
 BUF_X1 output154 (.A(net154),
    .Z(read_data[23]));
 BUF_X1 output155 (.A(net155),
    .Z(read_data[24]));
 BUF_X1 output156 (.A(net156),
    .Z(read_data[25]));
 BUF_X1 output157 (.A(net157),
    .Z(read_data[26]));
 BUF_X1 output158 (.A(net158),
    .Z(read_data[27]));
 BUF_X1 output159 (.A(net159),
    .Z(read_data[28]));
 BUF_X1 output160 (.A(net160),
    .Z(read_data[29]));
 BUF_X1 output161 (.A(net161),
    .Z(read_data[2]));
 BUF_X1 output162 (.A(net162),
    .Z(read_data[30]));
 BUF_X1 output163 (.A(net163),
    .Z(read_data[31]));
 BUF_X1 output164 (.A(net164),
    .Z(read_data[3]));
 BUF_X1 output165 (.A(net165),
    .Z(read_data[4]));
 BUF_X1 output166 (.A(net166),
    .Z(read_data[5]));
 BUF_X1 output167 (.A(net167),
    .Z(read_data[6]));
 BUF_X1 output168 (.A(net168),
    .Z(read_data[7]));
 BUF_X1 output169 (.A(net169),
    .Z(read_data[8]));
 BUF_X1 output170 (.A(net170),
    .Z(read_data[9]));
 BUF_X1 output171 (.A(net171),
    .Z(read_done));
 BUF_X1 output172 (.A(net172),
    .Z(read_err));
 BUF_X1 output173 (.A(net173),
    .Z(wb_adr_o[0]));
 BUF_X1 output174 (.A(net174),
    .Z(wb_adr_o[10]));
 BUF_X1 output175 (.A(net175),
    .Z(wb_adr_o[11]));
 BUF_X1 output176 (.A(net176),
    .Z(wb_adr_o[12]));
 BUF_X1 output177 (.A(net177),
    .Z(wb_adr_o[13]));
 BUF_X1 output178 (.A(net178),
    .Z(wb_adr_o[14]));
 BUF_X1 output179 (.A(net179),
    .Z(wb_adr_o[15]));
 BUF_X1 output180 (.A(net180),
    .Z(wb_adr_o[16]));
 BUF_X1 output181 (.A(net181),
    .Z(wb_adr_o[17]));
 BUF_X1 output182 (.A(net182),
    .Z(wb_adr_o[18]));
 BUF_X1 output183 (.A(net183),
    .Z(wb_adr_o[19]));
 BUF_X1 output184 (.A(net184),
    .Z(wb_adr_o[1]));
 BUF_X1 output185 (.A(net185),
    .Z(wb_adr_o[20]));
 BUF_X1 output186 (.A(net186),
    .Z(wb_adr_o[21]));
 BUF_X1 output187 (.A(net187),
    .Z(wb_adr_o[22]));
 BUF_X1 output188 (.A(net188),
    .Z(wb_adr_o[23]));
 BUF_X1 output189 (.A(net189),
    .Z(wb_adr_o[24]));
 BUF_X1 output190 (.A(net190),
    .Z(wb_adr_o[25]));
 BUF_X1 output191 (.A(net191),
    .Z(wb_adr_o[26]));
 BUF_X1 output192 (.A(net192),
    .Z(wb_adr_o[27]));
 BUF_X1 output193 (.A(net193),
    .Z(wb_adr_o[28]));
 BUF_X1 output194 (.A(net194),
    .Z(wb_adr_o[29]));
 BUF_X1 output195 (.A(net195),
    .Z(wb_adr_o[2]));
 BUF_X1 output196 (.A(net196),
    .Z(wb_adr_o[30]));
 BUF_X1 output197 (.A(net197),
    .Z(wb_adr_o[31]));
 BUF_X1 output198 (.A(net198),
    .Z(wb_adr_o[3]));
 BUF_X1 output199 (.A(net199),
    .Z(wb_adr_o[4]));
 BUF_X1 output200 (.A(net200),
    .Z(wb_adr_o[5]));
 BUF_X1 output201 (.A(net201),
    .Z(wb_adr_o[6]));
 BUF_X1 output202 (.A(net202),
    .Z(wb_adr_o[7]));
 BUF_X1 output203 (.A(net203),
    .Z(wb_adr_o[8]));
 BUF_X1 output204 (.A(net204),
    .Z(wb_adr_o[9]));
 BUF_X1 output205 (.A(net205),
    .Z(wb_cyc_o));
 BUF_X1 output206 (.A(net206),
    .Z(wb_dat_o[0]));
 BUF_X1 output207 (.A(net207),
    .Z(wb_dat_o[10]));
 BUF_X1 output208 (.A(net208),
    .Z(wb_dat_o[11]));
 BUF_X1 output209 (.A(net209),
    .Z(wb_dat_o[12]));
 BUF_X1 output210 (.A(net210),
    .Z(wb_dat_o[13]));
 BUF_X1 output211 (.A(net211),
    .Z(wb_dat_o[14]));
 BUF_X1 output212 (.A(net212),
    .Z(wb_dat_o[15]));
 BUF_X1 output213 (.A(net213),
    .Z(wb_dat_o[16]));
 BUF_X1 output214 (.A(net214),
    .Z(wb_dat_o[17]));
 BUF_X1 output215 (.A(net215),
    .Z(wb_dat_o[18]));
 BUF_X1 output216 (.A(net216),
    .Z(wb_dat_o[19]));
 BUF_X1 output217 (.A(net217),
    .Z(wb_dat_o[1]));
 BUF_X1 output218 (.A(net218),
    .Z(wb_dat_o[20]));
 BUF_X1 output219 (.A(net219),
    .Z(wb_dat_o[21]));
 BUF_X1 output220 (.A(net220),
    .Z(wb_dat_o[22]));
 BUF_X1 output221 (.A(net221),
    .Z(wb_dat_o[23]));
 BUF_X1 output222 (.A(net222),
    .Z(wb_dat_o[24]));
 BUF_X1 output223 (.A(net223),
    .Z(wb_dat_o[25]));
 BUF_X1 output224 (.A(net224),
    .Z(wb_dat_o[26]));
 BUF_X1 output225 (.A(net225),
    .Z(wb_dat_o[27]));
 BUF_X1 output226 (.A(net226),
    .Z(wb_dat_o[28]));
 BUF_X1 output227 (.A(net227),
    .Z(wb_dat_o[29]));
 BUF_X1 output228 (.A(net228),
    .Z(wb_dat_o[2]));
 BUF_X1 output229 (.A(net229),
    .Z(wb_dat_o[30]));
 BUF_X1 output230 (.A(net230),
    .Z(wb_dat_o[31]));
 BUF_X1 output231 (.A(net231),
    .Z(wb_dat_o[3]));
 BUF_X1 output232 (.A(net232),
    .Z(wb_dat_o[4]));
 BUF_X1 output233 (.A(net233),
    .Z(wb_dat_o[5]));
 BUF_X1 output234 (.A(net234),
    .Z(wb_dat_o[6]));
 BUF_X1 output235 (.A(net235),
    .Z(wb_dat_o[7]));
 BUF_X1 output236 (.A(net236),
    .Z(wb_dat_o[8]));
 BUF_X1 output237 (.A(net237),
    .Z(wb_dat_o[9]));
 BUF_X1 output238 (.A(net238),
    .Z(wb_sel_o[0]));
 BUF_X1 output239 (.A(net239),
    .Z(wb_sel_o[1]));
 BUF_X1 output240 (.A(net240),
    .Z(wb_sel_o[2]));
 BUF_X1 output241 (.A(net241),
    .Z(wb_sel_o[3]));
 BUF_X1 output242 (.A(net242),
    .Z(wb_stb_o));
 BUF_X1 output243 (.A(net243),
    .Z(wb_we_o));
 BUF_X1 output244 (.A(net244),
    .Z(write_done));
 BUF_X1 output245 (.A(net245),
    .Z(write_err));
 LOGIC0_X1 _814__246 (.Z(net246));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X1 clkload0 (.A(clknet_4_0_0_clk));
 CLKBUF_X1 clkload1 (.A(clknet_4_1_0_clk));
 INV_X1 clkload2 (.A(clknet_4_2_0_clk));
 INV_X2 clkload3 (.A(clknet_4_3_0_clk));
 INV_X2 clkload4 (.A(clknet_4_4_0_clk));
 INV_X4 clkload5 (.A(clknet_4_6_0_clk));
 INV_X2 clkload6 (.A(clknet_4_7_0_clk));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_10_0_clk));
 INV_X2 clkload10 (.A(clknet_4_11_0_clk));
 INV_X2 clkload11 (.A(clknet_4_12_0_clk));
 INV_X2 clkload12 (.A(clknet_4_13_0_clk));
 INV_X1 clkload13 (.A(clknet_4_14_0_clk));
 FILLCELL_X4 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_5 ();
 FILLCELL_X1 FILLER_0_7 ();
 FILLCELL_X4 FILLER_0_12 ();
 FILLCELL_X2 FILLER_0_16 ();
 FILLCELL_X1 FILLER_0_38 ();
 FILLCELL_X2 FILLER_0_68 ();
 FILLCELL_X1 FILLER_0_112 ();
 FILLCELL_X2 FILLER_0_116 ();
 FILLCELL_X1 FILLER_0_215 ();
 FILLCELL_X2 FILLER_0_233 ();
 FILLCELL_X1 FILLER_0_235 ();
 FILLCELL_X1 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_19 ();
 FILLCELL_X1 FILLER_1_38 ();
 FILLCELL_X1 FILLER_1_138 ();
 FILLCELL_X2 FILLER_1_197 ();
 FILLCELL_X2 FILLER_1_206 ();
 FILLCELL_X1 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_5 ();
 FILLCELL_X1 FILLER_2_30 ();
 FILLCELL_X1 FILLER_2_34 ();
 FILLCELL_X1 FILLER_2_39 ();
 FILLCELL_X1 FILLER_2_66 ();
 FILLCELL_X1 FILLER_2_91 ();
 FILLCELL_X2 FILLER_2_95 ();
 FILLCELL_X4 FILLER_2_121 ();
 FILLCELL_X2 FILLER_2_125 ();
 FILLCELL_X1 FILLER_2_127 ();
 FILLCELL_X2 FILLER_2_158 ();
 FILLCELL_X1 FILLER_2_160 ();
 FILLCELL_X1 FILLER_2_175 ();
 FILLCELL_X2 FILLER_2_203 ();
 FILLCELL_X2 FILLER_2_231 ();
 FILLCELL_X4 FILLER_3_22 ();
 FILLCELL_X2 FILLER_3_26 ();
 FILLCELL_X1 FILLER_3_28 ();
 FILLCELL_X1 FILLER_3_46 ();
 FILLCELL_X1 FILLER_3_54 ();
 FILLCELL_X8 FILLER_3_62 ();
 FILLCELL_X1 FILLER_3_70 ();
 FILLCELL_X8 FILLER_3_81 ();
 FILLCELL_X4 FILLER_3_89 ();
 FILLCELL_X2 FILLER_3_93 ();
 FILLCELL_X16 FILLER_3_106 ();
 FILLCELL_X4 FILLER_3_122 ();
 FILLCELL_X8 FILLER_3_146 ();
 FILLCELL_X4 FILLER_3_154 ();
 FILLCELL_X2 FILLER_3_158 ();
 FILLCELL_X1 FILLER_3_184 ();
 FILLCELL_X1 FILLER_3_189 ();
 FILLCELL_X1 FILLER_3_193 ();
 FILLCELL_X2 FILLER_3_227 ();
 FILLCELL_X8 FILLER_4_28 ();
 FILLCELL_X4 FILLER_4_36 ();
 FILLCELL_X1 FILLER_4_40 ();
 FILLCELL_X1 FILLER_4_45 ();
 FILLCELL_X1 FILLER_4_63 ();
 FILLCELL_X1 FILLER_4_67 ();
 FILLCELL_X2 FILLER_4_82 ();
 FILLCELL_X4 FILLER_4_91 ();
 FILLCELL_X32 FILLER_4_112 ();
 FILLCELL_X16 FILLER_4_144 ();
 FILLCELL_X2 FILLER_4_160 ();
 FILLCELL_X2 FILLER_4_169 ();
 FILLCELL_X1 FILLER_4_195 ();
 FILLCELL_X1 FILLER_4_206 ();
 FILLCELL_X1 FILLER_4_231 ();
 FILLCELL_X1 FILLER_4_235 ();
 FILLCELL_X2 FILLER_5_17 ();
 FILLCELL_X1 FILLER_5_22 ();
 FILLCELL_X16 FILLER_5_40 ();
 FILLCELL_X1 FILLER_5_56 ();
 FILLCELL_X1 FILLER_5_78 ();
 FILLCELL_X32 FILLER_5_96 ();
 FILLCELL_X2 FILLER_5_128 ();
 FILLCELL_X8 FILLER_5_137 ();
 FILLCELL_X4 FILLER_5_152 ();
 FILLCELL_X2 FILLER_5_156 ();
 FILLCELL_X1 FILLER_5_158 ();
 FILLCELL_X16 FILLER_5_176 ();
 FILLCELL_X8 FILLER_5_192 ();
 FILLCELL_X4 FILLER_5_200 ();
 FILLCELL_X2 FILLER_5_221 ();
 FILLCELL_X1 FILLER_5_223 ();
 FILLCELL_X1 FILLER_6_25 ();
 FILLCELL_X16 FILLER_6_37 ();
 FILLCELL_X8 FILLER_6_53 ();
 FILLCELL_X2 FILLER_6_61 ();
 FILLCELL_X1 FILLER_6_63 ();
 FILLCELL_X2 FILLER_6_86 ();
 FILLCELL_X2 FILLER_6_96 ();
 FILLCELL_X4 FILLER_6_102 ();
 FILLCELL_X2 FILLER_6_106 ();
 FILLCELL_X1 FILLER_6_108 ();
 FILLCELL_X4 FILLER_6_126 ();
 FILLCELL_X2 FILLER_6_130 ();
 FILLCELL_X8 FILLER_6_153 ();
 FILLCELL_X2 FILLER_6_161 ();
 FILLCELL_X1 FILLER_6_183 ();
 FILLCELL_X2 FILLER_6_201 ();
 FILLCELL_X1 FILLER_6_203 ();
 FILLCELL_X1 FILLER_6_207 ();
 FILLCELL_X1 FILLER_6_229 ();
 FILLCELL_X8 FILLER_7_25 ();
 FILLCELL_X4 FILLER_7_33 ();
 FILLCELL_X1 FILLER_7_37 ();
 FILLCELL_X4 FILLER_7_42 ();
 FILLCELL_X2 FILLER_7_46 ();
 FILLCELL_X1 FILLER_7_48 ();
 FILLCELL_X2 FILLER_7_57 ();
 FILLCELL_X4 FILLER_7_64 ();
 FILLCELL_X1 FILLER_7_68 ();
 FILLCELL_X1 FILLER_7_76 ();
 FILLCELL_X8 FILLER_7_97 ();
 FILLCELL_X2 FILLER_7_105 ();
 FILLCELL_X2 FILLER_7_111 ();
 FILLCELL_X2 FILLER_7_117 ();
 FILLCELL_X2 FILLER_7_130 ();
 FILLCELL_X4 FILLER_7_140 ();
 FILLCELL_X1 FILLER_7_144 ();
 FILLCELL_X1 FILLER_7_162 ();
 FILLCELL_X1 FILLER_7_167 ();
 FILLCELL_X4 FILLER_7_173 ();
 FILLCELL_X2 FILLER_7_177 ();
 FILLCELL_X1 FILLER_7_179 ();
 FILLCELL_X4 FILLER_7_187 ();
 FILLCELL_X2 FILLER_7_191 ();
 FILLCELL_X1 FILLER_7_197 ();
 FILLCELL_X1 FILLER_8_21 ();
 FILLCELL_X2 FILLER_8_28 ();
 FILLCELL_X1 FILLER_8_30 ();
 FILLCELL_X32 FILLER_8_42 ();
 FILLCELL_X4 FILLER_8_74 ();
 FILLCELL_X2 FILLER_8_78 ();
 FILLCELL_X1 FILLER_8_80 ();
 FILLCELL_X32 FILLER_8_85 ();
 FILLCELL_X4 FILLER_8_117 ();
 FILLCELL_X16 FILLER_8_138 ();
 FILLCELL_X8 FILLER_8_154 ();
 FILLCELL_X4 FILLER_8_162 ();
 FILLCELL_X2 FILLER_8_166 ();
 FILLCELL_X16 FILLER_8_192 ();
 FILLCELL_X8 FILLER_8_208 ();
 FILLCELL_X2 FILLER_8_216 ();
 FILLCELL_X1 FILLER_8_218 ();
 FILLCELL_X1 FILLER_8_222 ();
 FILLCELL_X1 FILLER_9_4 ();
 FILLCELL_X8 FILLER_9_29 ();
 FILLCELL_X32 FILLER_9_54 ();
 FILLCELL_X32 FILLER_9_86 ();
 FILLCELL_X32 FILLER_9_118 ();
 FILLCELL_X32 FILLER_9_150 ();
 FILLCELL_X4 FILLER_9_182 ();
 FILLCELL_X2 FILLER_9_196 ();
 FILLCELL_X1 FILLER_9_198 ();
 FILLCELL_X2 FILLER_9_209 ();
 FILLCELL_X2 FILLER_9_224 ();
 FILLCELL_X1 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_30 ();
 FILLCELL_X32 FILLER_10_62 ();
 FILLCELL_X8 FILLER_10_94 ();
 FILLCELL_X2 FILLER_10_102 ();
 FILLCELL_X1 FILLER_10_104 ();
 FILLCELL_X32 FILLER_10_109 ();
 FILLCELL_X32 FILLER_10_141 ();
 FILLCELL_X2 FILLER_10_173 ();
 FILLCELL_X1 FILLER_10_175 ();
 FILLCELL_X1 FILLER_10_232 ();
 FILLCELL_X2 FILLER_11_11 ();
 FILLCELL_X1 FILLER_11_13 ();
 FILLCELL_X8 FILLER_11_17 ();
 FILLCELL_X4 FILLER_11_39 ();
 FILLCELL_X2 FILLER_11_43 ();
 FILLCELL_X8 FILLER_11_47 ();
 FILLCELL_X2 FILLER_11_55 ();
 FILLCELL_X1 FILLER_11_57 ();
 FILLCELL_X16 FILLER_11_63 ();
 FILLCELL_X8 FILLER_11_79 ();
 FILLCELL_X1 FILLER_11_92 ();
 FILLCELL_X32 FILLER_11_98 ();
 FILLCELL_X32 FILLER_11_130 ();
 FILLCELL_X8 FILLER_11_162 ();
 FILLCELL_X1 FILLER_11_170 ();
 FILLCELL_X4 FILLER_11_175 ();
 FILLCELL_X4 FILLER_11_226 ();
 FILLCELL_X4 FILLER_12_57 ();
 FILLCELL_X2 FILLER_12_61 ();
 FILLCELL_X1 FILLER_12_63 ();
 FILLCELL_X32 FILLER_12_84 ();
 FILLCELL_X32 FILLER_12_116 ();
 FILLCELL_X16 FILLER_12_148 ();
 FILLCELL_X2 FILLER_12_198 ();
 FILLCELL_X1 FILLER_12_200 ();
 FILLCELL_X2 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_210 ();
 FILLCELL_X2 FILLER_12_221 ();
 FILLCELL_X2 FILLER_13_4 ();
 FILLCELL_X4 FILLER_13_40 ();
 FILLCELL_X1 FILLER_13_64 ();
 FILLCELL_X2 FILLER_13_74 ();
 FILLCELL_X32 FILLER_13_98 ();
 FILLCELL_X32 FILLER_13_130 ();
 FILLCELL_X16 FILLER_13_162 ();
 FILLCELL_X2 FILLER_13_178 ();
 FILLCELL_X1 FILLER_13_180 ();
 FILLCELL_X2 FILLER_13_185 ();
 FILLCELL_X1 FILLER_13_187 ();
 FILLCELL_X2 FILLER_13_195 ();
 FILLCELL_X1 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_228 ();
 FILLCELL_X2 FILLER_14_23 ();
 FILLCELL_X1 FILLER_14_25 ();
 FILLCELL_X2 FILLER_14_70 ();
 FILLCELL_X2 FILLER_14_93 ();
 FILLCELL_X2 FILLER_14_112 ();
 FILLCELL_X32 FILLER_14_118 ();
 FILLCELL_X32 FILLER_14_150 ();
 FILLCELL_X2 FILLER_14_182 ();
 FILLCELL_X8 FILLER_14_197 ();
 FILLCELL_X2 FILLER_14_205 ();
 FILLCELL_X1 FILLER_14_207 ();
 FILLCELL_X2 FILLER_14_213 ();
 FILLCELL_X1 FILLER_14_215 ();
 FILLCELL_X8 FILLER_15_25 ();
 FILLCELL_X4 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_62 ();
 FILLCELL_X16 FILLER_15_73 ();
 FILLCELL_X8 FILLER_15_89 ();
 FILLCELL_X4 FILLER_15_97 ();
 FILLCELL_X2 FILLER_15_101 ();
 FILLCELL_X32 FILLER_15_113 ();
 FILLCELL_X16 FILLER_15_145 ();
 FILLCELL_X1 FILLER_15_161 ();
 FILLCELL_X16 FILLER_15_169 ();
 FILLCELL_X8 FILLER_15_185 ();
 FILLCELL_X1 FILLER_15_193 ();
 FILLCELL_X1 FILLER_15_201 ();
 FILLCELL_X1 FILLER_15_206 ();
 FILLCELL_X1 FILLER_15_235 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X2 FILLER_16_49 ();
 FILLCELL_X1 FILLER_16_51 ();
 FILLCELL_X2 FILLER_16_64 ();
 FILLCELL_X1 FILLER_16_66 ();
 FILLCELL_X2 FILLER_16_90 ();
 FILLCELL_X1 FILLER_16_92 ();
 FILLCELL_X1 FILLER_16_97 ();
 FILLCELL_X1 FILLER_16_102 ();
 FILLCELL_X1 FILLER_16_106 ();
 FILLCELL_X2 FILLER_16_112 ();
 FILLCELL_X32 FILLER_16_128 ();
 FILLCELL_X16 FILLER_16_160 ();
 FILLCELL_X8 FILLER_16_176 ();
 FILLCELL_X2 FILLER_16_184 ();
 FILLCELL_X4 FILLER_16_190 ();
 FILLCELL_X2 FILLER_16_194 ();
 FILLCELL_X2 FILLER_16_213 ();
 FILLCELL_X1 FILLER_16_215 ();
 FILLCELL_X2 FILLER_16_221 ();
 FILLCELL_X1 FILLER_16_223 ();
 FILLCELL_X2 FILLER_16_230 ();
 FILLCELL_X1 FILLER_16_232 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X4 FILLER_17_17 ();
 FILLCELL_X32 FILLER_17_24 ();
 FILLCELL_X8 FILLER_17_56 ();
 FILLCELL_X2 FILLER_17_64 ();
 FILLCELL_X2 FILLER_17_71 ();
 FILLCELL_X1 FILLER_17_81 ();
 FILLCELL_X4 FILLER_17_84 ();
 FILLCELL_X2 FILLER_17_88 ();
 FILLCELL_X1 FILLER_17_90 ();
 FILLCELL_X2 FILLER_17_95 ();
 FILLCELL_X1 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_100 ();
 FILLCELL_X4 FILLER_17_108 ();
 FILLCELL_X2 FILLER_17_112 ();
 FILLCELL_X16 FILLER_17_116 ();
 FILLCELL_X16 FILLER_17_139 ();
 FILLCELL_X8 FILLER_17_155 ();
 FILLCELL_X1 FILLER_17_163 ();
 FILLCELL_X2 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_196 ();
 FILLCELL_X1 FILLER_17_198 ();
 FILLCELL_X8 FILLER_17_203 ();
 FILLCELL_X2 FILLER_17_211 ();
 FILLCELL_X2 FILLER_17_233 ();
 FILLCELL_X1 FILLER_17_235 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_9 ();
 FILLCELL_X2 FILLER_18_13 ();
 FILLCELL_X1 FILLER_18_15 ();
 FILLCELL_X16 FILLER_18_19 ();
 FILLCELL_X2 FILLER_18_35 ();
 FILLCELL_X2 FILLER_18_73 ();
 FILLCELL_X1 FILLER_18_75 ();
 FILLCELL_X1 FILLER_18_79 ();
 FILLCELL_X1 FILLER_18_104 ();
 FILLCELL_X2 FILLER_18_107 ();
 FILLCELL_X32 FILLER_18_126 ();
 FILLCELL_X32 FILLER_18_158 ();
 FILLCELL_X8 FILLER_18_190 ();
 FILLCELL_X1 FILLER_18_198 ();
 FILLCELL_X2 FILLER_18_234 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_3 ();
 FILLCELL_X8 FILLER_19_21 ();
 FILLCELL_X2 FILLER_19_29 ();
 FILLCELL_X1 FILLER_19_34 ();
 FILLCELL_X16 FILLER_19_38 ();
 FILLCELL_X2 FILLER_19_71 ();
 FILLCELL_X4 FILLER_19_108 ();
 FILLCELL_X1 FILLER_19_112 ();
 FILLCELL_X32 FILLER_19_149 ();
 FILLCELL_X16 FILLER_19_181 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_3 ();
 FILLCELL_X8 FILLER_20_25 ();
 FILLCELL_X4 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_37 ();
 FILLCELL_X1 FILLER_20_39 ();
 FILLCELL_X1 FILLER_20_74 ();
 FILLCELL_X1 FILLER_20_77 ();
 FILLCELL_X1 FILLER_20_86 ();
 FILLCELL_X32 FILLER_20_102 ();
 FILLCELL_X32 FILLER_20_134 ();
 FILLCELL_X8 FILLER_20_166 ();
 FILLCELL_X8 FILLER_20_178 ();
 FILLCELL_X4 FILLER_20_186 ();
 FILLCELL_X2 FILLER_20_200 ();
 FILLCELL_X1 FILLER_20_202 ();
 FILLCELL_X4 FILLER_20_217 ();
 FILLCELL_X2 FILLER_20_221 ();
 FILLCELL_X2 FILLER_20_233 ();
 FILLCELL_X1 FILLER_20_235 ();
 FILLCELL_X32 FILLER_21_18 ();
 FILLCELL_X4 FILLER_21_50 ();
 FILLCELL_X1 FILLER_21_54 ();
 FILLCELL_X8 FILLER_21_62 ();
 FILLCELL_X1 FILLER_21_70 ();
 FILLCELL_X1 FILLER_21_75 ();
 FILLCELL_X2 FILLER_21_87 ();
 FILLCELL_X32 FILLER_21_100 ();
 FILLCELL_X16 FILLER_21_132 ();
 FILLCELL_X4 FILLER_21_148 ();
 FILLCELL_X1 FILLER_21_152 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_208 ();
 FILLCELL_X2 FILLER_21_217 ();
 FILLCELL_X1 FILLER_22_7 ();
 FILLCELL_X8 FILLER_22_32 ();
 FILLCELL_X2 FILLER_22_40 ();
 FILLCELL_X1 FILLER_22_42 ();
 FILLCELL_X8 FILLER_22_67 ();
 FILLCELL_X2 FILLER_22_75 ();
 FILLCELL_X2 FILLER_22_83 ();
 FILLCELL_X2 FILLER_22_87 ();
 FILLCELL_X1 FILLER_22_89 ();
 FILLCELL_X1 FILLER_22_93 ();
 FILLCELL_X2 FILLER_22_98 ();
 FILLCELL_X1 FILLER_22_100 ();
 FILLCELL_X8 FILLER_22_118 ();
 FILLCELL_X4 FILLER_22_126 ();
 FILLCELL_X2 FILLER_22_130 ();
 FILLCELL_X1 FILLER_22_132 ();
 FILLCELL_X32 FILLER_22_137 ();
 FILLCELL_X16 FILLER_22_169 ();
 FILLCELL_X4 FILLER_22_185 ();
 FILLCELL_X1 FILLER_22_189 ();
 FILLCELL_X1 FILLER_22_201 ();
 FILLCELL_X1 FILLER_22_209 ();
 FILLCELL_X1 FILLER_22_227 ();
 FILLCELL_X2 FILLER_22_231 ();
 FILLCELL_X8 FILLER_23_35 ();
 FILLCELL_X16 FILLER_23_51 ();
 FILLCELL_X1 FILLER_23_67 ();
 FILLCELL_X4 FILLER_23_89 ();
 FILLCELL_X32 FILLER_23_101 ();
 FILLCELL_X8 FILLER_23_133 ();
 FILLCELL_X4 FILLER_23_141 ();
 FILLCELL_X2 FILLER_23_145 ();
 FILLCELL_X1 FILLER_23_147 ();
 FILLCELL_X1 FILLER_23_165 ();
 FILLCELL_X2 FILLER_23_187 ();
 FILLCELL_X1 FILLER_23_206 ();
 FILLCELL_X1 FILLER_23_224 ();
 FILLCELL_X2 FILLER_23_231 ();
 FILLCELL_X32 FILLER_24_18 ();
 FILLCELL_X8 FILLER_24_50 ();
 FILLCELL_X2 FILLER_24_58 ();
 FILLCELL_X1 FILLER_24_60 ();
 FILLCELL_X8 FILLER_24_64 ();
 FILLCELL_X4 FILLER_24_72 ();
 FILLCELL_X2 FILLER_24_76 ();
 FILLCELL_X8 FILLER_24_83 ();
 FILLCELL_X4 FILLER_24_91 ();
 FILLCELL_X16 FILLER_24_112 ();
 FILLCELL_X8 FILLER_24_128 ();
 FILLCELL_X1 FILLER_24_140 ();
 FILLCELL_X8 FILLER_24_143 ();
 FILLCELL_X2 FILLER_24_159 ();
 FILLCELL_X8 FILLER_24_168 ();
 FILLCELL_X2 FILLER_24_176 ();
 FILLCELL_X1 FILLER_24_178 ();
 FILLCELL_X4 FILLER_24_186 ();
 FILLCELL_X1 FILLER_24_190 ();
 FILLCELL_X2 FILLER_24_202 ();
 FILLCELL_X2 FILLER_24_217 ();
 FILLCELL_X2 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_3 ();
 FILLCELL_X8 FILLER_25_45 ();
 FILLCELL_X2 FILLER_25_53 ();
 FILLCELL_X1 FILLER_25_55 ();
 FILLCELL_X32 FILLER_25_79 ();
 FILLCELL_X2 FILLER_25_111 ();
 FILLCELL_X1 FILLER_25_113 ();
 FILLCELL_X2 FILLER_25_121 ();
 FILLCELL_X1 FILLER_25_123 ();
 FILLCELL_X4 FILLER_25_128 ();
 FILLCELL_X1 FILLER_25_158 ();
 FILLCELL_X2 FILLER_25_176 ();
 FILLCELL_X16 FILLER_25_183 ();
 FILLCELL_X2 FILLER_25_199 ();
 FILLCELL_X1 FILLER_25_201 ();
 FILLCELL_X1 FILLER_25_209 ();
 FILLCELL_X2 FILLER_25_214 ();
 FILLCELL_X4 FILLER_26_18 ();
 FILLCELL_X4 FILLER_26_26 ();
 FILLCELL_X1 FILLER_26_30 ();
 FILLCELL_X8 FILLER_26_48 ();
 FILLCELL_X16 FILLER_26_60 ();
 FILLCELL_X1 FILLER_26_76 ();
 FILLCELL_X8 FILLER_26_82 ();
 FILLCELL_X2 FILLER_26_90 ();
 FILLCELL_X2 FILLER_26_100 ();
 FILLCELL_X4 FILLER_26_136 ();
 FILLCELL_X1 FILLER_26_140 ();
 FILLCELL_X1 FILLER_26_165 ();
 FILLCELL_X8 FILLER_26_170 ();
 FILLCELL_X4 FILLER_26_178 ();
 FILLCELL_X2 FILLER_26_209 ();
 FILLCELL_X1 FILLER_26_235 ();
 FILLCELL_X8 FILLER_27_15 ();
 FILLCELL_X1 FILLER_27_23 ();
 FILLCELL_X4 FILLER_27_41 ();
 FILLCELL_X8 FILLER_27_69 ();
 FILLCELL_X2 FILLER_27_77 ();
 FILLCELL_X1 FILLER_27_79 ();
 FILLCELL_X4 FILLER_27_97 ();
 FILLCELL_X2 FILLER_27_101 ();
 FILLCELL_X4 FILLER_27_108 ();
 FILLCELL_X1 FILLER_27_112 ();
 FILLCELL_X4 FILLER_27_124 ();
 FILLCELL_X1 FILLER_27_128 ();
 FILLCELL_X8 FILLER_27_140 ();
 FILLCELL_X1 FILLER_27_148 ();
 FILLCELL_X2 FILLER_27_161 ();
 FILLCELL_X1 FILLER_27_201 ();
 FILLCELL_X1 FILLER_27_222 ();
 FILLCELL_X1 FILLER_27_226 ();
 FILLCELL_X16 FILLER_28_21 ();
 FILLCELL_X8 FILLER_28_37 ();
 FILLCELL_X1 FILLER_28_45 ();
 FILLCELL_X8 FILLER_28_63 ();
 FILLCELL_X2 FILLER_28_88 ();
 FILLCELL_X16 FILLER_28_101 ();
 FILLCELL_X8 FILLER_28_117 ();
 FILLCELL_X2 FILLER_28_125 ();
 FILLCELL_X1 FILLER_28_127 ();
 FILLCELL_X2 FILLER_28_145 ();
 FILLCELL_X4 FILLER_28_189 ();
 FILLCELL_X2 FILLER_28_193 ();
 FILLCELL_X1 FILLER_28_225 ();
 FILLCELL_X1 FILLER_28_229 ();
 FILLCELL_X1 FILLER_29_1 ();
 FILLCELL_X16 FILLER_29_5 ();
 FILLCELL_X4 FILLER_29_21 ();
 FILLCELL_X2 FILLER_29_42 ();
 FILLCELL_X1 FILLER_29_44 ();
 FILLCELL_X1 FILLER_29_70 ();
 FILLCELL_X1 FILLER_29_92 ();
 FILLCELL_X1 FILLER_29_96 ();
 FILLCELL_X8 FILLER_29_114 ();
 FILLCELL_X2 FILLER_29_122 ();
 FILLCELL_X8 FILLER_29_148 ();
 FILLCELL_X1 FILLER_29_156 ();
 FILLCELL_X1 FILLER_29_181 ();
 FILLCELL_X4 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_5 ();
 FILLCELL_X4 FILLER_30_23 ();
 FILLCELL_X1 FILLER_30_31 ();
 FILLCELL_X1 FILLER_30_42 ();
 FILLCELL_X2 FILLER_30_46 ();
 FILLCELL_X2 FILLER_30_55 ();
 FILLCELL_X1 FILLER_30_60 ();
 FILLCELL_X1 FILLER_30_116 ();
 FILLCELL_X2 FILLER_30_127 ();
 FILLCELL_X2 FILLER_30_168 ();
 FILLCELL_X2 FILLER_30_177 ();
 FILLCELL_X2 FILLER_30_217 ();
 FILLCELL_X2 FILLER_30_233 ();
 FILLCELL_X1 FILLER_30_235 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_5 ();
 FILLCELL_X8 FILLER_31_11 ();
 FILLCELL_X4 FILLER_31_19 ();
 FILLCELL_X1 FILLER_31_23 ();
 FILLCELL_X2 FILLER_31_28 ();
 FILLCELL_X1 FILLER_31_30 ();
 FILLCELL_X4 FILLER_31_47 ();
 FILLCELL_X1 FILLER_31_51 ();
 FILLCELL_X2 FILLER_31_115 ();
 FILLCELL_X1 FILLER_31_117 ();
 FILLCELL_X2 FILLER_31_124 ();
 FILLCELL_X1 FILLER_31_126 ();
 FILLCELL_X1 FILLER_31_136 ();
 FILLCELL_X1 FILLER_31_149 ();
 FILLCELL_X2 FILLER_31_190 ();
 FILLCELL_X1 FILLER_31_192 ();
 FILLCELL_X4 FILLER_31_231 ();
 FILLCELL_X1 FILLER_31_235 ();
endmodule
