module credit_based_fifo (clk,
    credit_return,
    empty,
    full,
    ready_in,
    ready_out,
    rst_n,
    valid_in,
    valid_out,
    credits_available,
    data_in,
    data_out,
    fifo_level);
 input clk;
 input credit_return;
 output empty;
 output full;
 input ready_in;
 output ready_out;
 input rst_n;
 input valid_in;
 output valid_out;
 output [4:0] credits_available;
 input [7:0] data_in;
 output [7:0] data_out;
 output [4:0] fifo_level;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \read_ptr[0] ;
 wire \read_ptr[1] ;
 wire \read_ptr[2] ;
 wire \read_ptr[3] ;
 wire \read_ptr[4] ;
 wire \write_ptr[0] ;
 wire \write_ptr[1] ;
 wire \write_ptr[2] ;
 wire \write_ptr[3] ;
 wire \write_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net36;

 sky130_fd_sc_hd__inv_1 _285_ (.A(_284_),
    .Y(net28));
 sky130_fd_sc_hd__xor2_2 _286_ (.A(\write_ptr[4] ),
    .B(\read_ptr[4] ),
    .X(_038_));
 sky130_fd_sc_hd__a21o_1 _287_ (.A1(_250_),
    .A2(_245_),
    .B1(_249_),
    .X(_039_));
 sky130_fd_sc_hd__a21oi_1 _288_ (.A1(_261_),
    .A2(_039_),
    .B1(_260_),
    .Y(_040_));
 sky130_fd_sc_hd__xnor2_2 _289_ (.A(_038_),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__clkinvlp_4 _290_ (.A(_041_),
    .Y(net32));
 sky130_fd_sc_hd__nand3b_1 _291_ (.A_N(_283_),
    .B(_251_),
    .C(_250_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_1 _292_ (.A1(_250_),
    .A2(_258_),
    .B1(_249_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_1 _293_ (.A(_250_),
    .B(_245_),
    .Y(_044_));
 sky130_fd_sc_hd__or2b_1 _294_ (.A(_284_),
    .B_N(net29),
    .X(_045_));
 sky130_fd_sc_hd__a2111oi_1 _295_ (.A1(_042_),
    .A2(_043_),
    .B1(_044_),
    .C1(_045_),
    .D1(_261_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_1 _296_ (.A(_044_),
    .Y(net30));
 sky130_fd_sc_hd__and3b_1 _297_ (.A_N(_284_),
    .B(net29),
    .C(_261_),
    .X(_047_));
 sky130_fd_sc_hd__and4_1 _298_ (.A(_042_),
    .B(_043_),
    .C(net30),
    .D(_047_),
    .X(_048_));
 sky130_fd_sc_hd__nor2_1 _299_ (.A(_046_),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__nand2_1 _300_ (.A(_041_),
    .B(_049_),
    .Y(net33));
 sky130_fd_sc_hd__or4_1 _301_ (.A(net17),
    .B(net18),
    .C(net16),
    .D(net15),
    .X(_050_));
 sky130_fd_sc_hd__nor2_2 _302_ (.A(net14),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2b_1 _303_ (.A(_051_),
    .B_N(net13),
    .Y(_052_));
 sky130_fd_sc_hd__and3_1 _304_ (.A(_041_),
    .B(_049_),
    .C(_052_),
    .X(_053_));
 sky130_fd_sc_hd__buf_6 _305_ (.A(_053_),
    .X(_253_));
 sky130_fd_sc_hd__inv_1 _306_ (.A(_253_),
    .Y(_255_));
 sky130_fd_sc_hd__nand4_1 _307_ (.A(_261_),
    .B(_250_),
    .C(_251_),
    .D(_284_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _308_ (.A(_038_),
    .B(_054_),
    .Y(net27));
 sky130_fd_sc_hd__inv_1 _309_ (.A(net11),
    .Y(_055_));
 sky130_fd_sc_hd__a21oi_4 _310_ (.A1(net35),
    .A2(_055_),
    .B1(net27),
    .Y(_056_));
 sky130_fd_sc_hd__and2_4 _311_ (.A(net12),
    .B(_056_),
    .X(_016_));
 sky130_fd_sc_hd__or2_2 _312_ (.A(_046_),
    .B(_048_),
    .X(_057_));
 sky130_fd_sc_hd__nor3_4 _313_ (.A(net32),
    .B(_057_),
    .C(_051_),
    .Y(_058_));
 sky130_fd_sc_hd__buf_6 _314_ (.A(_058_),
    .X(net34));
 sky130_fd_sc_hd__nand2_1 _315_ (.A(net13),
    .B(net12),
    .Y(_059_));
 sky130_fd_sc_hd__nor3_1 _316_ (.A(\write_ptr[3] ),
    .B(\write_ptr[2] ),
    .C(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__and3_4 _317_ (.A(_270_),
    .B(net34),
    .C(_060_),
    .X(_015_));
 sky130_fd_sc_hd__and3_4 _318_ (.A(_273_),
    .B(net34),
    .C(_060_),
    .X(_014_));
 sky130_fd_sc_hd__and3_4 _319_ (.A(_271_),
    .B(net34),
    .C(_060_),
    .X(_013_));
 sky130_fd_sc_hd__and3_4 _320_ (.A(_275_),
    .B(net34),
    .C(_060_),
    .X(_012_));
 sky130_fd_sc_hd__inv_1 _321_ (.A(\write_ptr[2] ),
    .Y(_061_));
 sky130_fd_sc_hd__nor3_1 _322_ (.A(\write_ptr[3] ),
    .B(_061_),
    .C(_059_),
    .Y(_062_));
 sky130_fd_sc_hd__and3_4 _323_ (.A(_270_),
    .B(net34),
    .C(_062_),
    .X(_011_));
 sky130_fd_sc_hd__and3_4 _324_ (.A(_273_),
    .B(net34),
    .C(_062_),
    .X(_010_));
 sky130_fd_sc_hd__and3_4 _325_ (.A(_271_),
    .B(net34),
    .C(_062_),
    .X(_009_));
 sky130_fd_sc_hd__and3_4 _326_ (.A(_275_),
    .B(net34),
    .C(_062_),
    .X(_008_));
 sky130_fd_sc_hd__nand3_1 _327_ (.A(net13),
    .B(net12),
    .C(\write_ptr[3] ),
    .Y(_063_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(\write_ptr[2] ),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__and3_4 _329_ (.A(_270_),
    .B(net34),
    .C(_064_),
    .X(_007_));
 sky130_fd_sc_hd__and3_4 _330_ (.A(_273_),
    .B(_058_),
    .C(_064_),
    .X(_006_));
 sky130_fd_sc_hd__and3_4 _331_ (.A(_271_),
    .B(_058_),
    .C(_064_),
    .X(_005_));
 sky130_fd_sc_hd__and3_4 _332_ (.A(_275_),
    .B(_058_),
    .C(_064_),
    .X(_004_));
 sky130_fd_sc_hd__nor2_1 _333_ (.A(_061_),
    .B(_063_),
    .Y(_065_));
 sky130_fd_sc_hd__and3_4 _334_ (.A(_270_),
    .B(_058_),
    .C(_065_),
    .X(_003_));
 sky130_fd_sc_hd__and3_4 _335_ (.A(_273_),
    .B(_058_),
    .C(_065_),
    .X(_002_));
 sky130_fd_sc_hd__and3_4 _336_ (.A(_275_),
    .B(_058_),
    .C(_065_),
    .X(_000_));
 sky130_fd_sc_hd__and3_4 _337_ (.A(_271_),
    .B(_058_),
    .C(_065_),
    .X(_001_));
 sky130_fd_sc_hd__buf_4 _338_ (.A(_267_),
    .X(_066_));
 sky130_fd_sc_hd__clkbuf_4 _339_ (.A(_265_),
    .X(_067_));
 sky130_fd_sc_hd__a22oi_1 _340_ (.A1(_066_),
    .A2(\mem[15][0] ),
    .B1(\mem[13][0] ),
    .B2(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__buf_4 _341_ (.A(_262_),
    .X(_069_));
 sky130_fd_sc_hd__nand2_1 _342_ (.A(\mem[8][0] ),
    .B(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__clkbuf_4 _343_ (.A(_267_),
    .X(_071_));
 sky130_fd_sc_hd__a222oi_1 _344_ (.A1(_071_),
    .A2(\mem[7][0] ),
    .B1(\mem[4][0] ),
    .B2(_262_),
    .C1(_067_),
    .C2(\mem[5][0] ),
    .Y(_072_));
 sky130_fd_sc_hd__clkbuf_4 _345_ (.A(_263_),
    .X(_073_));
 sky130_fd_sc_hd__buf_4 _346_ (.A(_073_),
    .X(_074_));
 sky130_fd_sc_hd__a22oi_1 _347_ (.A1(_066_),
    .A2(\mem[3][0] ),
    .B1(\mem[2][0] ),
    .B2(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__inv_1 _348_ (.A(\read_ptr[2] ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_1 _349_ (.A(\read_ptr[3] ),
    .Y(_077_));
 sky130_fd_sc_hd__buf_4 _350_ (.A(_077_),
    .X(_259_));
 sky130_fd_sc_hd__mux4_1 _351_ (.A0(_068_),
    .A1(_070_),
    .A2(_072_),
    .A3(_075_),
    .S0(_076_),
    .S1(_259_),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_4 _352_ (.A(\read_ptr[3] ),
    .X(_079_));
 sky130_fd_sc_hd__buf_4 _353_ (.A(\read_ptr[2] ),
    .X(_080_));
 sky130_fd_sc_hd__o21ai_1 _354_ (.A1(_079_),
    .A2(_080_),
    .B1(_069_),
    .Y(_081_));
 sky130_fd_sc_hd__nor3_1 _355_ (.A(_066_),
    .B(_073_),
    .C(_067_),
    .Y(_082_));
 sky130_fd_sc_hd__nand2_2 _356_ (.A(_081_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__buf_4 _357_ (.A(_083_),
    .X(_084_));
 sky130_fd_sc_hd__clkbuf_4 _358_ (.A(_080_),
    .X(_085_));
 sky130_fd_sc_hd__buf_4 _359_ (.A(_085_),
    .X(_086_));
 sky130_fd_sc_hd__buf_4 _360_ (.A(_262_),
    .X(_087_));
 sky130_fd_sc_hd__clkbuf_4 _361_ (.A(_073_),
    .X(_088_));
 sky130_fd_sc_hd__a22oi_1 _362_ (.A1(\mem[12][0] ),
    .A2(_087_),
    .B1(_088_),
    .B2(\mem[14][0] ),
    .Y(_089_));
 sky130_fd_sc_hd__nand3_1 _363_ (.A(_259_),
    .B(\mem[6][0] ),
    .C(_088_),
    .Y(_090_));
 sky130_fd_sc_hd__o21ai_0 _364_ (.A1(_259_),
    .A2(_089_),
    .B1(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__buf_4 _365_ (.A(_076_),
    .X(_248_));
 sky130_fd_sc_hd__buf_4 _366_ (.A(_067_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(\mem[1][0] ),
    .A1(\mem[9][0] ),
    .S(\read_ptr[3] ),
    .X(_093_));
 sky130_fd_sc_hd__a22o_1 _368_ (.A1(_066_),
    .A2(\mem[11][0] ),
    .B1(\mem[10][0] ),
    .B2(_074_),
    .X(_094_));
 sky130_fd_sc_hd__nor2b_1 _369_ (.A(_080_),
    .B_N(\read_ptr[3] ),
    .Y(_095_));
 sky130_fd_sc_hd__a32o_1 _370_ (.A1(_248_),
    .A2(_092_),
    .A3(_093_),
    .B1(_094_),
    .B2(_095_),
    .X(_096_));
 sky130_fd_sc_hd__a21oi_1 _371_ (.A1(_086_),
    .A2(_091_),
    .B1(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _372_ (.A(\mem[0][0] ),
    .B(_084_),
    .Y(_098_));
 sky130_fd_sc_hd__a31oi_1 _373_ (.A1(_078_),
    .A2(_084_),
    .A3(_097_),
    .B1(_098_),
    .Y(_235_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(\mem[2][1] ),
    .A1(\mem[6][1] ),
    .S(\read_ptr[2] ),
    .X(_099_));
 sky130_fd_sc_hd__a21oi_1 _375_ (.A1(_074_),
    .A2(_099_),
    .B1(_079_),
    .Y(_100_));
 sky130_fd_sc_hd__buf_4 _376_ (.A(_265_),
    .X(_101_));
 sky130_fd_sc_hd__a22oi_1 _377_ (.A1(\mem[4][1] ),
    .A2(_069_),
    .B1(_101_),
    .B2(\mem[5][1] ),
    .Y(_102_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\mem[10][1] ),
    .A1(\mem[14][1] ),
    .S(\read_ptr[2] ),
    .X(_103_));
 sky130_fd_sc_hd__nor2b_1 _379_ (.A(_080_),
    .B_N(_071_),
    .Y(_104_));
 sky130_fd_sc_hd__a221oi_2 _380_ (.A1(_074_),
    .A2(_103_),
    .B1(_104_),
    .B2(\mem[11][1] ),
    .C1(_077_),
    .Y(_105_));
 sky130_fd_sc_hd__a22oi_1 _381_ (.A1(_066_),
    .A2(\mem[15][1] ),
    .B1(\mem[13][1] ),
    .B2(_101_),
    .Y(_106_));
 sky130_fd_sc_hd__a22oi_1 _382_ (.A1(_100_),
    .A2(_102_),
    .B1(_105_),
    .B2(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o21ai_0 _383_ (.A1(_100_),
    .A2(_105_),
    .B1(_248_),
    .Y(_108_));
 sky130_fd_sc_hd__buf_4 _384_ (.A(_079_),
    .X(_109_));
 sky130_fd_sc_hd__nor2b_1 _385_ (.A(\read_ptr[3] ),
    .B_N(_071_),
    .Y(_110_));
 sky130_fd_sc_hd__a32oi_1 _386_ (.A1(_109_),
    .A2(\mem[12][1] ),
    .A3(_087_),
    .B1(_110_),
    .B2(\mem[7][1] ),
    .Y(_111_));
 sky130_fd_sc_hd__nand2_1 _387_ (.A(_086_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__a32oi_1 _388_ (.A1(_079_),
    .A2(\mem[8][1] ),
    .A3(_087_),
    .B1(_110_),
    .B2(\mem[3][1] ),
    .Y(_113_));
 sky130_fd_sc_hd__mux2_1 _389_ (.A0(\mem[1][1] ),
    .A1(\mem[9][1] ),
    .S(\read_ptr[3] ),
    .X(_114_));
 sky130_fd_sc_hd__nand2_1 _390_ (.A(_092_),
    .B(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__nand3_1 _391_ (.A(_248_),
    .B(_113_),
    .C(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__a22oi_1 _392_ (.A1(_107_),
    .A2(_108_),
    .B1(_112_),
    .B2(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _393_ (.A(\mem[0][1] ),
    .B(_084_),
    .Y(_118_));
 sky130_fd_sc_hd__a21oi_1 _394_ (.A1(_084_),
    .A2(_117_),
    .B1(_118_),
    .Y(_236_));
 sky130_fd_sc_hd__mux2i_1 _395_ (.A0(\mem[2][2] ),
    .A1(\mem[6][2] ),
    .S(_080_),
    .Y(_119_));
 sky130_fd_sc_hd__nand2_1 _396_ (.A(\mem[10][2] ),
    .B(_095_),
    .Y(_120_));
 sky130_fd_sc_hd__o21ai_0 _397_ (.A1(_079_),
    .A2(_119_),
    .B1(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__a22oi_1 _398_ (.A1(_066_),
    .A2(\mem[15][2] ),
    .B1(\mem[14][2] ),
    .B2(_074_),
    .Y(_122_));
 sky130_fd_sc_hd__a221oi_1 _399_ (.A1(\mem[4][2] ),
    .A2(_069_),
    .B1(_101_),
    .B2(\mem[5][2] ),
    .C1(_079_),
    .Y(_123_));
 sky130_fd_sc_hd__a21oi_1 _400_ (.A1(_109_),
    .A2(_122_),
    .B1(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__clkbuf_4 _401_ (.A(_080_),
    .X(_125_));
 sky130_fd_sc_hd__a32oi_1 _402_ (.A1(_079_),
    .A2(\mem[8][2] ),
    .A3(_087_),
    .B1(_110_),
    .B2(\mem[3][2] ),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _403_ (.A(_125_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__a221oi_1 _404_ (.A1(_088_),
    .A2(_121_),
    .B1(_124_),
    .B2(_086_),
    .C1(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__buf_4 _405_ (.A(_079_),
    .X(_129_));
 sky130_fd_sc_hd__nand2_1 _406_ (.A(\mem[1][2] ),
    .B(_092_),
    .Y(_130_));
 sky130_fd_sc_hd__clkbuf_4 _407_ (.A(_066_),
    .X(_131_));
 sky130_fd_sc_hd__nand3_1 _408_ (.A(_125_),
    .B(_131_),
    .C(\mem[7][2] ),
    .Y(_132_));
 sky130_fd_sc_hd__o21ai_0 _409_ (.A1(_125_),
    .A2(_130_),
    .B1(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__a221oi_1 _410_ (.A1(_066_),
    .A2(\mem[11][2] ),
    .B1(\mem[9][2] ),
    .B2(_101_),
    .C1(_085_),
    .Y(_134_));
 sky130_fd_sc_hd__a221oi_1 _411_ (.A1(\mem[12][2] ),
    .A2(_069_),
    .B1(_092_),
    .B2(\mem[13][2] ),
    .C1(_248_),
    .Y(_135_));
 sky130_fd_sc_hd__o21ai_0 _412_ (.A1(_134_),
    .A2(_135_),
    .B1(_109_),
    .Y(_136_));
 sky130_fd_sc_hd__o21ai_0 _413_ (.A1(_129_),
    .A2(_133_),
    .B1(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__nor2_1 _414_ (.A(\mem[0][2] ),
    .B(_084_),
    .Y(_138_));
 sky130_fd_sc_hd__a31oi_1 _415_ (.A1(_084_),
    .A2(_128_),
    .A3(_137_),
    .B1(_138_),
    .Y(_237_));
 sky130_fd_sc_hd__a222oi_1 _416_ (.A1(_071_),
    .A2(\mem[15][3] ),
    .B1(\mem[12][3] ),
    .B2(_262_),
    .C1(_067_),
    .C2(\mem[13][3] ),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _417_ (.A(\mem[10][3] ),
    .B(_074_),
    .Y(_140_));
 sky130_fd_sc_hd__a222oi_1 _418_ (.A1(_071_),
    .A2(\mem[7][3] ),
    .B1(\mem[6][3] ),
    .B2(_073_),
    .C1(_265_),
    .C2(\mem[5][3] ),
    .Y(_141_));
 sky130_fd_sc_hd__a222oi_1 _419_ (.A1(_071_),
    .A2(\mem[3][3] ),
    .B1(\mem[2][3] ),
    .B2(_073_),
    .C1(_067_),
    .C2(\mem[1][3] ),
    .Y(_142_));
 sky130_fd_sc_hd__mux4_1 _420_ (.A0(_139_),
    .A1(_140_),
    .A2(_141_),
    .A3(_142_),
    .S0(_076_),
    .S1(_259_),
    .X(_143_));
 sky130_fd_sc_hd__a22oi_1 _421_ (.A1(_066_),
    .A2(\mem[11][3] ),
    .B1(\mem[9][3] ),
    .B2(_101_),
    .Y(_144_));
 sky130_fd_sc_hd__nand3_1 _422_ (.A(_085_),
    .B(\mem[14][3] ),
    .C(_088_),
    .Y(_145_));
 sky130_fd_sc_hd__o21ai_0 _423_ (.A1(_085_),
    .A2(_144_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nand2_1 _424_ (.A(_085_),
    .B(\mem[4][3] ),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(\mem[8][3] ),
    .B(_095_),
    .Y(_148_));
 sky130_fd_sc_hd__o21ai_0 _426_ (.A1(_109_),
    .A2(_147_),
    .B1(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__a22oi_1 _427_ (.A1(_129_),
    .A2(_146_),
    .B1(_149_),
    .B2(_087_),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_1 _428_ (.A(\mem[0][3] ),
    .B(_084_),
    .Y(_151_));
 sky130_fd_sc_hd__a31oi_1 _429_ (.A1(_084_),
    .A2(_143_),
    .A3(_150_),
    .B1(_151_),
    .Y(_238_));
 sky130_fd_sc_hd__nand3_1 _430_ (.A(\mem[0][4] ),
    .B(_081_),
    .C(_082_),
    .Y(_152_));
 sky130_fd_sc_hd__a22oi_1 _431_ (.A1(_131_),
    .A2(\mem[7][4] ),
    .B1(\mem[6][4] ),
    .B2(_088_),
    .Y(_153_));
 sky130_fd_sc_hd__a221oi_1 _432_ (.A1(_131_),
    .A2(\mem[3][4] ),
    .B1(\mem[2][4] ),
    .B2(_088_),
    .C1(_085_),
    .Y(_154_));
 sky130_fd_sc_hd__a21oi_1 _433_ (.A1(_086_),
    .A2(_153_),
    .B1(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a221oi_1 _434_ (.A1(_131_),
    .A2(\mem[11][4] ),
    .B1(\mem[10][4] ),
    .B2(_088_),
    .C1(_125_),
    .Y(_156_));
 sky130_fd_sc_hd__a221oi_1 _435_ (.A1(_131_),
    .A2(\mem[15][4] ),
    .B1(\mem[13][4] ),
    .B2(_092_),
    .C1(_248_),
    .Y(_157_));
 sky130_fd_sc_hd__o21ai_0 _436_ (.A1(_156_),
    .A2(_157_),
    .B1(_129_),
    .Y(_158_));
 sky130_fd_sc_hd__o21ai_0 _437_ (.A1(_129_),
    .A2(_155_),
    .B1(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__a22oi_1 _438_ (.A1(\mem[8][4] ),
    .A2(_087_),
    .B1(_092_),
    .B2(\mem[9][4] ),
    .Y(_160_));
 sky130_fd_sc_hd__nand3_1 _439_ (.A(_259_),
    .B(\mem[1][4] ),
    .C(_092_),
    .Y(_161_));
 sky130_fd_sc_hd__o21ai_0 _440_ (.A1(_259_),
    .A2(_160_),
    .B1(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__a221oi_1 _441_ (.A1(\mem[4][4] ),
    .A2(_087_),
    .B1(_092_),
    .B2(\mem[5][4] ),
    .C1(_109_),
    .Y(_163_));
 sky130_fd_sc_hd__a221oi_1 _442_ (.A1(\mem[12][4] ),
    .A2(_087_),
    .B1(_088_),
    .B2(\mem[14][4] ),
    .C1(_259_),
    .Y(_164_));
 sky130_fd_sc_hd__o21ai_0 _443_ (.A1(_163_),
    .A2(_164_),
    .B1(_086_),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_0 _444_ (.A1(_086_),
    .A2(_162_),
    .B1(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__nand3_1 _445_ (.A(_152_),
    .B(_159_),
    .C(_166_),
    .Y(_239_));
 sky130_fd_sc_hd__a222oi_1 _446_ (.A1(_071_),
    .A2(\mem[15][5] ),
    .B1(\mem[12][5] ),
    .B2(_262_),
    .C1(_067_),
    .C2(\mem[13][5] ),
    .Y(_167_));
 sky130_fd_sc_hd__nor2_1 _447_ (.A(_248_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__a21oi_1 _448_ (.A1(\mem[11][5] ),
    .A2(_104_),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__a222oi_1 _449_ (.A1(\mem[6][5] ),
    .A2(_073_),
    .B1(_067_),
    .B2(\mem[5][5] ),
    .C1(\mem[4][5] ),
    .C2(_069_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _450_ (.A(_125_),
    .B(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__a222oi_1 _451_ (.A1(_066_),
    .A2(\mem[3][5] ),
    .B1(\mem[2][5] ),
    .B2(_073_),
    .C1(_067_),
    .C2(\mem[1][5] ),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(_248_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a21oi_1 _453_ (.A1(_171_),
    .A2(_173_),
    .B1(_109_),
    .Y(_174_));
 sky130_fd_sc_hd__a21oi_1 _454_ (.A1(_129_),
    .A2(_169_),
    .B1(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__a222oi_1 _455_ (.A1(\mem[10][5] ),
    .A2(_073_),
    .B1(_067_),
    .B2(\mem[9][5] ),
    .C1(\mem[8][5] ),
    .C2(_069_),
    .Y(_176_));
 sky130_fd_sc_hd__nand3_1 _456_ (.A(_085_),
    .B(\mem[14][5] ),
    .C(_088_),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_0 _457_ (.A1(_085_),
    .A2(_176_),
    .B1(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _458_ (.A(_129_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__nand4_1 _459_ (.A(_259_),
    .B(_086_),
    .C(_131_),
    .D(\mem[7][5] ),
    .Y(_180_));
 sky130_fd_sc_hd__nand3_1 _460_ (.A(_083_),
    .B(_179_),
    .C(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__o22a_1 _461_ (.A1(\mem[0][5] ),
    .A2(_083_),
    .B1(_175_),
    .B2(_181_),
    .X(_240_));
 sky130_fd_sc_hd__mux2i_1 _462_ (.A0(\mem[3][6] ),
    .A1(\mem[7][6] ),
    .S(_080_),
    .Y(_182_));
 sky130_fd_sc_hd__nand3_1 _463_ (.A(_109_),
    .B(_085_),
    .C(\mem[15][6] ),
    .Y(_183_));
 sky130_fd_sc_hd__o21ai_0 _464_ (.A1(_109_),
    .A2(_182_),
    .B1(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__a22oi_1 _465_ (.A1(\mem[12][6] ),
    .A2(_069_),
    .B1(_101_),
    .B2(\mem[13][6] ),
    .Y(_185_));
 sky130_fd_sc_hd__a21oi_1 _466_ (.A1(_131_),
    .A2(\mem[11][6] ),
    .B1(_085_),
    .Y(_186_));
 sky130_fd_sc_hd__a22oi_1 _467_ (.A1(\mem[10][6] ),
    .A2(_074_),
    .B1(_092_),
    .B2(\mem[9][6] ),
    .Y(_187_));
 sky130_fd_sc_hd__a22oi_1 _468_ (.A1(_125_),
    .A2(_185_),
    .B1(_186_),
    .B2(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__a22oi_1 _469_ (.A1(_131_),
    .A2(_184_),
    .B1(_188_),
    .B2(_129_),
    .Y(_189_));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(\mem[8][6] ),
    .B(_087_),
    .Y(_190_));
 sky130_fd_sc_hd__nand3_1 _471_ (.A(_125_),
    .B(\mem[14][6] ),
    .C(_088_),
    .Y(_191_));
 sky130_fd_sc_hd__o21ai_0 _472_ (.A1(_125_),
    .A2(_190_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__a222oi_1 _473_ (.A1(\mem[6][6] ),
    .A2(_073_),
    .B1(_101_),
    .B2(\mem[5][6] ),
    .C1(\mem[4][6] ),
    .C2(_069_),
    .Y(_193_));
 sky130_fd_sc_hd__a221oi_1 _474_ (.A1(\mem[2][6] ),
    .A2(_074_),
    .B1(_101_),
    .B2(\mem[1][6] ),
    .C1(_080_),
    .Y(_194_));
 sky130_fd_sc_hd__a211oi_1 _475_ (.A1(_125_),
    .A2(_193_),
    .B1(_194_),
    .C1(_109_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_1 _476_ (.A1(_129_),
    .A2(_192_),
    .B1(_195_),
    .Y(_196_));
 sky130_fd_sc_hd__nor2_1 _477_ (.A(\mem[0][6] ),
    .B(_083_),
    .Y(_197_));
 sky130_fd_sc_hd__a31oi_1 _478_ (.A1(_084_),
    .A2(_189_),
    .A3(_196_),
    .B1(_197_),
    .Y(_241_));
 sky130_fd_sc_hd__nand3_1 _479_ (.A(_079_),
    .B(\mem[8][7] ),
    .C(_087_),
    .Y(_198_));
 sky130_fd_sc_hd__nand3_1 _480_ (.A(_259_),
    .B(\mem[2][7] ),
    .C(_074_),
    .Y(_199_));
 sky130_fd_sc_hd__a21oi_1 _481_ (.A1(_198_),
    .A2(_199_),
    .B1(_125_),
    .Y(_200_));
 sky130_fd_sc_hd__a221oi_1 _482_ (.A1(\mem[6][7] ),
    .A2(_074_),
    .B1(_101_),
    .B2(\mem[5][7] ),
    .C1(_079_),
    .Y(_201_));
 sky130_fd_sc_hd__a221oi_1 _483_ (.A1(\mem[12][7] ),
    .A2(_069_),
    .B1(_101_),
    .B2(\mem[13][7] ),
    .C1(_077_),
    .Y(_202_));
 sky130_fd_sc_hd__nor3_1 _484_ (.A(_248_),
    .B(_201_),
    .C(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__a221oi_1 _485_ (.A1(_071_),
    .A2(\mem[11][7] ),
    .B1(\mem[10][7] ),
    .B2(_263_),
    .C1(_080_),
    .Y(_204_));
 sky130_fd_sc_hd__a221oi_1 _486_ (.A1(_071_),
    .A2(\mem[15][7] ),
    .B1(\mem[14][7] ),
    .B2(_073_),
    .C1(_076_),
    .Y(_205_));
 sky130_fd_sc_hd__or3_1 _487_ (.A(_077_),
    .B(_204_),
    .C(_205_),
    .X(_206_));
 sky130_fd_sc_hd__a221oi_1 _488_ (.A1(_267_),
    .A2(\mem[3][7] ),
    .B1(\mem[1][7] ),
    .B2(_265_),
    .C1(_080_),
    .Y(_207_));
 sky130_fd_sc_hd__a221oi_1 _489_ (.A1(_071_),
    .A2(\mem[7][7] ),
    .B1(\mem[4][7] ),
    .B2(_262_),
    .C1(_076_),
    .Y(_208_));
 sky130_fd_sc_hd__or3_1 _490_ (.A(\read_ptr[3] ),
    .B(_207_),
    .C(_208_),
    .X(_209_));
 sky130_fd_sc_hd__nand4_1 _491_ (.A(_109_),
    .B(_248_),
    .C(\mem[9][7] ),
    .D(_092_),
    .Y(_210_));
 sky130_fd_sc_hd__nand4_1 _492_ (.A(_083_),
    .B(_206_),
    .C(_209_),
    .D(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__o32a_1 _493_ (.A1(_200_),
    .A2(_203_),
    .A3(_211_),
    .B1(_084_),
    .B2(\mem[0][7] ),
    .X(_242_));
 sky130_fd_sc_hd__inv_1 _494_ (.A(net2),
    .Y(_252_));
 sky130_fd_sc_hd__inv_1 _495_ (.A(\read_ptr[0] ),
    .Y(_019_));
 sky130_fd_sc_hd__inv_1 _496_ (.A(\write_ptr[0] ),
    .Y(_017_));
 sky130_fd_sc_hd__inv_1 _497_ (.A(_283_),
    .Y(_244_));
 sky130_fd_sc_hd__clkinvlp_4 _498_ (.A(\read_ptr[1] ),
    .Y(_243_));
 sky130_fd_sc_hd__inv_1 _499_ (.A(\write_ptr[1] ),
    .Y(_269_));
 sky130_fd_sc_hd__a221o_2 _500_ (.A1(net18),
    .A2(_256_),
    .B1(_051_),
    .B2(_246_),
    .C1(_254_),
    .X(_212_));
 sky130_fd_sc_hd__xnor2_1 _501_ (.A(net14),
    .B(_212_),
    .Y(_022_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(_021_),
    .A1(net15),
    .S(_212_),
    .X(_023_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(_247_),
    .B(_280_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _504_ (.A(net16),
    .B(_212_),
    .Y(_214_));
 sky130_fd_sc_hd__o21ai_0 _505_ (.A1(_212_),
    .A2(_213_),
    .B1(_214_),
    .Y(_024_));
 sky130_fd_sc_hd__a21o_1 _506_ (.A1(net14),
    .A2(_278_),
    .B1(_277_),
    .X(_215_));
 sky130_fd_sc_hd__a21oi_1 _507_ (.A1(_280_),
    .A2(_215_),
    .B1(_279_),
    .Y(_216_));
 sky130_fd_sc_hd__xor2_1 _508_ (.A(_282_),
    .B(_216_),
    .X(_217_));
 sky130_fd_sc_hd__nand2_1 _509_ (.A(net17),
    .B(_212_),
    .Y(_218_));
 sky130_fd_sc_hd__o21ai_0 _510_ (.A1(_212_),
    .A2(_217_),
    .B1(_218_),
    .Y(_025_));
 sky130_fd_sc_hd__a21o_1 _511_ (.A1(_247_),
    .A2(_280_),
    .B1(_279_),
    .X(_219_));
 sky130_fd_sc_hd__a21oi_1 _512_ (.A1(_282_),
    .A2(_219_),
    .B1(_281_),
    .Y(_220_));
 sky130_fd_sc_hd__xor2_1 _513_ (.A(_246_),
    .B(_220_),
    .X(_221_));
 sky130_fd_sc_hd__nor2_1 _514_ (.A(_212_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__xor2_1 _515_ (.A(net18),
    .B(_222_),
    .X(_026_));
 sky130_fd_sc_hd__xnor2_1 _516_ (.A(_019_),
    .B(_056_),
    .Y(_027_));
 sky130_fd_sc_hd__nand2_1 _517_ (.A(_020_),
    .B(_056_),
    .Y(_223_));
 sky130_fd_sc_hd__o21ai_0 _518_ (.A1(_243_),
    .A2(_056_),
    .B1(_223_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _519_ (.A(_131_),
    .B(_056_),
    .Y(_224_));
 sky130_fd_sc_hd__xnor2_1 _520_ (.A(_086_),
    .B(_224_),
    .Y(_029_));
 sky130_fd_sc_hd__nand4_1 _521_ (.A(_086_),
    .B(\read_ptr[1] ),
    .C(\read_ptr[0] ),
    .D(_056_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_1 _522_ (.A(_129_),
    .B(_225_),
    .Y(_030_));
 sky130_fd_sc_hd__nand4_1 _523_ (.A(_129_),
    .B(_086_),
    .C(_131_),
    .D(_056_),
    .Y(_226_));
 sky130_fd_sc_hd__xnor2_1 _524_ (.A(\read_ptr[4] ),
    .B(_226_),
    .Y(_031_));
 sky130_fd_sc_hd__inv_1 _525_ (.A(net35),
    .Y(_227_));
 sky130_fd_sc_hd__o21ai_0 _526_ (.A1(_227_),
    .A2(net11),
    .B1(net27),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _527_ (.A(_017_),
    .B(_253_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(\write_ptr[1] ),
    .A1(_018_),
    .S(_253_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _529_ (.A(net13),
    .B(_275_),
    .Y(_228_));
 sky130_fd_sc_hd__nor4_1 _530_ (.A(net32),
    .B(_057_),
    .C(_051_),
    .D(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__xnor2_1 _531_ (.A(_061_),
    .B(_229_),
    .Y(_035_));
 sky130_fd_sc_hd__nand4_1 _532_ (.A(net13),
    .B(\write_ptr[2] ),
    .C(\write_ptr[1] ),
    .D(\write_ptr[0] ),
    .Y(_230_));
 sky130_fd_sc_hd__nor4_1 _533_ (.A(net32),
    .B(_057_),
    .C(_051_),
    .D(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__xor2_1 _534_ (.A(\write_ptr[3] ),
    .B(_231_),
    .X(_036_));
 sky130_fd_sc_hd__nand4_1 _535_ (.A(net13),
    .B(\write_ptr[3] ),
    .C(\write_ptr[2] ),
    .D(_275_),
    .Y(_232_));
 sky130_fd_sc_hd__nor4_1 _536_ (.A(net32),
    .B(_057_),
    .C(_051_),
    .D(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__xor2_1 _537_ (.A(\write_ptr[4] ),
    .B(_233_),
    .X(_037_));
 sky130_fd_sc_hd__nand2_1 _538_ (.A(_042_),
    .B(_043_),
    .Y(_234_));
 sky130_fd_sc_hd__xor2_1 _539_ (.A(_261_),
    .B(_234_),
    .X(net31));
 sky130_fd_sc_hd__fa_1 _540_ (.A(_243_),
    .B(\write_ptr[1] ),
    .CIN(_244_),
    .COUT(_245_),
    .SUM(net29));
 sky130_fd_sc_hd__fa_1 _541_ (.A(net14),
    .B(net15),
    .CIN(_246_),
    .COUT(_247_),
    .SUM(_021_));
 sky130_fd_sc_hd__ha_1 _542_ (.A(_248_),
    .B(\write_ptr[2] ),
    .COUT(_249_),
    .SUM(_250_));
 sky130_fd_sc_hd__ha_2 _543_ (.A(_252_),
    .B(_253_),
    .COUT(_246_),
    .SUM(_254_));
 sky130_fd_sc_hd__ha_1 _544_ (.A(net2),
    .B(_255_),
    .COUT(_256_),
    .SUM(_257_));
 sky130_fd_sc_hd__ha_1 _545_ (.A(_243_),
    .B(\write_ptr[1] ),
    .COUT(_258_),
    .SUM(_251_));
 sky130_fd_sc_hd__ha_1 _546_ (.A(_259_),
    .B(\write_ptr[3] ),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__ha_2 _547_ (.A(_019_),
    .B(_243_),
    .COUT(_262_),
    .SUM(_020_));
 sky130_fd_sc_hd__ha_1 _548_ (.A(_019_),
    .B(\read_ptr[1] ),
    .COUT(_263_),
    .SUM(_264_));
 sky130_fd_sc_hd__ha_1 _549_ (.A(\read_ptr[0] ),
    .B(_243_),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_1 _550_ (.A(\read_ptr[0] ),
    .B(\read_ptr[1] ),
    .COUT(_267_),
    .SUM(_268_));
 sky130_fd_sc_hd__ha_1 _551_ (.A(_017_),
    .B(_269_),
    .COUT(_270_),
    .SUM(_018_));
 sky130_fd_sc_hd__ha_1 _552_ (.A(_017_),
    .B(\write_ptr[1] ),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _553_ (.A(\write_ptr[0] ),
    .B(_269_),
    .COUT(_273_),
    .SUM(_274_));
 sky130_fd_sc_hd__ha_1 _554_ (.A(\write_ptr[0] ),
    .B(\write_ptr[1] ),
    .COUT(_275_),
    .SUM(_276_));
 sky130_fd_sc_hd__ha_1 _555_ (.A(net15),
    .B(_246_),
    .COUT(_277_),
    .SUM(_278_));
 sky130_fd_sc_hd__ha_1 _556_ (.A(net16),
    .B(_246_),
    .COUT(_279_),
    .SUM(_280_));
 sky130_fd_sc_hd__ha_1 _557_ (.A(net17),
    .B(_246_),
    .COUT(_281_),
    .SUM(_282_));
 sky130_fd_sc_hd__ha_1 _558_ (.A(\read_ptr[0] ),
    .B(_017_),
    .COUT(_283_),
    .SUM(_284_));
 sky130_fd_sc_hd__dfrtp_2 \credit_count[0]$_DFFE_PN0P_  (.D(_022_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \credit_count[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \credit_count[2]$_DFFE_PN0P_  (.D(_024_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \credit_count[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfstp_1 \credit_count[4]$_DFFE_PN1P_  (.D(_026_),
    .Q(net18),
    .SET_B(net12),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[0]$_DFFE_PP_  (.D(_235_),
    .DE(_016_),
    .Q(net19),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[1]$_DFFE_PP_  (.D(_236_),
    .DE(_016_),
    .Q(net20),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[2]$_DFFE_PP_  (.D(_237_),
    .DE(_016_),
    .Q(net21),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[3]$_DFFE_PP_  (.D(_238_),
    .DE(_016_),
    .Q(net22),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[4]$_DFFE_PP_  (.D(_239_),
    .DE(_016_),
    .Q(net23),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[5]$_DFFE_PP_  (.D(_240_),
    .DE(_016_),
    .Q(net24),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[6]$_DFFE_PP_  (.D(_241_),
    .DE(_016_),
    .Q(net25),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \data_out[7]$_DFFE_PP_  (.D(_242_),
    .DE(_016_),
    .Q(net26),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net3),
    .DE(_015_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net3),
    .DE(_005_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net3),
    .DE(_004_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net3),
    .DE(_003_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net3),
    .DE(_002_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net3),
    .DE(_001_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net3),
    .DE(_000_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net4),
    .DE(_000_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net5),
    .DE(_000_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net6),
    .DE(_000_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net7),
    .DE(_000_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net10),
    .DE(_000_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net3),
    .DE(_014_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net3),
    .DE(_013_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net3),
    .DE(_012_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net3),
    .DE(_011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net3),
    .DE(_010_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net3),
    .DE(_009_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net3),
    .DE(_008_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net3),
    .DE(_007_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net3),
    .DE(_006_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_ptr[0]$_DFFE_PN0P_  (.D(_027_),
    .Q(\read_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_ptr[1]$_DFFE_PN0P_  (.D(_028_),
    .Q(\read_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_ptr[2]$_DFFE_PN0P_  (.D(_029_),
    .Q(\read_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \read_ptr[3]$_DFFE_PN0P_  (.D(_030_),
    .Q(\read_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_ptr[4]$_DFFE_PN0P_  (.D(_031_),
    .Q(\read_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_out$_DFFE_PN0P_  (.D(_032_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_ptr[0]$_DFFE_PN0N_  (.D(_033_),
    .Q(\write_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \write_ptr[1]$_DFFE_PN0N_  (.D(_034_),
    .Q(\write_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \write_ptr[2]$_DFFE_PN0N_  (.D(_035_),
    .Q(\write_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \write_ptr[3]$_DFFE_PN0N_  (.D(_036_),
    .Q(\write_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_ptr[4]$_DFFE_PN0N_  (.D(_037_),
    .Q(\write_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__buf_6 hold1 (.A(net12),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_139 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(credit_return),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input2 (.A(data_in[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input3 (.A(data_in[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(data_in[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(data_in[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(data_in[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(data_in[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(data_in[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(data_in[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(ready_in),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(net36),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(valid_in),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(credits_available[0]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(credits_available[1]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(credits_available[2]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(credits_available[3]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(credits_available[4]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(fifo_level[0]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(fifo_level[1]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(fifo_level[2]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(fifo_level[3]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(fifo_level[4]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(ready_out));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(valid_out));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload13 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net36));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_231 ();
endmodule
