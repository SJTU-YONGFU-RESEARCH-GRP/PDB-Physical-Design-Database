module smart_fifo (almost_empty,
    almost_full,
    clear_errors,
    clk,
    empty,
    error_detected,
    full,
    overflow_detected,
    rd_en,
    rd_valid,
    rst_n,
    underflow_detected,
    wr_en,
    wr_ready,
    data_count,
    error_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clear_errors;
 input clk;
 output empty;
 output error_detected;
 output full;
 output overflow_detected;
 input rd_en;
 output rd_valid;
 input rst_n;
 output underflow_detected;
 input wr_en;
 output wr_ready;
 output [4:0] data_count;
 output [15:0] error_count;
 output [31:0] rd_data;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire \last_valid_data[0] ;
 wire \last_valid_data[10] ;
 wire \last_valid_data[11] ;
 wire \last_valid_data[12] ;
 wire \last_valid_data[13] ;
 wire \last_valid_data[14] ;
 wire \last_valid_data[15] ;
 wire \last_valid_data[16] ;
 wire \last_valid_data[17] ;
 wire \last_valid_data[18] ;
 wire \last_valid_data[19] ;
 wire \last_valid_data[1] ;
 wire \last_valid_data[20] ;
 wire \last_valid_data[21] ;
 wire \last_valid_data[22] ;
 wire \last_valid_data[23] ;
 wire \last_valid_data[24] ;
 wire \last_valid_data[25] ;
 wire \last_valid_data[26] ;
 wire \last_valid_data[27] ;
 wire \last_valid_data[28] ;
 wire \last_valid_data[29] ;
 wire \last_valid_data[2] ;
 wire \last_valid_data[30] ;
 wire \last_valid_data[31] ;
 wire \last_valid_data[3] ;
 wire \last_valid_data[4] ;
 wire \last_valid_data[5] ;
 wire \last_valid_data[6] ;
 wire \last_valid_data[7] ;
 wire \last_valid_data[8] ;
 wire \last_valid_data[9] ;
 wire last_valid_data_available;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;

 sky130_fd_sc_hd__inv_1 _0518_ (.A(_0517_),
    .Y(net38));
 sky130_fd_sc_hd__xor2_2 _0519_ (.A(_0505_),
    .B(_0497_),
    .X(net40));
 sky130_fd_sc_hd__nand3b_1 _0520_ (.A_N(_0516_),
    .B(_0502_),
    .C(_0505_),
    .Y(_0279_));
 sky130_fd_sc_hd__a21oi_1 _0521_ (.A1(_0505_),
    .A2(_0501_),
    .B1(_0504_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _0522_ (.A(_0279_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__xor2_1 _0523_ (.A(_0500_),
    .B(_0281_),
    .X(net41));
 sky130_fd_sc_hd__nand3_1 _0524_ (.A(_0500_),
    .B(_0505_),
    .C(_0497_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _0525_ (.A1(_0500_),
    .A2(_0504_),
    .B1(_0499_),
    .Y(_0283_));
 sky130_fd_sc_hd__xor2_2 _0526_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .X(_0284_));
 sky130_fd_sc_hd__a21oi_4 _0527_ (.A1(_0282_),
    .A2(_0283_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__and3_2 _0528_ (.A(_0282_),
    .B(_0283_),
    .C(_0284_),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_1 _0529_ (.A(_0285_),
    .B(_0286_),
    .Y(net42));
 sky130_fd_sc_hd__nand3b_1 _0530_ (.A_N(net39),
    .B(_0517_),
    .C(_0500_),
    .Y(_0287_));
 sky130_fd_sc_hd__a211o_1 _0531_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_0287_),
    .C1(net40),
    .X(_0288_));
 sky130_fd_sc_hd__nor3b_1 _0532_ (.A(_0500_),
    .B(net39),
    .C_N(_0517_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand4b_2 _0533_ (.A_N(net40),
    .B(_0279_),
    .C(_0280_),
    .D(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__a211oi_4 _0534_ (.A1(_0288_),
    .A2(_0290_),
    .B1(_0285_),
    .C1(_0286_),
    .Y(net61));
 sky130_fd_sc_hd__a2bb2oi_4 _0535_ (.A1_N(_0285_),
    .A2_N(_0286_),
    .B1(_0288_),
    .B2(_0290_),
    .Y(net43));
 sky130_fd_sc_hd__clkinv_4 _0536_ (.A(net43),
    .Y(_0291_));
 sky130_fd_sc_hd__buf_6 _0537_ (.A(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__buf_4 _0538_ (.A(_0292_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 _0539_ (.A(net133),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _0540_ (.A(_0293_),
    .B(net43),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_1 _0541_ (.A(_0294_),
    .Y(net96));
 sky130_fd_sc_hd__inv_1 _0542_ (.A(net60),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_0 _0543_ (.A1(_0295_),
    .A2(net2),
    .B1(_0294_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor2b_1 _0544_ (.A(\wr_ptr[2] ),
    .B_N(net35),
    .Y(_0296_));
 sky130_fd_sc_hd__nor2b_1 _0545_ (.A(\wr_ptr[3] ),
    .B_N(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__and2_4 _0546_ (.A(_0509_),
    .B(_0297_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_4 _0547_ (.A(_0512_),
    .B(_0297_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_4 _0548_ (.A(_0510_),
    .B(_0297_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_4 _0549_ (.A(_0514_),
    .B(_0297_),
    .X(_0010_));
 sky130_fd_sc_hd__nand2_1 _0550_ (.A(net35),
    .B(\wr_ptr[2] ),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _0551_ (.A(\wr_ptr[3] ),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__and2_4 _0552_ (.A(_0509_),
    .B(_0299_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_4 _0553_ (.A(_0512_),
    .B(_0299_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_4 _0554_ (.A(_0510_),
    .B(_0299_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_4 _0555_ (.A(_0514_),
    .B(_0299_),
    .X(_0014_));
 sky130_fd_sc_hd__and3_4 _0556_ (.A(\wr_ptr[3] ),
    .B(_0509_),
    .C(_0296_),
    .X(_0015_));
 sky130_fd_sc_hd__and3_4 _0557_ (.A(\wr_ptr[3] ),
    .B(_0512_),
    .C(_0296_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_4 _0558_ (.A(\wr_ptr[3] ),
    .B(_0510_),
    .C(_0296_),
    .X(_0002_));
 sky130_fd_sc_hd__and3_4 _0559_ (.A(\wr_ptr[3] ),
    .B(_0514_),
    .C(_0296_),
    .X(_0003_));
 sky130_fd_sc_hd__and3_1 _0560_ (.A(net35),
    .B(\wr_ptr[3] ),
    .C(\wr_ptr[2] ),
    .X(_0300_));
 sky130_fd_sc_hd__and2_4 _0561_ (.A(_0509_),
    .B(_0300_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_4 _0562_ (.A(_0512_),
    .B(_0300_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_4 _0563_ (.A(_0510_),
    .B(_0300_),
    .X(_0006_));
 sky130_fd_sc_hd__and2_4 _0564_ (.A(_0514_),
    .B(_0300_),
    .X(_0007_));
 sky130_fd_sc_hd__inv_1 _0565_ (.A(\rd_ptr[3] ),
    .Y(_0498_));
 sky130_fd_sc_hd__clkbuf_2 _0566_ (.A(\rd_ptr[1] ),
    .X(_0301_));
 sky130_fd_sc_hd__buf_4 _0567_ (.A(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__buf_6 _0568_ (.A(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__inv_1 _0569_ (.A(_0303_),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_1 _0570_ (.A(_0516_),
    .Y(_0496_));
 sky130_fd_sc_hd__buf_4 _0571_ (.A(\rd_ptr[2] ),
    .X(_0304_));
 sky130_fd_sc_hd__buf_4 _0572_ (.A(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__inv_1 _0573_ (.A(_0305_),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_1 _0574_ (.A(\wr_ptr[0] ),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_1 _0575_ (.A(\wr_ptr[1] ),
    .Y(_0508_));
 sky130_fd_sc_hd__xnor2_1 _0576_ (.A(net44),
    .B(_0294_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand4_2 _0577_ (.A(net55),
    .B(net56),
    .C(net57),
    .D(net58),
    .Y(_0306_));
 sky130_fd_sc_hd__and3_1 _0578_ (.A(net52),
    .B(net53),
    .C(net54),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _0579_ (.A(net59),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand2_2 _0580_ (.A(_0293_),
    .B(_0507_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor4_1 _0581_ (.A(_0292_),
    .B(_0306_),
    .C(_0308_),
    .D(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__xor2_1 _0582_ (.A(net45),
    .B(_0310_),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _0583_ (.A(net59),
    .B(net45),
    .Y(_0311_));
 sky130_fd_sc_hd__and3_1 _0584_ (.A(net44),
    .B(net51),
    .C(_0307_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_2 _0585_ (.A(_0293_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nor4_1 _0586_ (.A(_0291_),
    .B(_0306_),
    .C(_0311_),
    .D(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__xor2_1 _0587_ (.A(net46),
    .B(_0314_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _0588_ (.A(_0306_),
    .B(_0311_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand3_1 _0589_ (.A(net46),
    .B(_0307_),
    .C(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nor3_1 _0590_ (.A(_0292_),
    .B(_0309_),
    .C(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__xor2_1 _0591_ (.A(net47),
    .B(_0317_),
    .X(_0024_));
 sky130_fd_sc_hd__nand3_1 _0592_ (.A(net46),
    .B(net47),
    .C(_0315_),
    .Y(_0318_));
 sky130_fd_sc_hd__nor3_1 _0593_ (.A(_0292_),
    .B(_0313_),
    .C(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__xor2_1 _0594_ (.A(net48),
    .B(_0319_),
    .X(_0025_));
 sky130_fd_sc_hd__nand3_1 _0595_ (.A(net52),
    .B(net53),
    .C(net54),
    .Y(_0320_));
 sky130_fd_sc_hd__nand4_1 _0596_ (.A(net46),
    .B(net47),
    .C(net48),
    .D(_0315_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor4_1 _0597_ (.A(_0291_),
    .B(_0320_),
    .C(_0309_),
    .D(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__xor2_1 _0598_ (.A(net49),
    .B(_0322_),
    .X(_0026_));
 sky130_fd_sc_hd__nand3_1 _0599_ (.A(_0293_),
    .B(net49),
    .C(_0312_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor3_1 _0600_ (.A(_0292_),
    .B(_0321_),
    .C(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__xor2_1 _0601_ (.A(net50),
    .B(_0324_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0602_ (.A0(net51),
    .A1(_0020_),
    .S(net96),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_4 _0603_ (.A(_0291_),
    .X(_0325_));
 sky130_fd_sc_hd__nor2_1 _0604_ (.A(_0325_),
    .B(_0309_),
    .Y(_0326_));
 sky130_fd_sc_hd__xor2_1 _0605_ (.A(net52),
    .B(_0326_),
    .X(_0029_));
 sky130_fd_sc_hd__inv_1 _0606_ (.A(_0293_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand3_1 _0607_ (.A(net44),
    .B(net52),
    .C(net51),
    .Y(_0328_));
 sky130_fd_sc_hd__nor3_1 _0608_ (.A(_0327_),
    .B(_0325_),
    .C(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xor2_1 _0609_ (.A(net53),
    .B(_0329_),
    .X(_0030_));
 sky130_fd_sc_hd__nand2_1 _0610_ (.A(net52),
    .B(net53),
    .Y(_0330_));
 sky130_fd_sc_hd__nor3_1 _0611_ (.A(_0292_),
    .B(_0330_),
    .C(_0309_),
    .Y(_0331_));
 sky130_fd_sc_hd__xor2_1 _0612_ (.A(net54),
    .B(_0331_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_1 _0613_ (.A(_0325_),
    .B(_0313_),
    .Y(_0332_));
 sky130_fd_sc_hd__xor2_1 _0614_ (.A(net55),
    .B(_0332_),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_1 _0615_ (.A(net55),
    .B(_0307_),
    .Y(_0333_));
 sky130_fd_sc_hd__nor3_1 _0616_ (.A(_0292_),
    .B(_0309_),
    .C(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__xor2_1 _0617_ (.A(net56),
    .B(_0334_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _0618_ (.A(net55),
    .B(net56),
    .Y(_0335_));
 sky130_fd_sc_hd__nor3_1 _0619_ (.A(_0292_),
    .B(_0335_),
    .C(_0313_),
    .Y(_0336_));
 sky130_fd_sc_hd__xor2_1 _0620_ (.A(net57),
    .B(_0336_),
    .X(_0034_));
 sky130_fd_sc_hd__nand3_1 _0621_ (.A(net55),
    .B(net56),
    .C(net57),
    .Y(_0337_));
 sky130_fd_sc_hd__nor4_1 _0622_ (.A(_0291_),
    .B(_0320_),
    .C(_0337_),
    .D(_0309_),
    .Y(_0338_));
 sky130_fd_sc_hd__xor2_1 _0623_ (.A(net58),
    .B(_0338_),
    .X(_0035_));
 sky130_fd_sc_hd__nor3_1 _0624_ (.A(_0292_),
    .B(_0306_),
    .C(_0313_),
    .Y(_0339_));
 sky130_fd_sc_hd__xor2_1 _0625_ (.A(net59),
    .B(_0339_),
    .X(_0036_));
 sky130_fd_sc_hd__clkbuf_2 _0626_ (.A(\rd_ptr[0] ),
    .X(_0340_));
 sky130_fd_sc_hd__buf_6 _0627_ (.A(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_4 _0628_ (.A(_0304_),
    .X(_0342_));
 sky130_fd_sc_hd__mux4_1 _0629_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[4][0] ),
    .A3(\mem[5][0] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_0 _0630_ (.A(_0301_),
    .B(\rd_ptr[3] ),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_2 _0631_ (.A(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2b_2 _0632_ (.A_N(\rd_ptr[3] ),
    .B(_0301_),
    .Y(_0346_));
 sky130_fd_sc_hd__buf_4 _0633_ (.A(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__buf_6 _0634_ (.A(_0340_),
    .X(_0348_));
 sky130_fd_sc_hd__buf_6 _0635_ (.A(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_1 _0636_ (.A0(\mem[2][0] ),
    .A1(\mem[3][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_0349_),
    .S1(_0305_),
    .X(_0350_));
 sky130_fd_sc_hd__o22ai_1 _0637_ (.A1(_0343_),
    .A2(_0345_),
    .B1(_0347_),
    .B2(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__mux4_1 _0638_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S0(_0341_),
    .S1(_0302_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2b_2 _0639_ (.A_N(_0342_),
    .B(\rd_ptr[3] ),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_2 _0640_ (.A(_0342_),
    .B(\rd_ptr[3] ),
    .Y(_0354_));
 sky130_fd_sc_hd__buf_4 _0641_ (.A(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__mux4_1 _0642_ (.A0(\mem[12][0] ),
    .A1(\mem[13][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0356_));
 sky130_fd_sc_hd__o22ai_1 _0643_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0355_),
    .B2(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nor2_1 _0644_ (.A(_0351_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_8 _0645_ (.A(_0293_),
    .B(_0291_),
    .Y(_0359_));
 sky130_fd_sc_hd__buf_6 _0646_ (.A(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _0647_ (.A0(_0358_),
    .A1(\last_valid_data[0] ),
    .S(_0360_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_6 _0648_ (.A(_0348_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_8 _0649_ (.A(_0304_),
    .X(_0362_));
 sky130_fd_sc_hd__mux4_1 _0650_ (.A0(\mem[2][10] ),
    .A1(\mem[3][10] ),
    .A2(\mem[6][10] ),
    .A3(\mem[7][10] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_6 _0651_ (.A(_0348_),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_1 _0652_ (.A0(\mem[0][10] ),
    .A1(\mem[1][10] ),
    .A2(\mem[4][10] ),
    .A3(\mem[5][10] ),
    .S0(_0364_),
    .S1(_0305_),
    .X(_0365_));
 sky130_fd_sc_hd__buf_4 _0653_ (.A(_0345_),
    .X(_0366_));
 sky130_fd_sc_hd__o22ai_1 _0654_ (.A1(_0347_),
    .A2(_0363_),
    .B1(_0365_),
    .B2(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__buf_6 _0655_ (.A(_0348_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_8 _0656_ (.A(_0301_),
    .X(_0369_));
 sky130_fd_sc_hd__mux4_1 _0657_ (.A0(\mem[12][10] ),
    .A1(\mem[13][10] ),
    .A2(\mem[14][10] ),
    .A3(\mem[15][10] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__mux4_1 _0658_ (.A0(\mem[8][10] ),
    .A1(\mem[9][10] ),
    .A2(\mem[10][10] ),
    .A3(\mem[11][10] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0371_));
 sky130_fd_sc_hd__buf_4 _0659_ (.A(_0353_),
    .X(_0372_));
 sky130_fd_sc_hd__o22ai_1 _0660_ (.A1(_0355_),
    .A2(_0370_),
    .B1(_0371_),
    .B2(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__nor2_1 _0661_ (.A(_0367_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__mux2_1 _0662_ (.A0(_0374_),
    .A1(\last_valid_data[10] ),
    .S(_0360_),
    .X(_0038_));
 sky130_fd_sc_hd__mux4_1 _0663_ (.A0(\mem[2][11] ),
    .A1(\mem[3][11] ),
    .A2(\mem[6][11] ),
    .A3(\mem[7][11] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0375_));
 sky130_fd_sc_hd__mux4_1 _0664_ (.A0(\mem[0][11] ),
    .A1(\mem[1][11] ),
    .A2(\mem[4][11] ),
    .A3(\mem[5][11] ),
    .S0(_0364_),
    .S1(_0305_),
    .X(_0376_));
 sky130_fd_sc_hd__o22ai_1 _0665_ (.A1(_0347_),
    .A2(_0375_),
    .B1(_0376_),
    .B2(_0366_),
    .Y(_0377_));
 sky130_fd_sc_hd__mux4_1 _0666_ (.A0(\mem[12][11] ),
    .A1(\mem[13][11] ),
    .A2(\mem[14][11] ),
    .A3(\mem[15][11] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0378_));
 sky130_fd_sc_hd__mux4_1 _0667_ (.A0(\mem[8][11] ),
    .A1(\mem[9][11] ),
    .A2(\mem[10][11] ),
    .A3(\mem[11][11] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0379_));
 sky130_fd_sc_hd__o22ai_1 _0668_ (.A1(_0355_),
    .A2(_0378_),
    .B1(_0379_),
    .B2(_0372_),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _0669_ (.A(_0377_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__mux2_1 _0670_ (.A0(_0381_),
    .A1(\last_valid_data[11] ),
    .S(_0360_),
    .X(_0039_));
 sky130_fd_sc_hd__mux4_1 _0671_ (.A0(\mem[2][12] ),
    .A1(\mem[3][12] ),
    .A2(\mem[6][12] ),
    .A3(\mem[7][12] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0382_));
 sky130_fd_sc_hd__mux4_1 _0672_ (.A0(\mem[0][12] ),
    .A1(\mem[1][12] ),
    .A2(\mem[4][12] ),
    .A3(\mem[5][12] ),
    .S0(_0364_),
    .S1(_0305_),
    .X(_0383_));
 sky130_fd_sc_hd__o22ai_1 _0673_ (.A1(_0347_),
    .A2(_0382_),
    .B1(_0383_),
    .B2(_0366_),
    .Y(_0384_));
 sky130_fd_sc_hd__mux4_1 _0674_ (.A0(\mem[12][12] ),
    .A1(\mem[13][12] ),
    .A2(\mem[14][12] ),
    .A3(\mem[15][12] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0385_));
 sky130_fd_sc_hd__mux4_1 _0675_ (.A0(\mem[8][12] ),
    .A1(\mem[9][12] ),
    .A2(\mem[10][12] ),
    .A3(\mem[11][12] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0386_));
 sky130_fd_sc_hd__o22ai_1 _0676_ (.A1(_0355_),
    .A2(_0385_),
    .B1(_0386_),
    .B2(_0372_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _0677_ (.A(_0384_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__mux2_1 _0678_ (.A0(_0388_),
    .A1(\last_valid_data[12] ),
    .S(_0360_),
    .X(_0040_));
 sky130_fd_sc_hd__buf_6 _0679_ (.A(_0340_),
    .X(_0389_));
 sky130_fd_sc_hd__mux4_1 _0680_ (.A0(\mem[2][13] ),
    .A1(\mem[3][13] ),
    .A2(\mem[6][13] ),
    .A3(\mem[7][13] ),
    .S0(_0389_),
    .S1(_0362_),
    .X(_0390_));
 sky130_fd_sc_hd__mux4_1 _0681_ (.A0(\mem[0][13] ),
    .A1(\mem[1][13] ),
    .A2(\mem[4][13] ),
    .A3(\mem[5][13] ),
    .S0(_0364_),
    .S1(_0305_),
    .X(_0391_));
 sky130_fd_sc_hd__o22ai_1 _0682_ (.A1(_0347_),
    .A2(_0390_),
    .B1(_0391_),
    .B2(_0366_),
    .Y(_0392_));
 sky130_fd_sc_hd__mux4_1 _0683_ (.A0(\mem[12][13] ),
    .A1(\mem[13][13] ),
    .A2(\mem[14][13] ),
    .A3(\mem[15][13] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0393_));
 sky130_fd_sc_hd__mux4_1 _0684_ (.A0(\mem[8][13] ),
    .A1(\mem[9][13] ),
    .A2(\mem[10][13] ),
    .A3(\mem[11][13] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0394_));
 sky130_fd_sc_hd__o22ai_1 _0685_ (.A1(_0355_),
    .A2(_0393_),
    .B1(_0394_),
    .B2(_0372_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _0686_ (.A(_0392_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(_0396_),
    .A1(\last_valid_data[13] ),
    .S(_0360_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_4 _0688_ (.A(_0304_),
    .X(_0397_));
 sky130_fd_sc_hd__mux4_1 _0689_ (.A0(\mem[2][14] ),
    .A1(\mem[3][14] ),
    .A2(\mem[6][14] ),
    .A3(\mem[7][14] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_6 _0690_ (.A(_0348_),
    .X(_0399_));
 sky130_fd_sc_hd__mux4_1 _0691_ (.A0(\mem[0][14] ),
    .A1(\mem[1][14] ),
    .A2(\mem[4][14] ),
    .A3(\mem[5][14] ),
    .S0(_0399_),
    .S1(_0305_),
    .X(_0400_));
 sky130_fd_sc_hd__o22ai_1 _0692_ (.A1(_0347_),
    .A2(_0398_),
    .B1(_0400_),
    .B2(_0366_),
    .Y(_0401_));
 sky130_fd_sc_hd__mux4_1 _0693_ (.A0(\mem[12][14] ),
    .A1(\mem[13][14] ),
    .A2(\mem[14][14] ),
    .A3(\mem[15][14] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0402_));
 sky130_fd_sc_hd__mux4_1 _0694_ (.A0(\mem[8][14] ),
    .A1(\mem[9][14] ),
    .A2(\mem[10][14] ),
    .A3(\mem[11][14] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0403_));
 sky130_fd_sc_hd__o22ai_1 _0695_ (.A1(_0355_),
    .A2(_0402_),
    .B1(_0403_),
    .B2(_0372_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_1 _0696_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__mux2_1 _0697_ (.A0(_0405_),
    .A1(\last_valid_data[14] ),
    .S(_0360_),
    .X(_0042_));
 sky130_fd_sc_hd__mux4_1 _0698_ (.A0(\mem[2][15] ),
    .A1(\mem[3][15] ),
    .A2(\mem[6][15] ),
    .A3(\mem[7][15] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0406_));
 sky130_fd_sc_hd__buf_4 _0699_ (.A(_0304_),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _0700_ (.A0(\mem[0][15] ),
    .A1(\mem[1][15] ),
    .A2(\mem[4][15] ),
    .A3(\mem[5][15] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__o22ai_1 _0701_ (.A1(_0347_),
    .A2(_0406_),
    .B1(_0408_),
    .B2(_0366_),
    .Y(_0409_));
 sky130_fd_sc_hd__buf_6 _0702_ (.A(_0348_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_6 _0703_ (.A(_0301_),
    .X(_0411_));
 sky130_fd_sc_hd__mux4_1 _0704_ (.A0(\mem[12][15] ),
    .A1(\mem[13][15] ),
    .A2(\mem[14][15] ),
    .A3(\mem[15][15] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__mux4_1 _0705_ (.A0(\mem[8][15] ),
    .A1(\mem[9][15] ),
    .A2(\mem[10][15] ),
    .A3(\mem[11][15] ),
    .S0(_0349_),
    .S1(_0303_),
    .X(_0413_));
 sky130_fd_sc_hd__o22ai_1 _0706_ (.A1(_0355_),
    .A2(_0412_),
    .B1(_0413_),
    .B2(_0372_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor2_1 _0707_ (.A(_0409_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__mux2_1 _0708_ (.A0(_0415_),
    .A1(\last_valid_data[15] ),
    .S(_0360_),
    .X(_0043_));
 sky130_fd_sc_hd__mux4_1 _0709_ (.A0(\mem[2][16] ),
    .A1(\mem[3][16] ),
    .A2(\mem[6][16] ),
    .A3(\mem[7][16] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0416_));
 sky130_fd_sc_hd__mux4_1 _0710_ (.A0(\mem[0][16] ),
    .A1(\mem[1][16] ),
    .A2(\mem[4][16] ),
    .A3(\mem[5][16] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0417_));
 sky130_fd_sc_hd__o22ai_1 _0711_ (.A1(_0347_),
    .A2(_0416_),
    .B1(_0417_),
    .B2(_0366_),
    .Y(_0418_));
 sky130_fd_sc_hd__mux4_1 _0712_ (.A0(\mem[12][16] ),
    .A1(\mem[13][16] ),
    .A2(\mem[14][16] ),
    .A3(\mem[15][16] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_8 _0713_ (.A(_0348_),
    .X(_0420_));
 sky130_fd_sc_hd__buf_4 _0714_ (.A(_0302_),
    .X(_0421_));
 sky130_fd_sc_hd__mux4_1 _0715_ (.A0(\mem[8][16] ),
    .A1(\mem[9][16] ),
    .A2(\mem[10][16] ),
    .A3(\mem[11][16] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__o22ai_1 _0716_ (.A1(_0355_),
    .A2(_0419_),
    .B1(_0422_),
    .B2(_0372_),
    .Y(_0423_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(_0418_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__mux2_1 _0718_ (.A0(_0424_),
    .A1(\last_valid_data[16] ),
    .S(_0360_),
    .X(_0044_));
 sky130_fd_sc_hd__mux4_1 _0719_ (.A0(\mem[2][17] ),
    .A1(\mem[3][17] ),
    .A2(\mem[6][17] ),
    .A3(\mem[7][17] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0425_));
 sky130_fd_sc_hd__mux4_1 _0720_ (.A0(\mem[0][17] ),
    .A1(\mem[1][17] ),
    .A2(\mem[4][17] ),
    .A3(\mem[5][17] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0426_));
 sky130_fd_sc_hd__o22ai_1 _0721_ (.A1(_0347_),
    .A2(_0425_),
    .B1(_0426_),
    .B2(_0366_),
    .Y(_0427_));
 sky130_fd_sc_hd__mux4_1 _0722_ (.A0(\mem[12][17] ),
    .A1(\mem[13][17] ),
    .A2(\mem[14][17] ),
    .A3(\mem[15][17] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0428_));
 sky130_fd_sc_hd__mux4_1 _0723_ (.A0(\mem[8][17] ),
    .A1(\mem[9][17] ),
    .A2(\mem[10][17] ),
    .A3(\mem[11][17] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0429_));
 sky130_fd_sc_hd__o22ai_1 _0724_ (.A1(_0355_),
    .A2(_0428_),
    .B1(_0429_),
    .B2(_0372_),
    .Y(_0430_));
 sky130_fd_sc_hd__nor2_1 _0725_ (.A(_0427_),
    .B(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__buf_6 _0726_ (.A(_0359_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(_0431_),
    .A1(\last_valid_data[17] ),
    .S(_0432_),
    .X(_0045_));
 sky130_fd_sc_hd__mux4_1 _0728_ (.A0(\mem[2][18] ),
    .A1(\mem[3][18] ),
    .A2(\mem[6][18] ),
    .A3(\mem[7][18] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0433_));
 sky130_fd_sc_hd__mux4_1 _0729_ (.A0(\mem[0][18] ),
    .A1(\mem[1][18] ),
    .A2(\mem[4][18] ),
    .A3(\mem[5][18] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0434_));
 sky130_fd_sc_hd__o22ai_1 _0730_ (.A1(_0347_),
    .A2(_0433_),
    .B1(_0434_),
    .B2(_0366_),
    .Y(_0435_));
 sky130_fd_sc_hd__mux4_1 _0731_ (.A0(\mem[12][18] ),
    .A1(\mem[13][18] ),
    .A2(\mem[14][18] ),
    .A3(\mem[15][18] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0436_));
 sky130_fd_sc_hd__mux4_1 _0732_ (.A0(\mem[8][18] ),
    .A1(\mem[9][18] ),
    .A2(\mem[10][18] ),
    .A3(\mem[11][18] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0437_));
 sky130_fd_sc_hd__o22ai_1 _0733_ (.A1(_0355_),
    .A2(_0436_),
    .B1(_0437_),
    .B2(_0372_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_1 _0734_ (.A(_0435_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__mux2_1 _0735_ (.A0(_0439_),
    .A1(\last_valid_data[18] ),
    .S(_0432_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_6 _0736_ (.A(_0346_),
    .X(_0440_));
 sky130_fd_sc_hd__mux4_1 _0737_ (.A0(\mem[2][19] ),
    .A1(\mem[3][19] ),
    .A2(\mem[6][19] ),
    .A3(\mem[7][19] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0441_));
 sky130_fd_sc_hd__mux4_1 _0738_ (.A0(\mem[0][19] ),
    .A1(\mem[1][19] ),
    .A2(\mem[4][19] ),
    .A3(\mem[5][19] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0442_));
 sky130_fd_sc_hd__o22ai_1 _0739_ (.A1(_0440_),
    .A2(_0441_),
    .B1(_0442_),
    .B2(_0366_),
    .Y(_0443_));
 sky130_fd_sc_hd__buf_6 _0740_ (.A(_0354_),
    .X(_0444_));
 sky130_fd_sc_hd__mux4_1 _0741_ (.A0(\mem[12][19] ),
    .A1(\mem[13][19] ),
    .A2(\mem[14][19] ),
    .A3(\mem[15][19] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0445_));
 sky130_fd_sc_hd__mux4_1 _0742_ (.A0(\mem[8][19] ),
    .A1(\mem[9][19] ),
    .A2(\mem[10][19] ),
    .A3(\mem[11][19] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0446_));
 sky130_fd_sc_hd__o22ai_1 _0743_ (.A1(_0444_),
    .A2(_0445_),
    .B1(_0446_),
    .B2(_0372_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _0744_ (.A(_0443_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__mux2_1 _0745_ (.A0(_0448_),
    .A1(\last_valid_data[19] ),
    .S(_0432_),
    .X(_0047_));
 sky130_fd_sc_hd__mux4_1 _0746_ (.A0(\mem[2][1] ),
    .A1(\mem[3][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0449_));
 sky130_fd_sc_hd__mux4_1 _0747_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[4][1] ),
    .A3(\mem[5][1] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_4 _0748_ (.A(_0345_),
    .X(_0451_));
 sky130_fd_sc_hd__o22ai_2 _0749_ (.A1(_0440_),
    .A2(_0449_),
    .B1(_0450_),
    .B2(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__mux4_1 _0750_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0453_));
 sky130_fd_sc_hd__mux4_1 _0751_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0454_));
 sky130_fd_sc_hd__buf_6 _0752_ (.A(_0353_),
    .X(_0455_));
 sky130_fd_sc_hd__o22ai_1 _0753_ (.A1(_0444_),
    .A2(_0453_),
    .B1(_0454_),
    .B2(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nor2_1 _0754_ (.A(_0452_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(_0457_),
    .A1(\last_valid_data[1] ),
    .S(_0432_),
    .X(_0048_));
 sky130_fd_sc_hd__mux4_1 _0756_ (.A0(\mem[2][20] ),
    .A1(\mem[3][20] ),
    .A2(\mem[6][20] ),
    .A3(\mem[7][20] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0458_));
 sky130_fd_sc_hd__mux4_1 _0757_ (.A0(\mem[0][20] ),
    .A1(\mem[1][20] ),
    .A2(\mem[4][20] ),
    .A3(\mem[5][20] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0459_));
 sky130_fd_sc_hd__o22ai_2 _0758_ (.A1(_0440_),
    .A2(_0458_),
    .B1(_0459_),
    .B2(_0451_),
    .Y(_0460_));
 sky130_fd_sc_hd__mux4_1 _0759_ (.A0(\mem[12][20] ),
    .A1(\mem[13][20] ),
    .A2(\mem[14][20] ),
    .A3(\mem[15][20] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0461_));
 sky130_fd_sc_hd__mux4_1 _0760_ (.A0(\mem[8][20] ),
    .A1(\mem[9][20] ),
    .A2(\mem[10][20] ),
    .A3(\mem[11][20] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0462_));
 sky130_fd_sc_hd__o22ai_1 _0761_ (.A1(_0444_),
    .A2(_0461_),
    .B1(_0462_),
    .B2(_0455_),
    .Y(_0463_));
 sky130_fd_sc_hd__nor2_1 _0762_ (.A(_0460_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__mux2_1 _0763_ (.A0(_0464_),
    .A1(\last_valid_data[20] ),
    .S(_0432_),
    .X(_0049_));
 sky130_fd_sc_hd__mux4_1 _0764_ (.A0(\mem[2][21] ),
    .A1(\mem[3][21] ),
    .A2(\mem[6][21] ),
    .A3(\mem[7][21] ),
    .S0(_0389_),
    .S1(_0397_),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_1 _0765_ (.A0(\mem[0][21] ),
    .A1(\mem[1][21] ),
    .A2(\mem[4][21] ),
    .A3(\mem[5][21] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0466_));
 sky130_fd_sc_hd__o22ai_1 _0766_ (.A1(_0440_),
    .A2(_0465_),
    .B1(_0466_),
    .B2(_0451_),
    .Y(_0467_));
 sky130_fd_sc_hd__mux4_1 _0767_ (.A0(\mem[12][21] ),
    .A1(\mem[13][21] ),
    .A2(\mem[14][21] ),
    .A3(\mem[15][21] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0468_));
 sky130_fd_sc_hd__mux4_1 _0768_ (.A0(\mem[8][21] ),
    .A1(\mem[9][21] ),
    .A2(\mem[10][21] ),
    .A3(\mem[11][21] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0469_));
 sky130_fd_sc_hd__o22ai_1 _0769_ (.A1(_0444_),
    .A2(_0468_),
    .B1(_0469_),
    .B2(_0455_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_1 _0770_ (.A(_0467_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(_0471_),
    .A1(\last_valid_data[21] ),
    .S(_0432_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_6 _0772_ (.A(_0340_),
    .X(_0472_));
 sky130_fd_sc_hd__mux4_1 _0773_ (.A0(\mem[2][22] ),
    .A1(\mem[3][22] ),
    .A2(\mem[6][22] ),
    .A3(\mem[7][22] ),
    .S0(_0472_),
    .S1(_0397_),
    .X(_0473_));
 sky130_fd_sc_hd__mux4_1 _0774_ (.A0(\mem[0][22] ),
    .A1(\mem[1][22] ),
    .A2(\mem[4][22] ),
    .A3(\mem[5][22] ),
    .S0(_0399_),
    .S1(_0407_),
    .X(_0474_));
 sky130_fd_sc_hd__o22ai_1 _0775_ (.A1(_0440_),
    .A2(_0473_),
    .B1(_0474_),
    .B2(_0451_),
    .Y(_0475_));
 sky130_fd_sc_hd__mux4_1 _0776_ (.A0(\mem[12][22] ),
    .A1(\mem[13][22] ),
    .A2(\mem[14][22] ),
    .A3(\mem[15][22] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0476_));
 sky130_fd_sc_hd__mux4_1 _0777_ (.A0(\mem[8][22] ),
    .A1(\mem[9][22] ),
    .A2(\mem[10][22] ),
    .A3(\mem[11][22] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0477_));
 sky130_fd_sc_hd__o22ai_1 _0778_ (.A1(_0444_),
    .A2(_0476_),
    .B1(_0477_),
    .B2(_0455_),
    .Y(_0478_));
 sky130_fd_sc_hd__nor2_1 _0779_ (.A(_0475_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__mux2_1 _0780_ (.A0(_0479_),
    .A1(\last_valid_data[22] ),
    .S(_0432_),
    .X(_0051_));
 sky130_fd_sc_hd__buf_4 _0781_ (.A(_0304_),
    .X(_0480_));
 sky130_fd_sc_hd__mux4_1 _0782_ (.A0(\mem[2][23] ),
    .A1(\mem[3][23] ),
    .A2(\mem[6][23] ),
    .A3(\mem[7][23] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_8 _0783_ (.A(_0348_),
    .X(_0482_));
 sky130_fd_sc_hd__mux4_1 _0784_ (.A0(\mem[0][23] ),
    .A1(\mem[1][23] ),
    .A2(\mem[4][23] ),
    .A3(\mem[5][23] ),
    .S0(_0482_),
    .S1(_0407_),
    .X(_0483_));
 sky130_fd_sc_hd__o22ai_1 _0785_ (.A1(_0440_),
    .A2(_0481_),
    .B1(_0483_),
    .B2(_0451_),
    .Y(_0484_));
 sky130_fd_sc_hd__mux4_1 _0786_ (.A0(\mem[12][23] ),
    .A1(\mem[13][23] ),
    .A2(\mem[14][23] ),
    .A3(\mem[15][23] ),
    .S0(_0410_),
    .S1(_0411_),
    .X(_0485_));
 sky130_fd_sc_hd__mux4_1 _0787_ (.A0(\mem[8][23] ),
    .A1(\mem[9][23] ),
    .A2(\mem[10][23] ),
    .A3(\mem[11][23] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0486_));
 sky130_fd_sc_hd__o22ai_1 _0788_ (.A1(_0444_),
    .A2(_0485_),
    .B1(_0486_),
    .B2(_0455_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_1 _0789_ (.A(_0484_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(_0488_),
    .A1(\last_valid_data[23] ),
    .S(_0432_),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_1 _0791_ (.A0(\mem[2][24] ),
    .A1(\mem[3][24] ),
    .A2(\mem[6][24] ),
    .A3(\mem[7][24] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_6 _0792_ (.A(_0304_),
    .X(_0490_));
 sky130_fd_sc_hd__mux4_1 _0793_ (.A0(\mem[0][24] ),
    .A1(\mem[1][24] ),
    .A2(\mem[4][24] ),
    .A3(\mem[5][24] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o22ai_1 _0794_ (.A1(_0440_),
    .A2(_0489_),
    .B1(_0491_),
    .B2(_0451_),
    .Y(_0492_));
 sky130_fd_sc_hd__buf_6 _0795_ (.A(_0348_),
    .X(_0493_));
 sky130_fd_sc_hd__buf_6 _0796_ (.A(_0301_),
    .X(_0494_));
 sky130_fd_sc_hd__mux4_1 _0797_ (.A0(\mem[12][24] ),
    .A1(\mem[13][24] ),
    .A2(\mem[14][24] ),
    .A3(\mem[15][24] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0080_));
 sky130_fd_sc_hd__mux4_1 _0798_ (.A0(\mem[8][24] ),
    .A1(\mem[9][24] ),
    .A2(\mem[10][24] ),
    .A3(\mem[11][24] ),
    .S0(_0420_),
    .S1(_0421_),
    .X(_0081_));
 sky130_fd_sc_hd__o22ai_1 _0799_ (.A1(_0444_),
    .A2(_0080_),
    .B1(_0081_),
    .B2(_0455_),
    .Y(_0082_));
 sky130_fd_sc_hd__nor2_1 _0800_ (.A(_0492_),
    .B(_0082_),
    .Y(_0083_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(_0083_),
    .A1(\last_valid_data[24] ),
    .S(_0432_),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _0802_ (.A0(\mem[2][25] ),
    .A1(\mem[3][25] ),
    .A2(\mem[6][25] ),
    .A3(\mem[7][25] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0084_));
 sky130_fd_sc_hd__mux4_1 _0803_ (.A0(\mem[0][25] ),
    .A1(\mem[1][25] ),
    .A2(\mem[4][25] ),
    .A3(\mem[5][25] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0085_));
 sky130_fd_sc_hd__o22ai_1 _0804_ (.A1(_0440_),
    .A2(_0084_),
    .B1(_0085_),
    .B2(_0451_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux4_1 _0805_ (.A0(\mem[12][25] ),
    .A1(\mem[13][25] ),
    .A2(\mem[14][25] ),
    .A3(\mem[15][25] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0087_));
 sky130_fd_sc_hd__buf_4 _0806_ (.A(_0348_),
    .X(_0088_));
 sky130_fd_sc_hd__buf_4 _0807_ (.A(_0302_),
    .X(_0089_));
 sky130_fd_sc_hd__mux4_1 _0808_ (.A0(\mem[8][25] ),
    .A1(\mem[9][25] ),
    .A2(\mem[10][25] ),
    .A3(\mem[11][25] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__o22ai_1 _0809_ (.A1(_0444_),
    .A2(_0087_),
    .B1(_0090_),
    .B2(_0455_),
    .Y(_0091_));
 sky130_fd_sc_hd__nor2_1 _0810_ (.A(_0086_),
    .B(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__mux2_1 _0811_ (.A0(_0092_),
    .A1(\last_valid_data[25] ),
    .S(_0432_),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _0812_ (.A0(\mem[2][26] ),
    .A1(\mem[3][26] ),
    .A2(\mem[6][26] ),
    .A3(\mem[7][26] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _0813_ (.A0(\mem[0][26] ),
    .A1(\mem[1][26] ),
    .A2(\mem[4][26] ),
    .A3(\mem[5][26] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0094_));
 sky130_fd_sc_hd__o22ai_1 _0814_ (.A1(_0440_),
    .A2(_0093_),
    .B1(_0094_),
    .B2(_0451_),
    .Y(_0095_));
 sky130_fd_sc_hd__mux4_1 _0815_ (.A0(\mem[12][26] ),
    .A1(\mem[13][26] ),
    .A2(\mem[14][26] ),
    .A3(\mem[15][26] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0096_));
 sky130_fd_sc_hd__mux4_1 _0816_ (.A0(\mem[8][26] ),
    .A1(\mem[9][26] ),
    .A2(\mem[10][26] ),
    .A3(\mem[11][26] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0097_));
 sky130_fd_sc_hd__o22ai_2 _0817_ (.A1(_0444_),
    .A2(_0096_),
    .B1(_0097_),
    .B2(_0455_),
    .Y(_0098_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(_0095_),
    .B(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__buf_6 _0819_ (.A(_0359_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(_0099_),
    .A1(\last_valid_data[26] ),
    .S(_0100_),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _0821_ (.A0(\mem[2][27] ),
    .A1(\mem[3][27] ),
    .A2(\mem[6][27] ),
    .A3(\mem[7][27] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0101_));
 sky130_fd_sc_hd__mux4_1 _0822_ (.A0(\mem[0][27] ),
    .A1(\mem[1][27] ),
    .A2(\mem[4][27] ),
    .A3(\mem[5][27] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0102_));
 sky130_fd_sc_hd__o22ai_1 _0823_ (.A1(_0440_),
    .A2(_0101_),
    .B1(_0102_),
    .B2(_0451_),
    .Y(_0103_));
 sky130_fd_sc_hd__mux4_1 _0824_ (.A0(\mem[12][27] ),
    .A1(\mem[13][27] ),
    .A2(\mem[14][27] ),
    .A3(\mem[15][27] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0104_));
 sky130_fd_sc_hd__mux4_1 _0825_ (.A0(\mem[8][27] ),
    .A1(\mem[9][27] ),
    .A2(\mem[10][27] ),
    .A3(\mem[11][27] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0105_));
 sky130_fd_sc_hd__o22ai_1 _0826_ (.A1(_0444_),
    .A2(_0104_),
    .B1(_0105_),
    .B2(_0455_),
    .Y(_0106_));
 sky130_fd_sc_hd__nor2_1 _0827_ (.A(_0103_),
    .B(_0106_),
    .Y(_0107_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(_0107_),
    .A1(\last_valid_data[27] ),
    .S(_0100_),
    .X(_0056_));
 sky130_fd_sc_hd__buf_4 _0829_ (.A(_0346_),
    .X(_0108_));
 sky130_fd_sc_hd__mux4_1 _0830_ (.A0(\mem[2][28] ),
    .A1(\mem[3][28] ),
    .A2(\mem[6][28] ),
    .A3(\mem[7][28] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0109_));
 sky130_fd_sc_hd__mux4_1 _0831_ (.A0(\mem[0][28] ),
    .A1(\mem[1][28] ),
    .A2(\mem[4][28] ),
    .A3(\mem[5][28] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0110_));
 sky130_fd_sc_hd__o22ai_1 _0832_ (.A1(_0108_),
    .A2(_0109_),
    .B1(_0110_),
    .B2(_0451_),
    .Y(_0111_));
 sky130_fd_sc_hd__buf_4 _0833_ (.A(_0354_),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_1 _0834_ (.A0(\mem[12][28] ),
    .A1(\mem[13][28] ),
    .A2(\mem[14][28] ),
    .A3(\mem[15][28] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0113_));
 sky130_fd_sc_hd__mux4_1 _0835_ (.A0(\mem[8][28] ),
    .A1(\mem[9][28] ),
    .A2(\mem[10][28] ),
    .A3(\mem[11][28] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0114_));
 sky130_fd_sc_hd__o22ai_1 _0836_ (.A1(_0112_),
    .A2(_0113_),
    .B1(_0114_),
    .B2(_0455_),
    .Y(_0115_));
 sky130_fd_sc_hd__nor2_1 _0837_ (.A(_0111_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(_0116_),
    .A1(\last_valid_data[28] ),
    .S(_0100_),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _0839_ (.A0(\mem[2][29] ),
    .A1(\mem[3][29] ),
    .A2(\mem[6][29] ),
    .A3(\mem[7][29] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0117_));
 sky130_fd_sc_hd__mux4_1 _0840_ (.A0(\mem[0][29] ),
    .A1(\mem[1][29] ),
    .A2(\mem[4][29] ),
    .A3(\mem[5][29] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_8 _0841_ (.A(_0345_),
    .X(_0119_));
 sky130_fd_sc_hd__o22ai_1 _0842_ (.A1(_0108_),
    .A2(_0117_),
    .B1(_0118_),
    .B2(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__mux4_1 _0843_ (.A0(\mem[12][29] ),
    .A1(\mem[13][29] ),
    .A2(\mem[14][29] ),
    .A3(\mem[15][29] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0121_));
 sky130_fd_sc_hd__mux4_1 _0844_ (.A0(\mem[8][29] ),
    .A1(\mem[9][29] ),
    .A2(\mem[10][29] ),
    .A3(\mem[11][29] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0122_));
 sky130_fd_sc_hd__buf_4 _0845_ (.A(_0353_),
    .X(_0123_));
 sky130_fd_sc_hd__o22ai_1 _0846_ (.A1(_0112_),
    .A2(_0121_),
    .B1(_0122_),
    .B2(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0120_),
    .B(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(_0125_),
    .A1(\last_valid_data[29] ),
    .S(_0100_),
    .X(_0058_));
 sky130_fd_sc_hd__mux4_1 _0849_ (.A0(\mem[2][2] ),
    .A1(\mem[3][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0126_));
 sky130_fd_sc_hd__mux4_1 _0850_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[4][2] ),
    .A3(\mem[5][2] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0127_));
 sky130_fd_sc_hd__o22ai_1 _0851_ (.A1(_0108_),
    .A2(_0126_),
    .B1(_0127_),
    .B2(_0119_),
    .Y(_0128_));
 sky130_fd_sc_hd__mux4_1 _0852_ (.A0(\mem[12][2] ),
    .A1(\mem[13][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0129_));
 sky130_fd_sc_hd__mux4_1 _0853_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0130_));
 sky130_fd_sc_hd__o22ai_1 _0854_ (.A1(_0112_),
    .A2(_0129_),
    .B1(_0130_),
    .B2(_0123_),
    .Y(_0131_));
 sky130_fd_sc_hd__nor2_1 _0855_ (.A(_0128_),
    .B(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(_0132_),
    .A1(\last_valid_data[2] ),
    .S(_0100_),
    .X(_0059_));
 sky130_fd_sc_hd__mux4_1 _0857_ (.A0(\mem[2][30] ),
    .A1(\mem[3][30] ),
    .A2(\mem[6][30] ),
    .A3(\mem[7][30] ),
    .S0(_0472_),
    .S1(_0480_),
    .X(_0133_));
 sky130_fd_sc_hd__mux4_1 _0858_ (.A0(\mem[0][30] ),
    .A1(\mem[1][30] ),
    .A2(\mem[4][30] ),
    .A3(\mem[5][30] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0134_));
 sky130_fd_sc_hd__o22ai_1 _0859_ (.A1(_0108_),
    .A2(_0133_),
    .B1(_0134_),
    .B2(_0119_),
    .Y(_0135_));
 sky130_fd_sc_hd__mux4_1 _0860_ (.A0(\mem[12][30] ),
    .A1(\mem[13][30] ),
    .A2(\mem[14][30] ),
    .A3(\mem[15][30] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0136_));
 sky130_fd_sc_hd__mux4_1 _0861_ (.A0(\mem[8][30] ),
    .A1(\mem[9][30] ),
    .A2(\mem[10][30] ),
    .A3(\mem[11][30] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0137_));
 sky130_fd_sc_hd__o22ai_1 _0862_ (.A1(_0112_),
    .A2(_0136_),
    .B1(_0137_),
    .B2(_0123_),
    .Y(_0138_));
 sky130_fd_sc_hd__nor2_1 _0863_ (.A(_0135_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(_0139_),
    .A1(\last_valid_data[30] ),
    .S(_0100_),
    .X(_0060_));
 sky130_fd_sc_hd__mux4_1 _0865_ (.A0(\mem[2][31] ),
    .A1(\mem[3][31] ),
    .A2(\mem[6][31] ),
    .A3(\mem[7][31] ),
    .S0(_0341_),
    .S1(_0480_),
    .X(_0140_));
 sky130_fd_sc_hd__mux4_1 _0866_ (.A0(\mem[0][31] ),
    .A1(\mem[1][31] ),
    .A2(\mem[4][31] ),
    .A3(\mem[5][31] ),
    .S0(_0482_),
    .S1(_0490_),
    .X(_0141_));
 sky130_fd_sc_hd__o22ai_1 _0867_ (.A1(_0108_),
    .A2(_0140_),
    .B1(_0141_),
    .B2(_0119_),
    .Y(_0142_));
 sky130_fd_sc_hd__mux4_1 _0868_ (.A0(\mem[12][31] ),
    .A1(\mem[13][31] ),
    .A2(\mem[14][31] ),
    .A3(\mem[15][31] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0143_));
 sky130_fd_sc_hd__mux4_1 _0869_ (.A0(\mem[8][31] ),
    .A1(\mem[9][31] ),
    .A2(\mem[10][31] ),
    .A3(\mem[11][31] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0144_));
 sky130_fd_sc_hd__o22ai_1 _0870_ (.A1(_0112_),
    .A2(_0143_),
    .B1(_0144_),
    .B2(_0123_),
    .Y(_0145_));
 sky130_fd_sc_hd__nor2_1 _0871_ (.A(_0142_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__mux2_1 _0872_ (.A0(_0146_),
    .A1(\last_valid_data[31] ),
    .S(_0100_),
    .X(_0061_));
 sky130_fd_sc_hd__mux4_1 _0873_ (.A0(\mem[2][3] ),
    .A1(\mem[3][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0147_));
 sky130_fd_sc_hd__mux4_1 _0874_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[4][3] ),
    .A3(\mem[5][3] ),
    .S0(_0361_),
    .S1(_0490_),
    .X(_0148_));
 sky130_fd_sc_hd__o22ai_1 _0875_ (.A1(_0108_),
    .A2(_0147_),
    .B1(_0148_),
    .B2(_0119_),
    .Y(_0149_));
 sky130_fd_sc_hd__mux4_1 _0876_ (.A0(\mem[12][3] ),
    .A1(\mem[13][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_0493_),
    .S1(_0494_),
    .X(_0150_));
 sky130_fd_sc_hd__mux4_1 _0877_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0151_));
 sky130_fd_sc_hd__o22ai_1 _0878_ (.A1(_0112_),
    .A2(_0150_),
    .B1(_0151_),
    .B2(_0123_),
    .Y(_0152_));
 sky130_fd_sc_hd__nor2_1 _0879_ (.A(_0149_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(_0153_),
    .A1(\last_valid_data[3] ),
    .S(_0100_),
    .X(_0062_));
 sky130_fd_sc_hd__mux4_1 _0881_ (.A0(\mem[2][4] ),
    .A1(\mem[3][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0154_));
 sky130_fd_sc_hd__mux4_1 _0882_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[4][4] ),
    .A3(\mem[5][4] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0155_));
 sky130_fd_sc_hd__o22ai_1 _0883_ (.A1(_0108_),
    .A2(_0154_),
    .B1(_0155_),
    .B2(_0119_),
    .Y(_0156_));
 sky130_fd_sc_hd__mux4_1 _0884_ (.A0(\mem[12][4] ),
    .A1(\mem[13][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0157_));
 sky130_fd_sc_hd__mux4_1 _0885_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[11][4] ),
    .S0(_0088_),
    .S1(_0089_),
    .X(_0158_));
 sky130_fd_sc_hd__o22ai_1 _0886_ (.A1(_0112_),
    .A2(_0157_),
    .B1(_0158_),
    .B2(_0123_),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _0887_ (.A(_0156_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(_0160_),
    .A1(\last_valid_data[4] ),
    .S(_0100_),
    .X(_0063_));
 sky130_fd_sc_hd__mux4_1 _0889_ (.A0(\mem[2][5] ),
    .A1(\mem[3][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0161_));
 sky130_fd_sc_hd__mux4_1 _0890_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[4][5] ),
    .A3(\mem[5][5] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0162_));
 sky130_fd_sc_hd__o22ai_1 _0891_ (.A1(_0108_),
    .A2(_0161_),
    .B1(_0162_),
    .B2(_0119_),
    .Y(_0163_));
 sky130_fd_sc_hd__mux4_1 _0892_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0164_));
 sky130_fd_sc_hd__mux4_1 _0893_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0165_));
 sky130_fd_sc_hd__o22ai_1 _0894_ (.A1(_0112_),
    .A2(_0164_),
    .B1(_0165_),
    .B2(_0123_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0163_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(_0167_),
    .A1(\last_valid_data[5] ),
    .S(_0100_),
    .X(_0064_));
 sky130_fd_sc_hd__mux4_1 _0897_ (.A0(\mem[2][6] ),
    .A1(\mem[3][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0168_));
 sky130_fd_sc_hd__mux4_1 _0898_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[4][6] ),
    .A3(\mem[5][6] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0169_));
 sky130_fd_sc_hd__o22ai_1 _0899_ (.A1(_0108_),
    .A2(_0168_),
    .B1(_0169_),
    .B2(_0119_),
    .Y(_0170_));
 sky130_fd_sc_hd__mux4_1 _0900_ (.A0(\mem[12][6] ),
    .A1(\mem[13][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0171_));
 sky130_fd_sc_hd__mux4_1 _0901_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[10][6] ),
    .A3(\mem[11][6] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0172_));
 sky130_fd_sc_hd__o22ai_1 _0902_ (.A1(_0112_),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0123_),
    .Y(_0173_));
 sky130_fd_sc_hd__nor2_1 _0903_ (.A(_0170_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(_0174_),
    .A1(\last_valid_data[6] ),
    .S(_0359_),
    .X(_0065_));
 sky130_fd_sc_hd__mux4_1 _0905_ (.A0(\mem[2][7] ),
    .A1(\mem[3][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0175_));
 sky130_fd_sc_hd__mux4_1 _0906_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[4][7] ),
    .A3(\mem[5][7] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0176_));
 sky130_fd_sc_hd__o22ai_1 _0907_ (.A1(_0108_),
    .A2(_0175_),
    .B1(_0176_),
    .B2(_0119_),
    .Y(_0177_));
 sky130_fd_sc_hd__mux4_1 _0908_ (.A0(\mem[12][7] ),
    .A1(\mem[13][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0178_));
 sky130_fd_sc_hd__mux4_1 _0909_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[10][7] ),
    .A3(\mem[11][7] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0179_));
 sky130_fd_sc_hd__o22ai_1 _0910_ (.A1(_0112_),
    .A2(_0178_),
    .B1(_0179_),
    .B2(_0123_),
    .Y(_0180_));
 sky130_fd_sc_hd__nor2_1 _0911_ (.A(_0177_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(_0181_),
    .A1(\last_valid_data[7] ),
    .S(_0359_),
    .X(_0066_));
 sky130_fd_sc_hd__mux4_1 _0913_ (.A0(\mem[2][8] ),
    .A1(\mem[3][8] ),
    .A2(\mem[6][8] ),
    .A3(\mem[7][8] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0182_));
 sky130_fd_sc_hd__mux4_1 _0914_ (.A0(\mem[0][8] ),
    .A1(\mem[1][8] ),
    .A2(\mem[4][8] ),
    .A3(\mem[5][8] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0183_));
 sky130_fd_sc_hd__o22ai_1 _0915_ (.A1(_0346_),
    .A2(_0182_),
    .B1(_0183_),
    .B2(_0119_),
    .Y(_0184_));
 sky130_fd_sc_hd__mux4_1 _0916_ (.A0(\mem[12][8] ),
    .A1(\mem[13][8] ),
    .A2(\mem[14][8] ),
    .A3(\mem[15][8] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0185_));
 sky130_fd_sc_hd__mux4_1 _0917_ (.A0(\mem[8][8] ),
    .A1(\mem[9][8] ),
    .A2(\mem[10][8] ),
    .A3(\mem[11][8] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0186_));
 sky130_fd_sc_hd__o22ai_1 _0918_ (.A1(_0354_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0123_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0919_ (.A(_0184_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(_0188_),
    .A1(\last_valid_data[8] ),
    .S(_0359_),
    .X(_0067_));
 sky130_fd_sc_hd__mux4_1 _0921_ (.A0(\mem[2][9] ),
    .A1(\mem[3][9] ),
    .A2(\mem[6][9] ),
    .A3(\mem[7][9] ),
    .S0(_0341_),
    .S1(_0342_),
    .X(_0189_));
 sky130_fd_sc_hd__mux4_1 _0922_ (.A0(\mem[0][9] ),
    .A1(\mem[1][9] ),
    .A2(\mem[4][9] ),
    .A3(\mem[5][9] ),
    .S0(_0361_),
    .S1(_0362_),
    .X(_0190_));
 sky130_fd_sc_hd__o22ai_1 _0923_ (.A1(_0346_),
    .A2(_0189_),
    .B1(_0190_),
    .B2(_0345_),
    .Y(_0191_));
 sky130_fd_sc_hd__mux4_1 _0924_ (.A0(\mem[12][9] ),
    .A1(\mem[13][9] ),
    .A2(\mem[14][9] ),
    .A3(\mem[15][9] ),
    .S0(_0364_),
    .S1(_0302_),
    .X(_0192_));
 sky130_fd_sc_hd__mux4_1 _0925_ (.A0(\mem[8][9] ),
    .A1(\mem[9][9] ),
    .A2(\mem[10][9] ),
    .A3(\mem[11][9] ),
    .S0(_0368_),
    .S1(_0369_),
    .X(_0193_));
 sky130_fd_sc_hd__o22ai_1 _0926_ (.A1(_0354_),
    .A2(_0192_),
    .B1(_0193_),
    .B2(_0353_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _0927_ (.A(_0191_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(_0195_),
    .A1(\last_valid_data[9] ),
    .S(_0359_),
    .X(_0068_));
 sky130_fd_sc_hd__buf_2 _0929_ (.A(last_valid_data_available),
    .X(_0196_));
 sky130_fd_sc_hd__nand2b_1 _0930_ (.A_N(_0196_),
    .B(_0360_),
    .Y(_0069_));
 sky130_fd_sc_hd__xnor2_1 _0931_ (.A(_0349_),
    .B(_0360_),
    .Y(_0070_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(_0019_),
    .A1(_0303_),
    .S(_0359_),
    .X(_0071_));
 sky130_fd_sc_hd__nand3_1 _0933_ (.A(_0293_),
    .B(_0506_),
    .C(_0325_),
    .Y(_0197_));
 sky130_fd_sc_hd__xnor2_1 _0934_ (.A(_0305_),
    .B(_0197_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand3_1 _0935_ (.A(_0349_),
    .B(_0303_),
    .C(_0305_),
    .Y(_0198_));
 sky130_fd_sc_hd__nor3_1 _0936_ (.A(_0327_),
    .B(net43),
    .C(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__xnor2_1 _0937_ (.A(_0498_),
    .B(_0199_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand3_1 _0938_ (.A(_0305_),
    .B(\rd_ptr[3] ),
    .C(_0506_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor3_1 _0939_ (.A(_0327_),
    .B(net43),
    .C(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__xor2_1 _0940_ (.A(\rd_ptr[4] ),
    .B(_0201_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2b_1 _0941_ (.A_N(net61),
    .B(net35),
    .Y(_0202_));
 sky130_fd_sc_hd__xnor2_1 _0942_ (.A(\wr_ptr[0] ),
    .B(_0202_),
    .Y(_0075_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(_0018_),
    .A1(\wr_ptr[1] ),
    .S(_0202_),
    .X(_0076_));
 sky130_fd_sc_hd__nand3b_1 _0944_ (.A_N(net61),
    .B(_0514_),
    .C(net35),
    .Y(_0203_));
 sky130_fd_sc_hd__xnor2_1 _0945_ (.A(\wr_ptr[2] ),
    .B(_0203_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor4_1 _0946_ (.A(_0508_),
    .B(_0017_),
    .C(net61),
    .D(_0298_),
    .Y(_0204_));
 sky130_fd_sc_hd__xor2_1 _0947_ (.A(\wr_ptr[3] ),
    .B(_0204_),
    .X(_0078_));
 sky130_fd_sc_hd__nand2b_1 _0948_ (.A_N(net61),
    .B(_0007_),
    .Y(_0205_));
 sky130_fd_sc_hd__xnor2_1 _0949_ (.A(\wr_ptr[4] ),
    .B(_0205_),
    .Y(_0079_));
 sky130_fd_sc_hd__xor2_1 _0950_ (.A(_0517_),
    .B(net39),
    .X(_0206_));
 sky130_fd_sc_hd__nor4_1 _0951_ (.A(net40),
    .B(net41),
    .C(net42),
    .D(_0206_),
    .Y(net36));
 sky130_fd_sc_hd__a31o_1 _0952_ (.A1(net39),
    .A2(net40),
    .A3(net41),
    .B1(net42),
    .X(net37));
 sky130_fd_sc_hd__and2_0 _0953_ (.A(net35),
    .B(net61),
    .X(net62));
 sky130_fd_sc_hd__buf_4 _0954_ (.A(_0291_),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_8 _0955_ (.A(_0196_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _0956_ (.A(_0208_),
    .B(\last_valid_data[0] ),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _0957_ (.A(net95),
    .B(_0358_),
    .Y(_0210_));
 sky130_fd_sc_hd__o21ai_0 _0958_ (.A1(_0207_),
    .A2(_0209_),
    .B1(_0210_),
    .Y(net63));
 sky130_fd_sc_hd__nand2_1 _0959_ (.A(_0208_),
    .B(\last_valid_data[10] ),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _0960_ (.A(net95),
    .B(_0374_),
    .Y(_0212_));
 sky130_fd_sc_hd__o21ai_0 _0961_ (.A1(_0207_),
    .A2(_0211_),
    .B1(_0212_),
    .Y(net64));
 sky130_fd_sc_hd__nand2_1 _0962_ (.A(_0208_),
    .B(\last_valid_data[11] ),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _0963_ (.A(net95),
    .B(_0381_),
    .Y(_0214_));
 sky130_fd_sc_hd__o21ai_0 _0964_ (.A1(_0207_),
    .A2(_0213_),
    .B1(_0214_),
    .Y(net65));
 sky130_fd_sc_hd__nand2_1 _0965_ (.A(_0208_),
    .B(\last_valid_data[12] ),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _0966_ (.A(net95),
    .B(_0388_),
    .Y(_0216_));
 sky130_fd_sc_hd__o21ai_0 _0967_ (.A1(_0207_),
    .A2(_0215_),
    .B1(_0216_),
    .Y(net66));
 sky130_fd_sc_hd__nand2_1 _0968_ (.A(_0208_),
    .B(\last_valid_data[13] ),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _0969_ (.A(net95),
    .B(_0396_),
    .Y(_0218_));
 sky130_fd_sc_hd__o21ai_0 _0970_ (.A1(_0207_),
    .A2(_0217_),
    .B1(_0218_),
    .Y(net67));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(_0208_),
    .B(\last_valid_data[14] ),
    .Y(_0219_));
 sky130_fd_sc_hd__nand2_1 _0972_ (.A(net95),
    .B(_0405_),
    .Y(_0220_));
 sky130_fd_sc_hd__o21ai_0 _0973_ (.A1(_0207_),
    .A2(_0219_),
    .B1(_0220_),
    .Y(net68));
 sky130_fd_sc_hd__nand2_1 _0974_ (.A(_0208_),
    .B(\last_valid_data[15] ),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(net95),
    .B(_0415_),
    .Y(_0222_));
 sky130_fd_sc_hd__o21ai_0 _0976_ (.A1(_0207_),
    .A2(_0221_),
    .B1(_0222_),
    .Y(net69));
 sky130_fd_sc_hd__buf_6 _0977_ (.A(_0291_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _0978_ (.A(_0208_),
    .B(\last_valid_data[16] ),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(net95),
    .B(_0424_),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_1 _0980_ (.A1(_0223_),
    .A2(_0224_),
    .B1(_0225_),
    .Y(net70));
 sky130_fd_sc_hd__nand2_1 _0981_ (.A(_0208_),
    .B(\last_valid_data[17] ),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _0982_ (.A(net95),
    .B(_0431_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_1 _0983_ (.A1(_0223_),
    .A2(_0226_),
    .B1(_0227_),
    .Y(net71));
 sky130_fd_sc_hd__nand2_1 _0984_ (.A(_0208_),
    .B(\last_valid_data[18] ),
    .Y(_0228_));
 sky130_fd_sc_hd__buf_6 _0985_ (.A(_0325_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0986_ (.A(_0229_),
    .B(_0439_),
    .Y(_0230_));
 sky130_fd_sc_hd__o21ai_0 _0987_ (.A1(_0223_),
    .A2(_0228_),
    .B1(_0230_),
    .Y(net72));
 sky130_fd_sc_hd__buf_6 _0988_ (.A(_0196_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _0989_ (.A(_0231_),
    .B(\last_valid_data[19] ),
    .Y(_0232_));
 sky130_fd_sc_hd__nand2_1 _0990_ (.A(_0229_),
    .B(_0448_),
    .Y(_0233_));
 sky130_fd_sc_hd__o21ai_0 _0991_ (.A1(_0223_),
    .A2(_0232_),
    .B1(_0233_),
    .Y(net73));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(_0231_),
    .B(\last_valid_data[1] ),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0229_),
    .B(_0457_),
    .Y(_0235_));
 sky130_fd_sc_hd__o21ai_0 _0994_ (.A1(_0223_),
    .A2(_0234_),
    .B1(_0235_),
    .Y(net74));
 sky130_fd_sc_hd__nand2_1 _0995_ (.A(_0231_),
    .B(\last_valid_data[20] ),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0229_),
    .B(_0464_),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_0 _0997_ (.A1(_0223_),
    .A2(_0236_),
    .B1(_0237_),
    .Y(net75));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(_0231_),
    .B(\last_valid_data[21] ),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _0999_ (.A(_0229_),
    .B(_0471_),
    .Y(_0239_));
 sky130_fd_sc_hd__o21ai_0 _1000_ (.A1(_0223_),
    .A2(_0238_),
    .B1(_0239_),
    .Y(net76));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0231_),
    .B(\last_valid_data[22] ),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(_0229_),
    .B(_0479_),
    .Y(_0241_));
 sky130_fd_sc_hd__o21ai_0 _1003_ (.A1(_0223_),
    .A2(_0240_),
    .B1(_0241_),
    .Y(net77));
 sky130_fd_sc_hd__nand2_1 _1004_ (.A(_0231_),
    .B(\last_valid_data[23] ),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(_0229_),
    .B(_0488_),
    .Y(_0243_));
 sky130_fd_sc_hd__o21ai_0 _1006_ (.A1(_0223_),
    .A2(_0242_),
    .B1(_0243_),
    .Y(net78));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0231_),
    .B(\last_valid_data[24] ),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(_0229_),
    .B(_0083_),
    .Y(_0245_));
 sky130_fd_sc_hd__o21ai_1 _1009_ (.A1(_0223_),
    .A2(_0244_),
    .B1(_0245_),
    .Y(net79));
 sky130_fd_sc_hd__buf_4 _1010_ (.A(_0291_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _1011_ (.A(_0231_),
    .B(\last_valid_data[25] ),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _1012_ (.A(_0229_),
    .B(_0092_),
    .Y(_0248_));
 sky130_fd_sc_hd__o21ai_0 _1013_ (.A1(_0246_),
    .A2(_0247_),
    .B1(_0248_),
    .Y(net80));
 sky130_fd_sc_hd__nand2_1 _1014_ (.A(_0231_),
    .B(\last_valid_data[26] ),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(_0229_),
    .B(_0099_),
    .Y(_0250_));
 sky130_fd_sc_hd__o21ai_1 _1016_ (.A1(_0246_),
    .A2(_0249_),
    .B1(_0250_),
    .Y(net81));
 sky130_fd_sc_hd__nand2_1 _1017_ (.A(_0231_),
    .B(\last_valid_data[27] ),
    .Y(_0251_));
 sky130_fd_sc_hd__buf_4 _1018_ (.A(_0292_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _1019_ (.A(_0252_),
    .B(_0107_),
    .Y(_0253_));
 sky130_fd_sc_hd__o21ai_0 _1020_ (.A1(_0246_),
    .A2(_0251_),
    .B1(_0253_),
    .Y(net82));
 sky130_fd_sc_hd__buf_4 _1021_ (.A(_0196_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _1022_ (.A(_0254_),
    .B(\last_valid_data[28] ),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _1023_ (.A(_0252_),
    .B(_0116_),
    .Y(_0256_));
 sky130_fd_sc_hd__o21ai_0 _1024_ (.A1(_0246_),
    .A2(_0255_),
    .B1(_0256_),
    .Y(net83));
 sky130_fd_sc_hd__nand2_1 _1025_ (.A(_0254_),
    .B(\last_valid_data[29] ),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _1026_ (.A(_0252_),
    .B(_0125_),
    .Y(_0258_));
 sky130_fd_sc_hd__o21ai_0 _1027_ (.A1(_0246_),
    .A2(_0257_),
    .B1(_0258_),
    .Y(net84));
 sky130_fd_sc_hd__nand2_1 _1028_ (.A(_0254_),
    .B(\last_valid_data[2] ),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _1029_ (.A(_0252_),
    .B(_0132_),
    .Y(_0260_));
 sky130_fd_sc_hd__o21ai_0 _1030_ (.A1(_0246_),
    .A2(_0259_),
    .B1(_0260_),
    .Y(net85));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(_0254_),
    .B(\last_valid_data[30] ),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(_0252_),
    .B(_0139_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_0 _1033_ (.A1(_0246_),
    .A2(_0261_),
    .B1(_0262_),
    .Y(net86));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(_0254_),
    .B(\last_valid_data[31] ),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _1035_ (.A(_0252_),
    .B(_0146_),
    .Y(_0264_));
 sky130_fd_sc_hd__o21ai_0 _1036_ (.A1(_0246_),
    .A2(_0263_),
    .B1(_0264_),
    .Y(net87));
 sky130_fd_sc_hd__nand2_1 _1037_ (.A(_0254_),
    .B(\last_valid_data[3] ),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _1038_ (.A(_0252_),
    .B(_0153_),
    .Y(_0266_));
 sky130_fd_sc_hd__o21ai_0 _1039_ (.A1(_0246_),
    .A2(_0265_),
    .B1(_0266_),
    .Y(net88));
 sky130_fd_sc_hd__nand2_1 _1040_ (.A(_0254_),
    .B(\last_valid_data[4] ),
    .Y(_0267_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(_0252_),
    .B(_0160_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_1 _1042_ (.A1(_0246_),
    .A2(_0267_),
    .B1(_0268_),
    .Y(net89));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0254_),
    .B(\last_valid_data[5] ),
    .Y(_0269_));
 sky130_fd_sc_hd__nand2_1 _1044_ (.A(_0252_),
    .B(_0167_),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_0 _1045_ (.A1(_0325_),
    .A2(_0269_),
    .B1(_0270_),
    .Y(net90));
 sky130_fd_sc_hd__nand2_1 _1046_ (.A(_0254_),
    .B(\last_valid_data[6] ),
    .Y(_0271_));
 sky130_fd_sc_hd__nand2_1 _1047_ (.A(_0252_),
    .B(_0174_),
    .Y(_0272_));
 sky130_fd_sc_hd__o21ai_0 _1048_ (.A1(_0325_),
    .A2(_0271_),
    .B1(_0272_),
    .Y(net91));
 sky130_fd_sc_hd__nand2_1 _1049_ (.A(_0254_),
    .B(\last_valid_data[7] ),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _1050_ (.A(_0207_),
    .B(_0181_),
    .Y(_0274_));
 sky130_fd_sc_hd__o21ai_0 _1051_ (.A1(_0325_),
    .A2(_0273_),
    .B1(_0274_),
    .Y(net92));
 sky130_fd_sc_hd__nand2_1 _1052_ (.A(_0196_),
    .B(\last_valid_data[8] ),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_1 _1053_ (.A(_0207_),
    .B(_0188_),
    .Y(_0276_));
 sky130_fd_sc_hd__o21ai_1 _1054_ (.A1(_0325_),
    .A2(_0275_),
    .B1(_0276_),
    .Y(net93));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0196_),
    .B(\last_valid_data[9] ),
    .Y(_0277_));
 sky130_fd_sc_hd__nand2_1 _1056_ (.A(_0207_),
    .B(_0195_),
    .Y(_0278_));
 sky130_fd_sc_hd__o21ai_1 _1057_ (.A1(_0325_),
    .A2(_0277_),
    .B1(_0278_),
    .Y(net94));
 sky130_fd_sc_hd__inv_1 _1058_ (.A(net61),
    .Y(net97));
 sky130_fd_sc_hd__fa_2 _1059_ (.A(_0495_),
    .B(\wr_ptr[1] ),
    .CIN(_0496_),
    .COUT(_0497_),
    .SUM(net39));
 sky130_fd_sc_hd__ha_1 _1060_ (.A(_0498_),
    .B(\wr_ptr[3] ),
    .COUT(_0499_),
    .SUM(_0500_));
 sky130_fd_sc_hd__ha_1 _1061_ (.A(_0495_),
    .B(\wr_ptr[1] ),
    .COUT(_0501_),
    .SUM(_0502_));
 sky130_fd_sc_hd__ha_1 _1062_ (.A(_0503_),
    .B(\wr_ptr[2] ),
    .COUT(_0504_),
    .SUM(_0505_));
 sky130_fd_sc_hd__ha_1 _1063_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_0506_),
    .SUM(_0019_));
 sky130_fd_sc_hd__ha_1 _1064_ (.A(net44),
    .B(net51),
    .COUT(_0507_),
    .SUM(_0020_));
 sky130_fd_sc_hd__ha_1 _1065_ (.A(_0017_),
    .B(_0508_),
    .COUT(_0509_),
    .SUM(_0018_));
 sky130_fd_sc_hd__ha_1 _1066_ (.A(_0017_),
    .B(\wr_ptr[1] ),
    .COUT(_0510_),
    .SUM(_0511_));
 sky130_fd_sc_hd__ha_1 _1067_ (.A(\wr_ptr[0] ),
    .B(_0508_),
    .COUT(_0512_),
    .SUM(_0513_));
 sky130_fd_sc_hd__ha_1 _1068_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_0514_),
    .SUM(_0515_));
 sky130_fd_sc_hd__ha_1 _1069_ (.A(\rd_ptr[0] ),
    .B(_0017_),
    .COUT(_0516_),
    .SUM(_0517_));
 sky130_fd_sc_hd__dfrtp_2 \error_count[0]$_DFFE_PN0P_  (.D(_0021_),
    .Q(net44),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[10]$_DFFE_PN0P_  (.D(_0022_),
    .Q(net45),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[11]$_DFFE_PN0P_  (.D(_0023_),
    .Q(net46),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[12]$_DFFE_PN0P_  (.D(_0024_),
    .Q(net47),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[13]$_DFFE_PN0P_  (.D(_0025_),
    .Q(net48),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[14]$_DFFE_PN0P_  (.D(_0026_),
    .Q(net49),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[15]$_DFFE_PN0P_  (.D(_0027_),
    .Q(net50),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[1]$_DFFE_PN0P_  (.D(_0028_),
    .Q(net51),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[2]$_DFFE_PN0P_  (.D(_0029_),
    .Q(net52),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[3]$_DFFE_PN0P_  (.D(_0030_),
    .Q(net53),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[4]$_DFFE_PN0P_  (.D(_0031_),
    .Q(net54),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_2 \error_count[5]$_DFFE_PN0P_  (.D(_0032_),
    .Q(net55),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[6]$_DFFE_PN0P_  (.D(_0033_),
    .Q(net56),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[7]$_DFFE_PN0P_  (.D(_0034_),
    .Q(net57),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[8]$_DFFE_PN0P_  (.D(_0035_),
    .Q(net58),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_count[9]$_DFFE_PN0P_  (.D(_0036_),
    .Q(net59),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \error_detected$_DFF_PN0_  (.D(_0000_),
    .Q(net60),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[0]$_DFFE_PN0P_  (.D(_0037_),
    .Q(\last_valid_data[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[10]$_DFFE_PN0P_  (.D(_0038_),
    .Q(\last_valid_data[10] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[11]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\last_valid_data[11] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[12]$_DFFE_PN0P_  (.D(_0040_),
    .Q(\last_valid_data[12] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[13]$_DFFE_PN0P_  (.D(_0041_),
    .Q(\last_valid_data[13] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[14]$_DFFE_PN0P_  (.D(_0042_),
    .Q(\last_valid_data[14] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[15]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\last_valid_data[15] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[16]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\last_valid_data[16] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[17]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\last_valid_data[17] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[18]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\last_valid_data[18] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[19]$_DFFE_PN0P_  (.D(_0047_),
    .Q(\last_valid_data[19] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[1]$_DFFE_PN0P_  (.D(_0048_),
    .Q(\last_valid_data[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[20]$_DFFE_PN0P_  (.D(_0049_),
    .Q(\last_valid_data[20] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[21]$_DFFE_PN0P_  (.D(_0050_),
    .Q(\last_valid_data[21] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[22]$_DFFE_PN0P_  (.D(_0051_),
    .Q(\last_valid_data[22] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[23]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\last_valid_data[23] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[24]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\last_valid_data[24] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[25]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\last_valid_data[25] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[26]$_DFFE_PN0P_  (.D(_0055_),
    .Q(\last_valid_data[26] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[27]$_DFFE_PN0P_  (.D(_0056_),
    .Q(\last_valid_data[27] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[28]$_DFFE_PN0P_  (.D(_0057_),
    .Q(\last_valid_data[28] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[29]$_DFFE_PN0P_  (.D(_0058_),
    .Q(\last_valid_data[29] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[2]$_DFFE_PN0P_  (.D(_0059_),
    .Q(\last_valid_data[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[30]$_DFFE_PN0P_  (.D(_0060_),
    .Q(\last_valid_data[30] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[31]$_DFFE_PN0P_  (.D(_0061_),
    .Q(\last_valid_data[31] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[3]$_DFFE_PN0P_  (.D(_0062_),
    .Q(\last_valid_data[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[4]$_DFFE_PN0P_  (.D(_0063_),
    .Q(\last_valid_data[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[5]$_DFFE_PN0P_  (.D(_0064_),
    .Q(\last_valid_data[5] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[6]$_DFFE_PN0P_  (.D(_0065_),
    .Q(\last_valid_data[6] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[7]$_DFFE_PN0P_  (.D(_0066_),
    .Q(\last_valid_data[7] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[8]$_DFFE_PN0P_  (.D(_0067_),
    .Q(\last_valid_data[8] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data[9]$_DFFE_PN0P_  (.D(_0068_),
    .Q(\last_valid_data[9] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \last_valid_data_available$_DFFE_PN0P_  (.D(_0069_),
    .Q(last_valid_data_available),
    .RESET_B(net1),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net3),
    .DE(_0001_),
    .Q(\mem[0][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][10]$_DFFE_PP_  (.D(net4),
    .DE(_0001_),
    .Q(\mem[0][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][11]$_DFFE_PP_  (.D(net5),
    .DE(_0001_),
    .Q(\mem[0][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][12]$_DFFE_PP_  (.D(net6),
    .DE(_0001_),
    .Q(\mem[0][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][13]$_DFFE_PP_  (.D(net7),
    .DE(_0001_),
    .Q(\mem[0][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][14]$_DFFE_PP_  (.D(net8),
    .DE(_0001_),
    .Q(\mem[0][14] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][15]$_DFFE_PP_  (.D(net9),
    .DE(_0001_),
    .Q(\mem[0][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][16]$_DFFE_PP_  (.D(net10),
    .DE(_0001_),
    .Q(\mem[0][16] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][17]$_DFFE_PP_  (.D(net11),
    .DE(_0001_),
    .Q(\mem[0][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][18]$_DFFE_PP_  (.D(net12),
    .DE(_0001_),
    .Q(\mem[0][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][19]$_DFFE_PP_  (.D(net13),
    .DE(_0001_),
    .Q(\mem[0][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net14),
    .DE(_0001_),
    .Q(\mem[0][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][20]$_DFFE_PP_  (.D(net15),
    .DE(_0001_),
    .Q(\mem[0][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][21]$_DFFE_PP_  (.D(net16),
    .DE(_0001_),
    .Q(\mem[0][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][22]$_DFFE_PP_  (.D(net17),
    .DE(_0001_),
    .Q(\mem[0][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][23]$_DFFE_PP_  (.D(net18),
    .DE(_0001_),
    .Q(\mem[0][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][24]$_DFFE_PP_  (.D(net19),
    .DE(_0001_),
    .Q(\mem[0][24] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][25]$_DFFE_PP_  (.D(net20),
    .DE(_0001_),
    .Q(\mem[0][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][26]$_DFFE_PP_  (.D(net21),
    .DE(_0001_),
    .Q(\mem[0][26] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][27]$_DFFE_PP_  (.D(net22),
    .DE(_0001_),
    .Q(\mem[0][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][28]$_DFFE_PP_  (.D(net23),
    .DE(_0001_),
    .Q(\mem[0][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][29]$_DFFE_PP_  (.D(net24),
    .DE(_0001_),
    .Q(\mem[0][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net25),
    .DE(_0001_),
    .Q(\mem[0][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][30]$_DFFE_PP_  (.D(net26),
    .DE(_0001_),
    .Q(\mem[0][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][31]$_DFFE_PP_  (.D(net27),
    .DE(_0001_),
    .Q(\mem[0][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net28),
    .DE(_0001_),
    .Q(\mem[0][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net29),
    .DE(_0001_),
    .Q(\mem[0][4] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net30),
    .DE(_0001_),
    .Q(\mem[0][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net31),
    .DE(_0001_),
    .Q(\mem[0][6] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net32),
    .DE(_0001_),
    .Q(\mem[0][7] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][8]$_DFFE_PP_  (.D(net33),
    .DE(_0001_),
    .Q(\mem[0][8] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][9]$_DFFE_PP_  (.D(net34),
    .DE(_0001_),
    .Q(\mem[0][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net3),
    .DE(_0002_),
    .Q(\mem[10][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][10]$_DFFE_PP_  (.D(net4),
    .DE(_0002_),
    .Q(\mem[10][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][11]$_DFFE_PP_  (.D(net5),
    .DE(_0002_),
    .Q(\mem[10][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][12]$_DFFE_PP_  (.D(net6),
    .DE(_0002_),
    .Q(\mem[10][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][13]$_DFFE_PP_  (.D(net7),
    .DE(_0002_),
    .Q(\mem[10][13] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][14]$_DFFE_PP_  (.D(net8),
    .DE(_0002_),
    .Q(\mem[10][14] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][15]$_DFFE_PP_  (.D(net9),
    .DE(_0002_),
    .Q(\mem[10][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][16]$_DFFE_PP_  (.D(net10),
    .DE(_0002_),
    .Q(\mem[10][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][17]$_DFFE_PP_  (.D(net11),
    .DE(_0002_),
    .Q(\mem[10][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][18]$_DFFE_PP_  (.D(net12),
    .DE(_0002_),
    .Q(\mem[10][18] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][19]$_DFFE_PP_  (.D(net13),
    .DE(_0002_),
    .Q(\mem[10][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net14),
    .DE(_0002_),
    .Q(\mem[10][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][20]$_DFFE_PP_  (.D(net15),
    .DE(_0002_),
    .Q(\mem[10][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][21]$_DFFE_PP_  (.D(net16),
    .DE(_0002_),
    .Q(\mem[10][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][22]$_DFFE_PP_  (.D(net17),
    .DE(_0002_),
    .Q(\mem[10][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][23]$_DFFE_PP_  (.D(net18),
    .DE(_0002_),
    .Q(\mem[10][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][24]$_DFFE_PP_  (.D(net19),
    .DE(_0002_),
    .Q(\mem[10][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][25]$_DFFE_PP_  (.D(net20),
    .DE(_0002_),
    .Q(\mem[10][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][26]$_DFFE_PP_  (.D(net21),
    .DE(_0002_),
    .Q(\mem[10][26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][27]$_DFFE_PP_  (.D(net22),
    .DE(_0002_),
    .Q(\mem[10][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][28]$_DFFE_PP_  (.D(net23),
    .DE(_0002_),
    .Q(\mem[10][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][29]$_DFFE_PP_  (.D(net24),
    .DE(_0002_),
    .Q(\mem[10][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net25),
    .DE(_0002_),
    .Q(\mem[10][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][30]$_DFFE_PP_  (.D(net26),
    .DE(_0002_),
    .Q(\mem[10][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][31]$_DFFE_PP_  (.D(net27),
    .DE(_0002_),
    .Q(\mem[10][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net28),
    .DE(_0002_),
    .Q(\mem[10][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net29),
    .DE(_0002_),
    .Q(\mem[10][4] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net30),
    .DE(_0002_),
    .Q(\mem[10][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net31),
    .DE(_0002_),
    .Q(\mem[10][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net32),
    .DE(_0002_),
    .Q(\mem[10][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][8]$_DFFE_PP_  (.D(net33),
    .DE(_0002_),
    .Q(\mem[10][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][9]$_DFFE_PP_  (.D(net34),
    .DE(_0002_),
    .Q(\mem[10][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net3),
    .DE(_0003_),
    .Q(\mem[11][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][10]$_DFFE_PP_  (.D(net4),
    .DE(_0003_),
    .Q(\mem[11][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][11]$_DFFE_PP_  (.D(net5),
    .DE(_0003_),
    .Q(\mem[11][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][12]$_DFFE_PP_  (.D(net6),
    .DE(_0003_),
    .Q(\mem[11][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][13]$_DFFE_PP_  (.D(net7),
    .DE(_0003_),
    .Q(\mem[11][13] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][14]$_DFFE_PP_  (.D(net8),
    .DE(_0003_),
    .Q(\mem[11][14] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][15]$_DFFE_PP_  (.D(net9),
    .DE(_0003_),
    .Q(\mem[11][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][16]$_DFFE_PP_  (.D(net10),
    .DE(_0003_),
    .Q(\mem[11][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][17]$_DFFE_PP_  (.D(net11),
    .DE(_0003_),
    .Q(\mem[11][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][18]$_DFFE_PP_  (.D(net12),
    .DE(_0003_),
    .Q(\mem[11][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][19]$_DFFE_PP_  (.D(net13),
    .DE(_0003_),
    .Q(\mem[11][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net14),
    .DE(_0003_),
    .Q(\mem[11][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][20]$_DFFE_PP_  (.D(net15),
    .DE(_0003_),
    .Q(\mem[11][20] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][21]$_DFFE_PP_  (.D(net16),
    .DE(_0003_),
    .Q(\mem[11][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][22]$_DFFE_PP_  (.D(net17),
    .DE(_0003_),
    .Q(\mem[11][22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][23]$_DFFE_PP_  (.D(net18),
    .DE(_0003_),
    .Q(\mem[11][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][24]$_DFFE_PP_  (.D(net19),
    .DE(_0003_),
    .Q(\mem[11][24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][25]$_DFFE_PP_  (.D(net20),
    .DE(_0003_),
    .Q(\mem[11][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][26]$_DFFE_PP_  (.D(net21),
    .DE(_0003_),
    .Q(\mem[11][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][27]$_DFFE_PP_  (.D(net22),
    .DE(_0003_),
    .Q(\mem[11][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][28]$_DFFE_PP_  (.D(net23),
    .DE(_0003_),
    .Q(\mem[11][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][29]$_DFFE_PP_  (.D(net24),
    .DE(_0003_),
    .Q(\mem[11][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net25),
    .DE(_0003_),
    .Q(\mem[11][2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][30]$_DFFE_PP_  (.D(net26),
    .DE(_0003_),
    .Q(\mem[11][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][31]$_DFFE_PP_  (.D(net27),
    .DE(_0003_),
    .Q(\mem[11][31] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net28),
    .DE(_0003_),
    .Q(\mem[11][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net29),
    .DE(_0003_),
    .Q(\mem[11][4] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net30),
    .DE(_0003_),
    .Q(\mem[11][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net31),
    .DE(_0003_),
    .Q(\mem[11][6] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net32),
    .DE(_0003_),
    .Q(\mem[11][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][8]$_DFFE_PP_  (.D(net33),
    .DE(_0003_),
    .Q(\mem[11][8] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][9]$_DFFE_PP_  (.D(net34),
    .DE(_0003_),
    .Q(\mem[11][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net3),
    .DE(_0004_),
    .Q(\mem[12][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][10]$_DFFE_PP_  (.D(net4),
    .DE(_0004_),
    .Q(\mem[12][10] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][11]$_DFFE_PP_  (.D(net5),
    .DE(_0004_),
    .Q(\mem[12][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][12]$_DFFE_PP_  (.D(net6),
    .DE(_0004_),
    .Q(\mem[12][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][13]$_DFFE_PP_  (.D(net7),
    .DE(_0004_),
    .Q(\mem[12][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][14]$_DFFE_PP_  (.D(net8),
    .DE(_0004_),
    .Q(\mem[12][14] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][15]$_DFFE_PP_  (.D(net9),
    .DE(_0004_),
    .Q(\mem[12][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][16]$_DFFE_PP_  (.D(net10),
    .DE(_0004_),
    .Q(\mem[12][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][17]$_DFFE_PP_  (.D(net11),
    .DE(_0004_),
    .Q(\mem[12][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][18]$_DFFE_PP_  (.D(net12),
    .DE(_0004_),
    .Q(\mem[12][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][19]$_DFFE_PP_  (.D(net13),
    .DE(_0004_),
    .Q(\mem[12][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net14),
    .DE(_0004_),
    .Q(\mem[12][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][20]$_DFFE_PP_  (.D(net15),
    .DE(_0004_),
    .Q(\mem[12][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][21]$_DFFE_PP_  (.D(net16),
    .DE(_0004_),
    .Q(\mem[12][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][22]$_DFFE_PP_  (.D(net17),
    .DE(_0004_),
    .Q(\mem[12][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][23]$_DFFE_PP_  (.D(net18),
    .DE(_0004_),
    .Q(\mem[12][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][24]$_DFFE_PP_  (.D(net19),
    .DE(_0004_),
    .Q(\mem[12][24] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][25]$_DFFE_PP_  (.D(net20),
    .DE(_0004_),
    .Q(\mem[12][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][26]$_DFFE_PP_  (.D(net21),
    .DE(_0004_),
    .Q(\mem[12][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][27]$_DFFE_PP_  (.D(net22),
    .DE(_0004_),
    .Q(\mem[12][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][28]$_DFFE_PP_  (.D(net23),
    .DE(_0004_),
    .Q(\mem[12][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][29]$_DFFE_PP_  (.D(net24),
    .DE(_0004_),
    .Q(\mem[12][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net25),
    .DE(_0004_),
    .Q(\mem[12][2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][30]$_DFFE_PP_  (.D(net26),
    .DE(_0004_),
    .Q(\mem[12][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][31]$_DFFE_PP_  (.D(net27),
    .DE(_0004_),
    .Q(\mem[12][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net28),
    .DE(_0004_),
    .Q(\mem[12][3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net29),
    .DE(_0004_),
    .Q(\mem[12][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net30),
    .DE(_0004_),
    .Q(\mem[12][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net31),
    .DE(_0004_),
    .Q(\mem[12][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net32),
    .DE(_0004_),
    .Q(\mem[12][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][8]$_DFFE_PP_  (.D(net33),
    .DE(_0004_),
    .Q(\mem[12][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][9]$_DFFE_PP_  (.D(net34),
    .DE(_0004_),
    .Q(\mem[12][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net3),
    .DE(_0005_),
    .Q(\mem[13][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][10]$_DFFE_PP_  (.D(net4),
    .DE(_0005_),
    .Q(\mem[13][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][11]$_DFFE_PP_  (.D(net5),
    .DE(_0005_),
    .Q(\mem[13][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][12]$_DFFE_PP_  (.D(net6),
    .DE(_0005_),
    .Q(\mem[13][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][13]$_DFFE_PP_  (.D(net7),
    .DE(_0005_),
    .Q(\mem[13][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][14]$_DFFE_PP_  (.D(net8),
    .DE(_0005_),
    .Q(\mem[13][14] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][15]$_DFFE_PP_  (.D(net9),
    .DE(_0005_),
    .Q(\mem[13][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][16]$_DFFE_PP_  (.D(net10),
    .DE(_0005_),
    .Q(\mem[13][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][17]$_DFFE_PP_  (.D(net11),
    .DE(_0005_),
    .Q(\mem[13][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][18]$_DFFE_PP_  (.D(net12),
    .DE(_0005_),
    .Q(\mem[13][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][19]$_DFFE_PP_  (.D(net13),
    .DE(_0005_),
    .Q(\mem[13][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net14),
    .DE(_0005_),
    .Q(\mem[13][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][20]$_DFFE_PP_  (.D(net15),
    .DE(_0005_),
    .Q(\mem[13][20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][21]$_DFFE_PP_  (.D(net16),
    .DE(_0005_),
    .Q(\mem[13][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][22]$_DFFE_PP_  (.D(net17),
    .DE(_0005_),
    .Q(\mem[13][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][23]$_DFFE_PP_  (.D(net18),
    .DE(_0005_),
    .Q(\mem[13][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][24]$_DFFE_PP_  (.D(net19),
    .DE(_0005_),
    .Q(\mem[13][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][25]$_DFFE_PP_  (.D(net20),
    .DE(_0005_),
    .Q(\mem[13][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][26]$_DFFE_PP_  (.D(net21),
    .DE(_0005_),
    .Q(\mem[13][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][27]$_DFFE_PP_  (.D(net22),
    .DE(_0005_),
    .Q(\mem[13][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][28]$_DFFE_PP_  (.D(net23),
    .DE(_0005_),
    .Q(\mem[13][28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][29]$_DFFE_PP_  (.D(net24),
    .DE(_0005_),
    .Q(\mem[13][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net25),
    .DE(_0005_),
    .Q(\mem[13][2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][30]$_DFFE_PP_  (.D(net26),
    .DE(_0005_),
    .Q(\mem[13][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][31]$_DFFE_PP_  (.D(net27),
    .DE(_0005_),
    .Q(\mem[13][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net28),
    .DE(_0005_),
    .Q(\mem[13][3] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net29),
    .DE(_0005_),
    .Q(\mem[13][4] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net30),
    .DE(_0005_),
    .Q(\mem[13][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net31),
    .DE(_0005_),
    .Q(\mem[13][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net32),
    .DE(_0005_),
    .Q(\mem[13][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][8]$_DFFE_PP_  (.D(net33),
    .DE(_0005_),
    .Q(\mem[13][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][9]$_DFFE_PP_  (.D(net34),
    .DE(_0005_),
    .Q(\mem[13][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net3),
    .DE(_0006_),
    .Q(\mem[14][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][10]$_DFFE_PP_  (.D(net4),
    .DE(_0006_),
    .Q(\mem[14][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][11]$_DFFE_PP_  (.D(net5),
    .DE(_0006_),
    .Q(\mem[14][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][12]$_DFFE_PP_  (.D(net6),
    .DE(_0006_),
    .Q(\mem[14][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][13]$_DFFE_PP_  (.D(net7),
    .DE(_0006_),
    .Q(\mem[14][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][14]$_DFFE_PP_  (.D(net8),
    .DE(_0006_),
    .Q(\mem[14][14] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][15]$_DFFE_PP_  (.D(net9),
    .DE(_0006_),
    .Q(\mem[14][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][16]$_DFFE_PP_  (.D(net10),
    .DE(_0006_),
    .Q(\mem[14][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][17]$_DFFE_PP_  (.D(net11),
    .DE(_0006_),
    .Q(\mem[14][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][18]$_DFFE_PP_  (.D(net12),
    .DE(_0006_),
    .Q(\mem[14][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][19]$_DFFE_PP_  (.D(net13),
    .DE(_0006_),
    .Q(\mem[14][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net14),
    .DE(_0006_),
    .Q(\mem[14][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][20]$_DFFE_PP_  (.D(net15),
    .DE(_0006_),
    .Q(\mem[14][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][21]$_DFFE_PP_  (.D(net16),
    .DE(_0006_),
    .Q(\mem[14][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][22]$_DFFE_PP_  (.D(net17),
    .DE(_0006_),
    .Q(\mem[14][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][23]$_DFFE_PP_  (.D(net18),
    .DE(_0006_),
    .Q(\mem[14][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][24]$_DFFE_PP_  (.D(net19),
    .DE(_0006_),
    .Q(\mem[14][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][25]$_DFFE_PP_  (.D(net20),
    .DE(_0006_),
    .Q(\mem[14][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][26]$_DFFE_PP_  (.D(net21),
    .DE(_0006_),
    .Q(\mem[14][26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][27]$_DFFE_PP_  (.D(net22),
    .DE(_0006_),
    .Q(\mem[14][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][28]$_DFFE_PP_  (.D(net23),
    .DE(_0006_),
    .Q(\mem[14][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][29]$_DFFE_PP_  (.D(net24),
    .DE(_0006_),
    .Q(\mem[14][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net25),
    .DE(_0006_),
    .Q(\mem[14][2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][30]$_DFFE_PP_  (.D(net26),
    .DE(_0006_),
    .Q(\mem[14][30] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][31]$_DFFE_PP_  (.D(net27),
    .DE(_0006_),
    .Q(\mem[14][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net28),
    .DE(_0006_),
    .Q(\mem[14][3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net29),
    .DE(_0006_),
    .Q(\mem[14][4] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net30),
    .DE(_0006_),
    .Q(\mem[14][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net31),
    .DE(_0006_),
    .Q(\mem[14][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net32),
    .DE(_0006_),
    .Q(\mem[14][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][8]$_DFFE_PP_  (.D(net33),
    .DE(_0006_),
    .Q(\mem[14][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][9]$_DFFE_PP_  (.D(net34),
    .DE(_0006_),
    .Q(\mem[14][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net3),
    .DE(_0007_),
    .Q(\mem[15][0] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][10]$_DFFE_PP_  (.D(net4),
    .DE(_0007_),
    .Q(\mem[15][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][11]$_DFFE_PP_  (.D(net5),
    .DE(_0007_),
    .Q(\mem[15][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][12]$_DFFE_PP_  (.D(net6),
    .DE(_0007_),
    .Q(\mem[15][12] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][13]$_DFFE_PP_  (.D(net7),
    .DE(_0007_),
    .Q(\mem[15][13] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][14]$_DFFE_PP_  (.D(net8),
    .DE(_0007_),
    .Q(\mem[15][14] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][15]$_DFFE_PP_  (.D(net9),
    .DE(_0007_),
    .Q(\mem[15][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][16]$_DFFE_PP_  (.D(net10),
    .DE(_0007_),
    .Q(\mem[15][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][17]$_DFFE_PP_  (.D(net11),
    .DE(_0007_),
    .Q(\mem[15][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][18]$_DFFE_PP_  (.D(net12),
    .DE(_0007_),
    .Q(\mem[15][18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][19]$_DFFE_PP_  (.D(net13),
    .DE(_0007_),
    .Q(\mem[15][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net14),
    .DE(_0007_),
    .Q(\mem[15][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][20]$_DFFE_PP_  (.D(net15),
    .DE(_0007_),
    .Q(\mem[15][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][21]$_DFFE_PP_  (.D(net16),
    .DE(_0007_),
    .Q(\mem[15][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][22]$_DFFE_PP_  (.D(net17),
    .DE(_0007_),
    .Q(\mem[15][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][23]$_DFFE_PP_  (.D(net18),
    .DE(_0007_),
    .Q(\mem[15][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][24]$_DFFE_PP_  (.D(net19),
    .DE(_0007_),
    .Q(\mem[15][24] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][25]$_DFFE_PP_  (.D(net20),
    .DE(_0007_),
    .Q(\mem[15][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][26]$_DFFE_PP_  (.D(net21),
    .DE(_0007_),
    .Q(\mem[15][26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][27]$_DFFE_PP_  (.D(net22),
    .DE(_0007_),
    .Q(\mem[15][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][28]$_DFFE_PP_  (.D(net23),
    .DE(_0007_),
    .Q(\mem[15][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][29]$_DFFE_PP_  (.D(net24),
    .DE(_0007_),
    .Q(\mem[15][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net25),
    .DE(_0007_),
    .Q(\mem[15][2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][30]$_DFFE_PP_  (.D(net26),
    .DE(_0007_),
    .Q(\mem[15][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][31]$_DFFE_PP_  (.D(net27),
    .DE(_0007_),
    .Q(\mem[15][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net28),
    .DE(_0007_),
    .Q(\mem[15][3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net29),
    .DE(_0007_),
    .Q(\mem[15][4] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net30),
    .DE(_0007_),
    .Q(\mem[15][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net31),
    .DE(_0007_),
    .Q(\mem[15][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net32),
    .DE(_0007_),
    .Q(\mem[15][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][8]$_DFFE_PP_  (.D(net33),
    .DE(_0007_),
    .Q(\mem[15][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][9]$_DFFE_PP_  (.D(net34),
    .DE(_0007_),
    .Q(\mem[15][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net3),
    .DE(_0008_),
    .Q(\mem[1][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][10]$_DFFE_PP_  (.D(net4),
    .DE(_0008_),
    .Q(\mem[1][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][11]$_DFFE_PP_  (.D(net5),
    .DE(_0008_),
    .Q(\mem[1][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][12]$_DFFE_PP_  (.D(net6),
    .DE(_0008_),
    .Q(\mem[1][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][13]$_DFFE_PP_  (.D(net7),
    .DE(_0008_),
    .Q(\mem[1][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][14]$_DFFE_PP_  (.D(net8),
    .DE(_0008_),
    .Q(\mem[1][14] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][15]$_DFFE_PP_  (.D(net9),
    .DE(_0008_),
    .Q(\mem[1][15] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][16]$_DFFE_PP_  (.D(net10),
    .DE(_0008_),
    .Q(\mem[1][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][17]$_DFFE_PP_  (.D(net11),
    .DE(_0008_),
    .Q(\mem[1][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][18]$_DFFE_PP_  (.D(net12),
    .DE(_0008_),
    .Q(\mem[1][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][19]$_DFFE_PP_  (.D(net13),
    .DE(_0008_),
    .Q(\mem[1][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net14),
    .DE(_0008_),
    .Q(\mem[1][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][20]$_DFFE_PP_  (.D(net15),
    .DE(_0008_),
    .Q(\mem[1][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][21]$_DFFE_PP_  (.D(net16),
    .DE(_0008_),
    .Q(\mem[1][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][22]$_DFFE_PP_  (.D(net17),
    .DE(_0008_),
    .Q(\mem[1][22] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][23]$_DFFE_PP_  (.D(net18),
    .DE(_0008_),
    .Q(\mem[1][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][24]$_DFFE_PP_  (.D(net19),
    .DE(_0008_),
    .Q(\mem[1][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][25]$_DFFE_PP_  (.D(net20),
    .DE(_0008_),
    .Q(\mem[1][25] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][26]$_DFFE_PP_  (.D(net21),
    .DE(_0008_),
    .Q(\mem[1][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][27]$_DFFE_PP_  (.D(net22),
    .DE(_0008_),
    .Q(\mem[1][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][28]$_DFFE_PP_  (.D(net23),
    .DE(_0008_),
    .Q(\mem[1][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][29]$_DFFE_PP_  (.D(net24),
    .DE(_0008_),
    .Q(\mem[1][29] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net25),
    .DE(_0008_),
    .Q(\mem[1][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][30]$_DFFE_PP_  (.D(net26),
    .DE(_0008_),
    .Q(\mem[1][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][31]$_DFFE_PP_  (.D(net27),
    .DE(_0008_),
    .Q(\mem[1][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net28),
    .DE(_0008_),
    .Q(\mem[1][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net29),
    .DE(_0008_),
    .Q(\mem[1][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net30),
    .DE(_0008_),
    .Q(\mem[1][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net31),
    .DE(_0008_),
    .Q(\mem[1][6] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net32),
    .DE(_0008_),
    .Q(\mem[1][7] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][8]$_DFFE_PP_  (.D(net33),
    .DE(_0008_),
    .Q(\mem[1][8] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][9]$_DFFE_PP_  (.D(net34),
    .DE(_0008_),
    .Q(\mem[1][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net3),
    .DE(_0009_),
    .Q(\mem[2][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][10]$_DFFE_PP_  (.D(net4),
    .DE(_0009_),
    .Q(\mem[2][10] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][11]$_DFFE_PP_  (.D(net5),
    .DE(_0009_),
    .Q(\mem[2][11] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][12]$_DFFE_PP_  (.D(net6),
    .DE(_0009_),
    .Q(\mem[2][12] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][13]$_DFFE_PP_  (.D(net7),
    .DE(_0009_),
    .Q(\mem[2][13] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][14]$_DFFE_PP_  (.D(net8),
    .DE(_0009_),
    .Q(\mem[2][14] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][15]$_DFFE_PP_  (.D(net9),
    .DE(_0009_),
    .Q(\mem[2][15] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][16]$_DFFE_PP_  (.D(net10),
    .DE(_0009_),
    .Q(\mem[2][16] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][17]$_DFFE_PP_  (.D(net11),
    .DE(_0009_),
    .Q(\mem[2][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][18]$_DFFE_PP_  (.D(net12),
    .DE(_0009_),
    .Q(\mem[2][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][19]$_DFFE_PP_  (.D(net13),
    .DE(_0009_),
    .Q(\mem[2][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net14),
    .DE(_0009_),
    .Q(\mem[2][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][20]$_DFFE_PP_  (.D(net15),
    .DE(_0009_),
    .Q(\mem[2][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][21]$_DFFE_PP_  (.D(net16),
    .DE(_0009_),
    .Q(\mem[2][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][22]$_DFFE_PP_  (.D(net17),
    .DE(_0009_),
    .Q(\mem[2][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][23]$_DFFE_PP_  (.D(net18),
    .DE(_0009_),
    .Q(\mem[2][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][24]$_DFFE_PP_  (.D(net19),
    .DE(_0009_),
    .Q(\mem[2][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][25]$_DFFE_PP_  (.D(net20),
    .DE(_0009_),
    .Q(\mem[2][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][26]$_DFFE_PP_  (.D(net21),
    .DE(_0009_),
    .Q(\mem[2][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][27]$_DFFE_PP_  (.D(net22),
    .DE(_0009_),
    .Q(\mem[2][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][28]$_DFFE_PP_  (.D(net23),
    .DE(_0009_),
    .Q(\mem[2][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][29]$_DFFE_PP_  (.D(net24),
    .DE(_0009_),
    .Q(\mem[2][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net25),
    .DE(_0009_),
    .Q(\mem[2][2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][30]$_DFFE_PP_  (.D(net26),
    .DE(_0009_),
    .Q(\mem[2][30] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][31]$_DFFE_PP_  (.D(net27),
    .DE(_0009_),
    .Q(\mem[2][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net28),
    .DE(_0009_),
    .Q(\mem[2][3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net29),
    .DE(_0009_),
    .Q(\mem[2][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net30),
    .DE(_0009_),
    .Q(\mem[2][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net31),
    .DE(_0009_),
    .Q(\mem[2][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net32),
    .DE(_0009_),
    .Q(\mem[2][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][8]$_DFFE_PP_  (.D(net33),
    .DE(_0009_),
    .Q(\mem[2][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][9]$_DFFE_PP_  (.D(net34),
    .DE(_0009_),
    .Q(\mem[2][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net3),
    .DE(_0010_),
    .Q(\mem[3][0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][10]$_DFFE_PP_  (.D(net4),
    .DE(_0010_),
    .Q(\mem[3][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][11]$_DFFE_PP_  (.D(net5),
    .DE(_0010_),
    .Q(\mem[3][11] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][12]$_DFFE_PP_  (.D(net6),
    .DE(_0010_),
    .Q(\mem[3][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][13]$_DFFE_PP_  (.D(net7),
    .DE(_0010_),
    .Q(\mem[3][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][14]$_DFFE_PP_  (.D(net8),
    .DE(_0010_),
    .Q(\mem[3][14] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][15]$_DFFE_PP_  (.D(net9),
    .DE(_0010_),
    .Q(\mem[3][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][16]$_DFFE_PP_  (.D(net10),
    .DE(_0010_),
    .Q(\mem[3][16] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][17]$_DFFE_PP_  (.D(net11),
    .DE(_0010_),
    .Q(\mem[3][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][18]$_DFFE_PP_  (.D(net12),
    .DE(_0010_),
    .Q(\mem[3][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][19]$_DFFE_PP_  (.D(net13),
    .DE(_0010_),
    .Q(\mem[3][19] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net14),
    .DE(_0010_),
    .Q(\mem[3][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][20]$_DFFE_PP_  (.D(net15),
    .DE(_0010_),
    .Q(\mem[3][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][21]$_DFFE_PP_  (.D(net16),
    .DE(_0010_),
    .Q(\mem[3][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][22]$_DFFE_PP_  (.D(net17),
    .DE(_0010_),
    .Q(\mem[3][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][23]$_DFFE_PP_  (.D(net18),
    .DE(_0010_),
    .Q(\mem[3][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][24]$_DFFE_PP_  (.D(net19),
    .DE(_0010_),
    .Q(\mem[3][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][25]$_DFFE_PP_  (.D(net20),
    .DE(_0010_),
    .Q(\mem[3][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][26]$_DFFE_PP_  (.D(net21),
    .DE(_0010_),
    .Q(\mem[3][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][27]$_DFFE_PP_  (.D(net22),
    .DE(_0010_),
    .Q(\mem[3][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][28]$_DFFE_PP_  (.D(net23),
    .DE(_0010_),
    .Q(\mem[3][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][29]$_DFFE_PP_  (.D(net24),
    .DE(_0010_),
    .Q(\mem[3][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net25),
    .DE(_0010_),
    .Q(\mem[3][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][30]$_DFFE_PP_  (.D(net26),
    .DE(_0010_),
    .Q(\mem[3][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][31]$_DFFE_PP_  (.D(net27),
    .DE(_0010_),
    .Q(\mem[3][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net28),
    .DE(_0010_),
    .Q(\mem[3][3] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net29),
    .DE(_0010_),
    .Q(\mem[3][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net30),
    .DE(_0010_),
    .Q(\mem[3][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net31),
    .DE(_0010_),
    .Q(\mem[3][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net32),
    .DE(_0010_),
    .Q(\mem[3][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][8]$_DFFE_PP_  (.D(net33),
    .DE(_0010_),
    .Q(\mem[3][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][9]$_DFFE_PP_  (.D(net34),
    .DE(_0010_),
    .Q(\mem[3][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net3),
    .DE(_0011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][10]$_DFFE_PP_  (.D(net4),
    .DE(_0011_),
    .Q(\mem[4][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][11]$_DFFE_PP_  (.D(net5),
    .DE(_0011_),
    .Q(\mem[4][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][12]$_DFFE_PP_  (.D(net6),
    .DE(_0011_),
    .Q(\mem[4][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][13]$_DFFE_PP_  (.D(net7),
    .DE(_0011_),
    .Q(\mem[4][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][14]$_DFFE_PP_  (.D(net8),
    .DE(_0011_),
    .Q(\mem[4][14] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][15]$_DFFE_PP_  (.D(net9),
    .DE(_0011_),
    .Q(\mem[4][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][16]$_DFFE_PP_  (.D(net10),
    .DE(_0011_),
    .Q(\mem[4][16] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][17]$_DFFE_PP_  (.D(net11),
    .DE(_0011_),
    .Q(\mem[4][17] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][18]$_DFFE_PP_  (.D(net12),
    .DE(_0011_),
    .Q(\mem[4][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][19]$_DFFE_PP_  (.D(net13),
    .DE(_0011_),
    .Q(\mem[4][19] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net14),
    .DE(_0011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][20]$_DFFE_PP_  (.D(net15),
    .DE(_0011_),
    .Q(\mem[4][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][21]$_DFFE_PP_  (.D(net16),
    .DE(_0011_),
    .Q(\mem[4][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][22]$_DFFE_PP_  (.D(net17),
    .DE(_0011_),
    .Q(\mem[4][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][23]$_DFFE_PP_  (.D(net18),
    .DE(_0011_),
    .Q(\mem[4][23] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][24]$_DFFE_PP_  (.D(net19),
    .DE(_0011_),
    .Q(\mem[4][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][25]$_DFFE_PP_  (.D(net20),
    .DE(_0011_),
    .Q(\mem[4][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][26]$_DFFE_PP_  (.D(net21),
    .DE(_0011_),
    .Q(\mem[4][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][27]$_DFFE_PP_  (.D(net22),
    .DE(_0011_),
    .Q(\mem[4][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][28]$_DFFE_PP_  (.D(net23),
    .DE(_0011_),
    .Q(\mem[4][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][29]$_DFFE_PP_  (.D(net24),
    .DE(_0011_),
    .Q(\mem[4][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net25),
    .DE(_0011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][30]$_DFFE_PP_  (.D(net26),
    .DE(_0011_),
    .Q(\mem[4][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][31]$_DFFE_PP_  (.D(net27),
    .DE(_0011_),
    .Q(\mem[4][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net28),
    .DE(_0011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net29),
    .DE(_0011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net30),
    .DE(_0011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net31),
    .DE(_0011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net32),
    .DE(_0011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][8]$_DFFE_PP_  (.D(net33),
    .DE(_0011_),
    .Q(\mem[4][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][9]$_DFFE_PP_  (.D(net34),
    .DE(_0011_),
    .Q(\mem[4][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net3),
    .DE(_0012_),
    .Q(\mem[5][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][10]$_DFFE_PP_  (.D(net4),
    .DE(_0012_),
    .Q(\mem[5][10] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][11]$_DFFE_PP_  (.D(net5),
    .DE(_0012_),
    .Q(\mem[5][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][12]$_DFFE_PP_  (.D(net6),
    .DE(_0012_),
    .Q(\mem[5][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][13]$_DFFE_PP_  (.D(net7),
    .DE(_0012_),
    .Q(\mem[5][13] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][14]$_DFFE_PP_  (.D(net8),
    .DE(_0012_),
    .Q(\mem[5][14] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][15]$_DFFE_PP_  (.D(net9),
    .DE(_0012_),
    .Q(\mem[5][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][16]$_DFFE_PP_  (.D(net10),
    .DE(_0012_),
    .Q(\mem[5][16] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][17]$_DFFE_PP_  (.D(net11),
    .DE(_0012_),
    .Q(\mem[5][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][18]$_DFFE_PP_  (.D(net12),
    .DE(_0012_),
    .Q(\mem[5][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][19]$_DFFE_PP_  (.D(net13),
    .DE(_0012_),
    .Q(\mem[5][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net14),
    .DE(_0012_),
    .Q(\mem[5][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][20]$_DFFE_PP_  (.D(net15),
    .DE(_0012_),
    .Q(\mem[5][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][21]$_DFFE_PP_  (.D(net16),
    .DE(_0012_),
    .Q(\mem[5][21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][22]$_DFFE_PP_  (.D(net17),
    .DE(_0012_),
    .Q(\mem[5][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][23]$_DFFE_PP_  (.D(net18),
    .DE(_0012_),
    .Q(\mem[5][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][24]$_DFFE_PP_  (.D(net19),
    .DE(_0012_),
    .Q(\mem[5][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][25]$_DFFE_PP_  (.D(net20),
    .DE(_0012_),
    .Q(\mem[5][25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][26]$_DFFE_PP_  (.D(net21),
    .DE(_0012_),
    .Q(\mem[5][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][27]$_DFFE_PP_  (.D(net22),
    .DE(_0012_),
    .Q(\mem[5][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][28]$_DFFE_PP_  (.D(net23),
    .DE(_0012_),
    .Q(\mem[5][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][29]$_DFFE_PP_  (.D(net24),
    .DE(_0012_),
    .Q(\mem[5][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net25),
    .DE(_0012_),
    .Q(\mem[5][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][30]$_DFFE_PP_  (.D(net26),
    .DE(_0012_),
    .Q(\mem[5][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][31]$_DFFE_PP_  (.D(net27),
    .DE(_0012_),
    .Q(\mem[5][31] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net28),
    .DE(_0012_),
    .Q(\mem[5][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net29),
    .DE(_0012_),
    .Q(\mem[5][4] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net30),
    .DE(_0012_),
    .Q(\mem[5][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net31),
    .DE(_0012_),
    .Q(\mem[5][6] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net32),
    .DE(_0012_),
    .Q(\mem[5][7] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][8]$_DFFE_PP_  (.D(net33),
    .DE(_0012_),
    .Q(\mem[5][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][9]$_DFFE_PP_  (.D(net34),
    .DE(_0012_),
    .Q(\mem[5][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net3),
    .DE(_0013_),
    .Q(\mem[6][0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][10]$_DFFE_PP_  (.D(net4),
    .DE(_0013_),
    .Q(\mem[6][10] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][11]$_DFFE_PP_  (.D(net5),
    .DE(_0013_),
    .Q(\mem[6][11] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][12]$_DFFE_PP_  (.D(net6),
    .DE(_0013_),
    .Q(\mem[6][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][13]$_DFFE_PP_  (.D(net7),
    .DE(_0013_),
    .Q(\mem[6][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][14]$_DFFE_PP_  (.D(net8),
    .DE(_0013_),
    .Q(\mem[6][14] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][15]$_DFFE_PP_  (.D(net9),
    .DE(_0013_),
    .Q(\mem[6][15] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][16]$_DFFE_PP_  (.D(net10),
    .DE(_0013_),
    .Q(\mem[6][16] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][17]$_DFFE_PP_  (.D(net11),
    .DE(_0013_),
    .Q(\mem[6][17] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][18]$_DFFE_PP_  (.D(net12),
    .DE(_0013_),
    .Q(\mem[6][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][19]$_DFFE_PP_  (.D(net13),
    .DE(_0013_),
    .Q(\mem[6][19] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net14),
    .DE(_0013_),
    .Q(\mem[6][1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][20]$_DFFE_PP_  (.D(net15),
    .DE(_0013_),
    .Q(\mem[6][20] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][21]$_DFFE_PP_  (.D(net16),
    .DE(_0013_),
    .Q(\mem[6][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][22]$_DFFE_PP_  (.D(net17),
    .DE(_0013_),
    .Q(\mem[6][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][23]$_DFFE_PP_  (.D(net18),
    .DE(_0013_),
    .Q(\mem[6][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][24]$_DFFE_PP_  (.D(net19),
    .DE(_0013_),
    .Q(\mem[6][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][25]$_DFFE_PP_  (.D(net20),
    .DE(_0013_),
    .Q(\mem[6][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][26]$_DFFE_PP_  (.D(net21),
    .DE(_0013_),
    .Q(\mem[6][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][27]$_DFFE_PP_  (.D(net22),
    .DE(_0013_),
    .Q(\mem[6][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][28]$_DFFE_PP_  (.D(net23),
    .DE(_0013_),
    .Q(\mem[6][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][29]$_DFFE_PP_  (.D(net24),
    .DE(_0013_),
    .Q(\mem[6][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net25),
    .DE(_0013_),
    .Q(\mem[6][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][30]$_DFFE_PP_  (.D(net26),
    .DE(_0013_),
    .Q(\mem[6][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][31]$_DFFE_PP_  (.D(net27),
    .DE(_0013_),
    .Q(\mem[6][31] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net28),
    .DE(_0013_),
    .Q(\mem[6][3] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net29),
    .DE(_0013_),
    .Q(\mem[6][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net30),
    .DE(_0013_),
    .Q(\mem[6][5] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net31),
    .DE(_0013_),
    .Q(\mem[6][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net32),
    .DE(_0013_),
    .Q(\mem[6][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][8]$_DFFE_PP_  (.D(net33),
    .DE(_0013_),
    .Q(\mem[6][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][9]$_DFFE_PP_  (.D(net34),
    .DE(_0013_),
    .Q(\mem[6][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net3),
    .DE(_0014_),
    .Q(\mem[7][0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][10]$_DFFE_PP_  (.D(net4),
    .DE(_0014_),
    .Q(\mem[7][10] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][11]$_DFFE_PP_  (.D(net5),
    .DE(_0014_),
    .Q(\mem[7][11] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][12]$_DFFE_PP_  (.D(net6),
    .DE(_0014_),
    .Q(\mem[7][12] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][13]$_DFFE_PP_  (.D(net7),
    .DE(_0014_),
    .Q(\mem[7][13] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][14]$_DFFE_PP_  (.D(net8),
    .DE(_0014_),
    .Q(\mem[7][14] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][15]$_DFFE_PP_  (.D(net9),
    .DE(_0014_),
    .Q(\mem[7][15] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][16]$_DFFE_PP_  (.D(net10),
    .DE(_0014_),
    .Q(\mem[7][16] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][17]$_DFFE_PP_  (.D(net11),
    .DE(_0014_),
    .Q(\mem[7][17] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][18]$_DFFE_PP_  (.D(net12),
    .DE(_0014_),
    .Q(\mem[7][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][19]$_DFFE_PP_  (.D(net13),
    .DE(_0014_),
    .Q(\mem[7][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net14),
    .DE(_0014_),
    .Q(\mem[7][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][20]$_DFFE_PP_  (.D(net15),
    .DE(_0014_),
    .Q(\mem[7][20] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][21]$_DFFE_PP_  (.D(net16),
    .DE(_0014_),
    .Q(\mem[7][21] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][22]$_DFFE_PP_  (.D(net17),
    .DE(_0014_),
    .Q(\mem[7][22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][23]$_DFFE_PP_  (.D(net18),
    .DE(_0014_),
    .Q(\mem[7][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][24]$_DFFE_PP_  (.D(net19),
    .DE(_0014_),
    .Q(\mem[7][24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][25]$_DFFE_PP_  (.D(net20),
    .DE(_0014_),
    .Q(\mem[7][25] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][26]$_DFFE_PP_  (.D(net21),
    .DE(_0014_),
    .Q(\mem[7][26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][27]$_DFFE_PP_  (.D(net22),
    .DE(_0014_),
    .Q(\mem[7][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][28]$_DFFE_PP_  (.D(net23),
    .DE(_0014_),
    .Q(\mem[7][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][29]$_DFFE_PP_  (.D(net24),
    .DE(_0014_),
    .Q(\mem[7][29] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net25),
    .DE(_0014_),
    .Q(\mem[7][2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][30]$_DFFE_PP_  (.D(net26),
    .DE(_0014_),
    .Q(\mem[7][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][31]$_DFFE_PP_  (.D(net27),
    .DE(_0014_),
    .Q(\mem[7][31] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net28),
    .DE(_0014_),
    .Q(\mem[7][3] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net29),
    .DE(_0014_),
    .Q(\mem[7][4] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net30),
    .DE(_0014_),
    .Q(\mem[7][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net31),
    .DE(_0014_),
    .Q(\mem[7][6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net32),
    .DE(_0014_),
    .Q(\mem[7][7] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][8]$_DFFE_PP_  (.D(net33),
    .DE(_0014_),
    .Q(\mem[7][8] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][9]$_DFFE_PP_  (.D(net34),
    .DE(_0014_),
    .Q(\mem[7][9] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net3),
    .DE(_0015_),
    .Q(\mem[8][0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][10]$_DFFE_PP_  (.D(net4),
    .DE(_0015_),
    .Q(\mem[8][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][11]$_DFFE_PP_  (.D(net5),
    .DE(_0015_),
    .Q(\mem[8][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][12]$_DFFE_PP_  (.D(net6),
    .DE(_0015_),
    .Q(\mem[8][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][13]$_DFFE_PP_  (.D(net7),
    .DE(_0015_),
    .Q(\mem[8][13] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][14]$_DFFE_PP_  (.D(net8),
    .DE(_0015_),
    .Q(\mem[8][14] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][15]$_DFFE_PP_  (.D(net9),
    .DE(_0015_),
    .Q(\mem[8][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][16]$_DFFE_PP_  (.D(net10),
    .DE(_0015_),
    .Q(\mem[8][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][17]$_DFFE_PP_  (.D(net11),
    .DE(_0015_),
    .Q(\mem[8][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][18]$_DFFE_PP_  (.D(net12),
    .DE(_0015_),
    .Q(\mem[8][18] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][19]$_DFFE_PP_  (.D(net13),
    .DE(_0015_),
    .Q(\mem[8][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net14),
    .DE(_0015_),
    .Q(\mem[8][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][20]$_DFFE_PP_  (.D(net15),
    .DE(_0015_),
    .Q(\mem[8][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][21]$_DFFE_PP_  (.D(net16),
    .DE(_0015_),
    .Q(\mem[8][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][22]$_DFFE_PP_  (.D(net17),
    .DE(_0015_),
    .Q(\mem[8][22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][23]$_DFFE_PP_  (.D(net18),
    .DE(_0015_),
    .Q(\mem[8][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][24]$_DFFE_PP_  (.D(net19),
    .DE(_0015_),
    .Q(\mem[8][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][25]$_DFFE_PP_  (.D(net20),
    .DE(_0015_),
    .Q(\mem[8][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][26]$_DFFE_PP_  (.D(net21),
    .DE(_0015_),
    .Q(\mem[8][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][27]$_DFFE_PP_  (.D(net22),
    .DE(_0015_),
    .Q(\mem[8][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][28]$_DFFE_PP_  (.D(net23),
    .DE(_0015_),
    .Q(\mem[8][28] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][29]$_DFFE_PP_  (.D(net24),
    .DE(_0015_),
    .Q(\mem[8][29] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net25),
    .DE(_0015_),
    .Q(\mem[8][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][30]$_DFFE_PP_  (.D(net26),
    .DE(_0015_),
    .Q(\mem[8][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][31]$_DFFE_PP_  (.D(net27),
    .DE(_0015_),
    .Q(\mem[8][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net28),
    .DE(_0015_),
    .Q(\mem[8][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net29),
    .DE(_0015_),
    .Q(\mem[8][4] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net30),
    .DE(_0015_),
    .Q(\mem[8][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net31),
    .DE(_0015_),
    .Q(\mem[8][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net32),
    .DE(_0015_),
    .Q(\mem[8][7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][8]$_DFFE_PP_  (.D(net33),
    .DE(_0015_),
    .Q(\mem[8][8] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][9]$_DFFE_PP_  (.D(net34),
    .DE(_0015_),
    .Q(\mem[8][9] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net3),
    .DE(_0016_),
    .Q(\mem[9][0] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][10]$_DFFE_PP_  (.D(net4),
    .DE(_0016_),
    .Q(\mem[9][10] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][11]$_DFFE_PP_  (.D(net5),
    .DE(_0016_),
    .Q(\mem[9][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][12]$_DFFE_PP_  (.D(net6),
    .DE(_0016_),
    .Q(\mem[9][12] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][13]$_DFFE_PP_  (.D(net7),
    .DE(_0016_),
    .Q(\mem[9][13] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][14]$_DFFE_PP_  (.D(net8),
    .DE(_0016_),
    .Q(\mem[9][14] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][15]$_DFFE_PP_  (.D(net9),
    .DE(_0016_),
    .Q(\mem[9][15] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][16]$_DFFE_PP_  (.D(net10),
    .DE(_0016_),
    .Q(\mem[9][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][17]$_DFFE_PP_  (.D(net11),
    .DE(_0016_),
    .Q(\mem[9][17] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][18]$_DFFE_PP_  (.D(net12),
    .DE(_0016_),
    .Q(\mem[9][18] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][19]$_DFFE_PP_  (.D(net13),
    .DE(_0016_),
    .Q(\mem[9][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net14),
    .DE(_0016_),
    .Q(\mem[9][1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][20]$_DFFE_PP_  (.D(net15),
    .DE(_0016_),
    .Q(\mem[9][20] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][21]$_DFFE_PP_  (.D(net16),
    .DE(_0016_),
    .Q(\mem[9][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][22]$_DFFE_PP_  (.D(net17),
    .DE(_0016_),
    .Q(\mem[9][22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][23]$_DFFE_PP_  (.D(net18),
    .DE(_0016_),
    .Q(\mem[9][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][24]$_DFFE_PP_  (.D(net19),
    .DE(_0016_),
    .Q(\mem[9][24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][25]$_DFFE_PP_  (.D(net20),
    .DE(_0016_),
    .Q(\mem[9][25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][26]$_DFFE_PP_  (.D(net21),
    .DE(_0016_),
    .Q(\mem[9][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][27]$_DFFE_PP_  (.D(net22),
    .DE(_0016_),
    .Q(\mem[9][27] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][28]$_DFFE_PP_  (.D(net23),
    .DE(_0016_),
    .Q(\mem[9][28] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][29]$_DFFE_PP_  (.D(net24),
    .DE(_0016_),
    .Q(\mem[9][29] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net25),
    .DE(_0016_),
    .Q(\mem[9][2] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][30]$_DFFE_PP_  (.D(net26),
    .DE(_0016_),
    .Q(\mem[9][30] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][31]$_DFFE_PP_  (.D(net27),
    .DE(_0016_),
    .Q(\mem[9][31] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net28),
    .DE(_0016_),
    .Q(\mem[9][3] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net29),
    .DE(_0016_),
    .Q(\mem[9][4] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net30),
    .DE(_0016_),
    .Q(\mem[9][5] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net31),
    .DE(_0016_),
    .Q(\mem[9][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net32),
    .DE(_0016_),
    .Q(\mem[9][7] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][8]$_DFFE_PP_  (.D(net33),
    .DE(_0016_),
    .Q(\mem[9][8] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][9]$_DFFE_PP_  (.D(net34),
    .DE(_0016_),
    .Q(\mem[9][9] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr[0]$_DFFE_PN0P_  (.D(_0070_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_0071_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_0072_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr[3]$_DFFE_PN0P_  (.D(_0073_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_0074_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_0075_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_0076_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0P_  (.D(_0077_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr[3]$_DFFE_PN0P_  (.D(_0078_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_0079_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net98),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_524 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(net99),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input2 (.A(net105),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(net122),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input4 (.A(net129),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(net118),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(net115),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(net119),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(net123),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input9 (.A(net102),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(net124),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(net125),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(net127),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(net112),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(net114),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(net109),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(net108),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(net117),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input18 (.A(net101),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input19 (.A(net100),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input20 (.A(net103),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(net106),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(net113),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input23 (.A(net104),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(net132),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(net120),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(net116),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(net126),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(net131),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input29 (.A(net110),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(net128),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(net130),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input32 (.A(net107),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input33 (.A(net111),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(net121),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net36),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net37),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net38),
    .X(data_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net39),
    .X(data_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net40),
    .X(data_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net41),
    .X(data_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net42),
    .X(data_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net43),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net44),
    .X(error_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net45),
    .X(error_count[10]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net46),
    .X(error_count[11]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net47),
    .X(error_count[12]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net48),
    .X(error_count[13]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net49),
    .X(error_count[14]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net50),
    .X(error_count[15]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net51),
    .X(error_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net52),
    .X(error_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net53),
    .X(error_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net54),
    .X(error_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net55),
    .X(error_count[5]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net56),
    .X(error_count[6]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net57),
    .X(error_count[7]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net58),
    .X(error_count[8]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net59),
    .X(error_count[9]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net60),
    .X(error_detected));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net61),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net62),
    .X(overflow_detected));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net63),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net64),
    .X(rd_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net65),
    .X(rd_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net66),
    .X(rd_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net67),
    .X(rd_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(rd_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(rd_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(rd_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(rd_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(rd_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(rd_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(rd_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(rd_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(rd_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(rd_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(rd_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(rd_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(rd_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(rd_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(rd_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(rd_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(rd_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(rd_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(rd_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(rd_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(rd_valid));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(underflow_detected));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(wr_ready));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload4 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__bufinv_16 clkload5 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload8 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload10 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload11 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload13 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload16 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload17 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__bufinv_16 clkload19 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload20 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload21 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload22 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_1 clkload23 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__bufinv_16 clkload25 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload27 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_2 clkload28 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_2 clkload29 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinv_1 clkload30 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_1 clkload31 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_2 clkload33 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__bufinv_16 clkload34 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__bufinv_16 clkload35 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload36 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload37 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkinv_1 clkload38 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_1 clkload39 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_2 clkload41 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__bufinv_16 clkload42 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__bufinv_16 clkload43 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinv_1 clkload44 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload45 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload46 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_2 clkload48 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(clear_errors),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(wr_data[25]),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(wr_data[24]),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(wr_data[16]),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(wr_data[26]),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(wr_data[29]),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(wr_data[0]),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(wr_data[27]),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(wr_data[8]),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(wr_data[22]),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(wr_data[21]),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(wr_data[5]),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(wr_data[9]),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(wr_data[1]),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(wr_data[28]),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(wr_data[20]),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(wr_data[13]),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(wr_data[31]),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(wr_data[23]),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(wr_data[12]),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(wr_data[14]),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(wr_data[30]),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(wr_en),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(wr_data[10]),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(wr_data[15]),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(wr_data[17]),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(wr_data[18]),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(wr_data[3]),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(wr_data[19]),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(wr_data[6]),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(wr_data[11]),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(wr_data[7]),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(wr_data[4]),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(wr_data[2]),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(rd_en),
    .X(net133));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_429 ();
endmodule
