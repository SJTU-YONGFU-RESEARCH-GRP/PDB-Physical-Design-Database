module showahead_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    peek_en,
    rd_en,
    rst_n,
    valid,
    wr_en,
    data_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input peek_en;
 input rd_en;
 input rst_n;
 output valid;
 input wr_en;
 output [4:0] data_count;
 output [7:0] rd_data;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net30;
 wire net31;

 sky130_fd_sc_hd__inv_1 _131_ (.A(_130_),
    .Y(net14));
 sky130_fd_sc_hd__inv_1 _132_ (.A(_114_),
    .Y(_029_));
 sky130_fd_sc_hd__nand2_1 _133_ (.A(_119_),
    .B(_116_),
    .Y(_030_));
 sky130_fd_sc_hd__a21oi_1 _134_ (.A1(_119_),
    .A2(_115_),
    .B1(_118_),
    .Y(_031_));
 sky130_fd_sc_hd__o21ai_2 _135_ (.A1(_129_),
    .A2(_030_),
    .B1(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _136_ (.A(_029_),
    .B(_032_),
    .Y(net17));
 sky130_fd_sc_hd__xor2_2 _137_ (.A(_119_),
    .B(_111_),
    .X(net16));
 sky130_fd_sc_hd__a21o_1 _138_ (.A1(_119_),
    .A2(_111_),
    .B1(_118_),
    .X(_033_));
 sky130_fd_sc_hd__a21oi_1 _139_ (.A1(_114_),
    .A2(_033_),
    .B1(_113_),
    .Y(_034_));
 sky130_fd_sc_hd__xnor2_1 _140_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Y(_035_));
 sky130_fd_sc_hd__xor2_2 _141_ (.A(_034_),
    .B(_035_),
    .X(_036_));
 sky130_fd_sc_hd__inv_2 _142_ (.A(_036_),
    .Y(net18));
 sky130_fd_sc_hd__nor4_1 _143_ (.A(_114_),
    .B(net14),
    .C(net15),
    .D(net16),
    .Y(_037_));
 sky130_fd_sc_hd__nor4_1 _144_ (.A(_029_),
    .B(net14),
    .C(net15),
    .D(net16),
    .Y(_038_));
 sky130_fd_sc_hd__mux2_4 _145_ (.A0(_037_),
    .A1(_038_),
    .S(_032_),
    .X(_039_));
 sky130_fd_sc_hd__and2_0 _146_ (.A(net18),
    .B(_039_),
    .X(net20));
 sky130_fd_sc_hd__and2_0 _147_ (.A(_036_),
    .B(_039_),
    .X(_040_));
 sky130_fd_sc_hd__buf_4 _148_ (.A(_040_),
    .X(net19));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .Y(_041_));
 sky130_fd_sc_hd__a21boi_2 _150_ (.A1(net18),
    .A2(_039_),
    .B1_N(net11),
    .Y(_042_));
 sky130_fd_sc_hd__and3_4 _151_ (.A(_122_),
    .B(_041_),
    .C(_042_),
    .X(_000_));
 sky130_fd_sc_hd__and3_4 _152_ (.A(_125_),
    .B(_041_),
    .C(_042_),
    .X(_007_));
 sky130_fd_sc_hd__and3_4 _153_ (.A(_123_),
    .B(_041_),
    .C(_042_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _154_ (.A(net11),
    .B(_127_),
    .Y(_043_));
 sky130_fd_sc_hd__a21oi_2 _155_ (.A1(net18),
    .A2(_039_),
    .B1(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__and2_4 _156_ (.A(_041_),
    .B(_044_),
    .X(_009_));
 sky130_fd_sc_hd__buf_4 _157_ (.A(_042_),
    .X(_045_));
 sky130_fd_sc_hd__nor2b_1 _158_ (.A(\wr_ptr[3] ),
    .B_N(\wr_ptr[2] ),
    .Y(_046_));
 sky130_fd_sc_hd__and3_4 _159_ (.A(_122_),
    .B(_045_),
    .C(_046_),
    .X(_010_));
 sky130_fd_sc_hd__and3_4 _160_ (.A(_125_),
    .B(_045_),
    .C(_046_),
    .X(_011_));
 sky130_fd_sc_hd__and3_4 _161_ (.A(_123_),
    .B(_045_),
    .C(_046_),
    .X(_012_));
 sky130_fd_sc_hd__and2_4 _162_ (.A(_044_),
    .B(_046_),
    .X(_013_));
 sky130_fd_sc_hd__nor2b_2 _163_ (.A(\wr_ptr[2] ),
    .B_N(\wr_ptr[3] ),
    .Y(_047_));
 sky130_fd_sc_hd__and3_4 _164_ (.A(_122_),
    .B(_045_),
    .C(_047_),
    .X(_014_));
 sky130_fd_sc_hd__and3_4 _165_ (.A(_125_),
    .B(_045_),
    .C(_047_),
    .X(_015_));
 sky130_fd_sc_hd__and3_4 _166_ (.A(_123_),
    .B(_045_),
    .C(_047_),
    .X(_001_));
 sky130_fd_sc_hd__and2_4 _167_ (.A(_044_),
    .B(_047_),
    .X(_002_));
 sky130_fd_sc_hd__and2_1 _168_ (.A(\wr_ptr[3] ),
    .B(\wr_ptr[2] ),
    .X(_048_));
 sky130_fd_sc_hd__and3_4 _169_ (.A(_122_),
    .B(_045_),
    .C(_048_),
    .X(_003_));
 sky130_fd_sc_hd__and3_4 _170_ (.A(_125_),
    .B(_045_),
    .C(_048_),
    .X(_004_));
 sky130_fd_sc_hd__and3_2 _171_ (.A(_123_),
    .B(_045_),
    .C(_048_),
    .X(_005_));
 sky130_fd_sc_hd__nand3_1 _172_ (.A(net11),
    .B(_127_),
    .C(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__a21oi_4 _173_ (.A1(net18),
    .A2(_039_),
    .B1(_049_),
    .Y(_006_));
 sky130_fd_sc_hd__inv_6 _174_ (.A(\rd_ptr[3] ),
    .Y(_112_));
 sky130_fd_sc_hd__buf_6 _175_ (.A(\rd_ptr[1] ),
    .X(_050_));
 sky130_fd_sc_hd__inv_1 _176_ (.A(_050_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_1 _177_ (.A(_129_),
    .Y(_110_));
 sky130_fd_sc_hd__buf_6 _178_ (.A(\rd_ptr[2] ),
    .X(_051_));
 sky130_fd_sc_hd__buf_6 _179_ (.A(_051_),
    .X(_052_));
 sky130_fd_sc_hd__inv_1 _180_ (.A(_052_),
    .Y(_117_));
 sky130_fd_sc_hd__inv_1 _181_ (.A(\wr_ptr[0] ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_1 _182_ (.A(\wr_ptr[1] ),
    .Y(_121_));
 sky130_fd_sc_hd__buf_6 _183_ (.A(\rd_ptr[0] ),
    .X(_053_));
 sky130_fd_sc_hd__buf_8 _184_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__a21boi_1 _185_ (.A1(_036_),
    .A2(_039_),
    .B1_N(net2),
    .Y(_055_));
 sky130_fd_sc_hd__xor2_1 _186_ (.A(_054_),
    .B(_055_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _187_ (.A0(_050_),
    .A1(_018_),
    .S(_055_),
    .X(_020_));
 sky130_fd_sc_hd__nand2_1 _188_ (.A(net2),
    .B(_120_),
    .Y(_056_));
 sky130_fd_sc_hd__a21oi_1 _189_ (.A1(_036_),
    .A2(_039_),
    .B1(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__xnor2_1 _190_ (.A(_117_),
    .B(_057_),
    .Y(_021_));
 sky130_fd_sc_hd__nand4_1 _191_ (.A(net2),
    .B(_054_),
    .C(_050_),
    .D(_052_),
    .Y(_058_));
 sky130_fd_sc_hd__a21oi_1 _192_ (.A1(_036_),
    .A2(_039_),
    .B1(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__xnor2_1 _193_ (.A(_112_),
    .B(_059_),
    .Y(_022_));
 sky130_fd_sc_hd__nand4_1 _194_ (.A(net2),
    .B(_052_),
    .C(\rd_ptr[3] ),
    .D(_120_),
    .Y(_060_));
 sky130_fd_sc_hd__a21oi_1 _195_ (.A1(_036_),
    .A2(_039_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__xor2_1 _196_ (.A(\rd_ptr[4] ),
    .B(_061_),
    .X(_023_));
 sky130_fd_sc_hd__xnor2_1 _197_ (.A(_016_),
    .B(_045_),
    .Y(_024_));
 sky130_fd_sc_hd__mux2_1 _198_ (.A0(\wr_ptr[1] ),
    .A1(_017_),
    .S(_042_),
    .X(_025_));
 sky130_fd_sc_hd__xor2_1 _199_ (.A(\wr_ptr[2] ),
    .B(_044_),
    .X(_026_));
 sky130_fd_sc_hd__nand4_1 _200_ (.A(net11),
    .B(\wr_ptr[2] ),
    .C(\wr_ptr[1] ),
    .D(\wr_ptr[0] ),
    .Y(_062_));
 sky130_fd_sc_hd__a21oi_1 _201_ (.A1(net18),
    .A2(_039_),
    .B1(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__xor2_1 _202_ (.A(\wr_ptr[3] ),
    .B(_063_),
    .X(_027_));
 sky130_fd_sc_hd__xor2_1 _203_ (.A(\wr_ptr[4] ),
    .B(_006_),
    .X(_028_));
 sky130_fd_sc_hd__inv_1 _204_ (.A(net19),
    .Y(net29));
 sky130_fd_sc_hd__xor2_1 _205_ (.A(_130_),
    .B(net15),
    .X(_064_));
 sky130_fd_sc_hd__nor4_1 _206_ (.A(net17),
    .B(net16),
    .C(net18),
    .D(_064_),
    .Y(net12));
 sky130_fd_sc_hd__a31o_1 _207_ (.A1(net15),
    .A2(net17),
    .A3(net16),
    .B1(net18),
    .X(net13));
 sky130_fd_sc_hd__buf_8 _208_ (.A(_053_),
    .X(_065_));
 sky130_fd_sc_hd__buf_4 _209_ (.A(_051_),
    .X(_066_));
 sky130_fd_sc_hd__mux4_1 _210_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[12][0] ),
    .A3(\mem[13][0] ),
    .S0(_065_),
    .S1(_066_),
    .X(_067_));
 sky130_fd_sc_hd__buf_16 _211_ (.A(_053_),
    .X(_068_));
 sky130_fd_sc_hd__buf_4 _212_ (.A(_051_),
    .X(_069_));
 sky130_fd_sc_hd__mux4_1 _213_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[4][0] ),
    .A3(\mem[5][0] ),
    .S0(_068_),
    .S1(_069_),
    .X(_070_));
 sky130_fd_sc_hd__mux4_1 _214_ (.A0(\mem[10][0] ),
    .A1(\mem[11][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(_065_),
    .S1(_066_),
    .X(_071_));
 sky130_fd_sc_hd__mux4_1 _215_ (.A0(\mem[2][0] ),
    .A1(\mem[3][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(_054_),
    .S1(_052_),
    .X(_072_));
 sky130_fd_sc_hd__mux4_1 _216_ (.A0(_067_),
    .A1(_070_),
    .A2(_071_),
    .A3(_072_),
    .S0(_112_),
    .S1(_050_),
    .X(_073_));
 sky130_fd_sc_hd__nor2b_1 _217_ (.A(net19),
    .B_N(_073_),
    .Y(net21));
 sky130_fd_sc_hd__mux4_1 _218_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[12][1] ),
    .A3(\mem[13][1] ),
    .S0(_065_),
    .S1(_066_),
    .X(_074_));
 sky130_fd_sc_hd__mux4_1 _219_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[4][1] ),
    .A3(\mem[5][1] ),
    .S0(_068_),
    .S1(_069_),
    .X(_075_));
 sky130_fd_sc_hd__mux4_1 _220_ (.A0(\mem[10][1] ),
    .A1(\mem[11][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(_065_),
    .S1(_069_),
    .X(_076_));
 sky130_fd_sc_hd__mux4_2 _221_ (.A0(\mem[2][1] ),
    .A1(\mem[3][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(_054_),
    .S1(_052_),
    .X(_077_));
 sky130_fd_sc_hd__mux4_1 _222_ (.A0(_074_),
    .A1(_075_),
    .A2(_076_),
    .A3(_077_),
    .S0(_112_),
    .S1(_050_),
    .X(_078_));
 sky130_fd_sc_hd__nor2b_1 _223_ (.A(net19),
    .B_N(_078_),
    .Y(net22));
 sky130_fd_sc_hd__mux4_1 _224_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[12][2] ),
    .A3(\mem[13][2] ),
    .S0(_065_),
    .S1(_066_),
    .X(_079_));
 sky130_fd_sc_hd__mux4_1 _225_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[4][2] ),
    .A3(\mem[5][2] ),
    .S0(_068_),
    .S1(_069_),
    .X(_080_));
 sky130_fd_sc_hd__mux4_1 _226_ (.A0(\mem[10][2] ),
    .A1(\mem[11][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(_068_),
    .S1(_069_),
    .X(_081_));
 sky130_fd_sc_hd__mux4_1 _227_ (.A0(\mem[2][2] ),
    .A1(\mem[3][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(_054_),
    .S1(_052_),
    .X(_082_));
 sky130_fd_sc_hd__mux4_1 _228_ (.A0(_079_),
    .A1(_080_),
    .A2(_081_),
    .A3(_082_),
    .S0(_112_),
    .S1(_050_),
    .X(_083_));
 sky130_fd_sc_hd__nor2b_1 _229_ (.A(net19),
    .B_N(_083_),
    .Y(net23));
 sky130_fd_sc_hd__mux4_1 _230_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[12][3] ),
    .A3(\mem[13][3] ),
    .S0(_065_),
    .S1(_066_),
    .X(_084_));
 sky130_fd_sc_hd__mux4_1 _231_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[4][3] ),
    .A3(\mem[5][3] ),
    .S0(_068_),
    .S1(_051_),
    .X(_085_));
 sky130_fd_sc_hd__mux4_1 _232_ (.A0(\mem[10][3] ),
    .A1(\mem[11][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(_068_),
    .S1(_069_),
    .X(_086_));
 sky130_fd_sc_hd__mux4_2 _233_ (.A0(\mem[2][3] ),
    .A1(\mem[3][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(_054_),
    .S1(_052_),
    .X(_087_));
 sky130_fd_sc_hd__mux4_1 _234_ (.A0(_084_),
    .A1(_085_),
    .A2(_086_),
    .A3(_087_),
    .S0(_112_),
    .S1(_050_),
    .X(_088_));
 sky130_fd_sc_hd__nor2b_1 _235_ (.A(net19),
    .B_N(_088_),
    .Y(net24));
 sky130_fd_sc_hd__mux4_1 _236_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[12][4] ),
    .A3(\mem[13][4] ),
    .S0(_065_),
    .S1(_066_),
    .X(_089_));
 sky130_fd_sc_hd__mux4_1 _237_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[4][4] ),
    .A3(\mem[5][4] ),
    .S0(_053_),
    .S1(_051_),
    .X(_090_));
 sky130_fd_sc_hd__mux4_1 _238_ (.A0(\mem[10][4] ),
    .A1(\mem[11][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(_068_),
    .S1(_069_),
    .X(_091_));
 sky130_fd_sc_hd__mux4_4 _239_ (.A0(\mem[2][4] ),
    .A1(\mem[3][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(_054_),
    .S1(_052_),
    .X(_092_));
 sky130_fd_sc_hd__mux4_1 _240_ (.A0(_089_),
    .A1(_090_),
    .A2(_091_),
    .A3(_092_),
    .S0(_112_),
    .S1(_050_),
    .X(_093_));
 sky130_fd_sc_hd__nor2b_1 _241_ (.A(net19),
    .B_N(_093_),
    .Y(net25));
 sky130_fd_sc_hd__mux4_1 _242_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[12][5] ),
    .A3(\mem[13][5] ),
    .S0(_065_),
    .S1(_066_),
    .X(_094_));
 sky130_fd_sc_hd__mux4_1 _243_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[4][5] ),
    .A3(\mem[5][5] ),
    .S0(_053_),
    .S1(_051_),
    .X(_095_));
 sky130_fd_sc_hd__mux4_2 _244_ (.A0(\mem[10][5] ),
    .A1(\mem[11][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(_068_),
    .S1(_069_),
    .X(_096_));
 sky130_fd_sc_hd__mux4_2 _245_ (.A0(\mem[2][5] ),
    .A1(\mem[3][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(_054_),
    .S1(_052_),
    .X(_097_));
 sky130_fd_sc_hd__mux4_1 _246_ (.A0(_094_),
    .A1(_095_),
    .A2(_096_),
    .A3(_097_),
    .S0(_112_),
    .S1(_050_),
    .X(_098_));
 sky130_fd_sc_hd__nor2b_1 _247_ (.A(net19),
    .B_N(_098_),
    .Y(net26));
 sky130_fd_sc_hd__mux4_1 _248_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[12][6] ),
    .A3(\mem[13][6] ),
    .S0(_065_),
    .S1(_066_),
    .X(_099_));
 sky130_fd_sc_hd__mux4_1 _249_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[4][6] ),
    .A3(\mem[5][6] ),
    .S0(_053_),
    .S1(_051_),
    .X(_100_));
 sky130_fd_sc_hd__mux4_4 _250_ (.A0(\mem[10][6] ),
    .A1(\mem[11][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(_068_),
    .S1(_069_),
    .X(_101_));
 sky130_fd_sc_hd__mux4_2 _251_ (.A0(\mem[2][6] ),
    .A1(\mem[3][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(_054_),
    .S1(_052_),
    .X(_102_));
 sky130_fd_sc_hd__mux4_1 _252_ (.A0(_099_),
    .A1(_100_),
    .A2(_101_),
    .A3(_102_),
    .S0(_112_),
    .S1(_050_),
    .X(_103_));
 sky130_fd_sc_hd__nor2b_1 _253_ (.A(net19),
    .B_N(_103_),
    .Y(net27));
 sky130_fd_sc_hd__mux4_1 _254_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[12][7] ),
    .A3(\mem[13][7] ),
    .S0(_065_),
    .S1(_066_),
    .X(_104_));
 sky130_fd_sc_hd__mux4_1 _255_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[4][7] ),
    .A3(\mem[5][7] ),
    .S0(_053_),
    .S1(_051_),
    .X(_105_));
 sky130_fd_sc_hd__mux4_2 _256_ (.A0(\mem[10][7] ),
    .A1(\mem[11][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(_068_),
    .S1(_069_),
    .X(_106_));
 sky130_fd_sc_hd__mux4_1 _257_ (.A0(\mem[2][7] ),
    .A1(\mem[3][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(_054_),
    .S1(_066_),
    .X(_107_));
 sky130_fd_sc_hd__mux4_1 _258_ (.A0(_104_),
    .A1(_105_),
    .A2(_106_),
    .A3(_107_),
    .S0(_112_),
    .S1(\rd_ptr[1] ),
    .X(_108_));
 sky130_fd_sc_hd__nor2b_1 _259_ (.A(net19),
    .B_N(_108_),
    .Y(net28));
 sky130_fd_sc_hd__fa_2 _260_ (.A(_109_),
    .B(\wr_ptr[1] ),
    .CIN(_110_),
    .COUT(_111_),
    .SUM(net15));
 sky130_fd_sc_hd__ha_1 _261_ (.A(_112_),
    .B(\wr_ptr[3] ),
    .COUT(_113_),
    .SUM(_114_));
 sky130_fd_sc_hd__ha_1 _262_ (.A(_109_),
    .B(\wr_ptr[1] ),
    .COUT(_115_),
    .SUM(_116_));
 sky130_fd_sc_hd__ha_1 _263_ (.A(_117_),
    .B(\wr_ptr[2] ),
    .COUT(_118_),
    .SUM(_119_));
 sky130_fd_sc_hd__ha_1 _264_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_120_),
    .SUM(_018_));
 sky130_fd_sc_hd__ha_1 _265_ (.A(_016_),
    .B(_121_),
    .COUT(_122_),
    .SUM(_017_));
 sky130_fd_sc_hd__ha_1 _266_ (.A(_016_),
    .B(\wr_ptr[1] ),
    .COUT(_123_),
    .SUM(_124_));
 sky130_fd_sc_hd__ha_1 _267_ (.A(\wr_ptr[0] ),
    .B(_121_),
    .COUT(_125_),
    .SUM(_126_));
 sky130_fd_sc_hd__ha_1 _268_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_127_),
    .SUM(_128_));
 sky130_fd_sc_hd__ha_1 _269_ (.A(\rd_ptr[0] ),
    .B(_016_),
    .COUT(_129_),
    .SUM(_130_));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net3),
    .DE(_000_),
    .Q(\mem[0][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net4),
    .DE(_000_),
    .Q(\mem[0][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net5),
    .DE(_000_),
    .Q(\mem[0][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net6),
    .DE(_000_),
    .Q(\mem[0][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net7),
    .DE(_000_),
    .Q(\mem[0][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\mem[0][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\mem[0][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net10),
    .DE(_000_),
    .Q(\mem[0][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net3),
    .DE(_001_),
    .Q(\mem[10][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\mem[10][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\mem[10][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\mem[10][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\mem[10][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\mem[10][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\mem[10][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net10),
    .DE(_001_),
    .Q(\mem[10][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net3),
    .DE(_002_),
    .Q(\mem[11][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\mem[11][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\mem[11][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\mem[11][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\mem[11][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\mem[11][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\mem[11][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net10),
    .DE(_002_),
    .Q(\mem[11][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net3),
    .DE(_003_),
    .Q(\mem[12][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\mem[12][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\mem[12][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\mem[12][3] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\mem[12][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\mem[12][5] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\mem[12][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net10),
    .DE(_003_),
    .Q(\mem[12][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net3),
    .DE(_004_),
    .Q(\mem[13][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\mem[13][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\mem[13][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\mem[13][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\mem[13][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\mem[13][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\mem[13][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net10),
    .DE(_004_),
    .Q(\mem[13][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net3),
    .DE(_005_),
    .Q(\mem[14][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\mem[14][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\mem[14][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\mem[14][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\mem[14][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\mem[14][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\mem[14][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net10),
    .DE(_005_),
    .Q(\mem[14][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net3),
    .DE(_006_),
    .Q(\mem[15][0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\mem[15][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\mem[15][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\mem[15][3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\mem[15][4] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\mem[15][5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\mem[15][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net10),
    .DE(_006_),
    .Q(\mem[15][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net3),
    .DE(_007_),
    .Q(\mem[1][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\mem[1][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\mem[1][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\mem[1][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\mem[1][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\mem[1][5] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\mem[1][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net10),
    .DE(_007_),
    .Q(\mem[1][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net3),
    .DE(_008_),
    .Q(\mem[2][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\mem[2][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\mem[2][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\mem[2][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\mem[2][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\mem[2][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\mem[2][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net10),
    .DE(_008_),
    .Q(\mem[2][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net3),
    .DE(_009_),
    .Q(\mem[3][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\mem[3][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\mem[3][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\mem[3][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\mem[3][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\mem[3][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\mem[3][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net10),
    .DE(_009_),
    .Q(\mem[3][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net3),
    .DE(_010_),
    .Q(\mem[4][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\mem[4][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\mem[4][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\mem[4][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\mem[4][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\mem[4][5] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\mem[4][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net10),
    .DE(_010_),
    .Q(\mem[4][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net3),
    .DE(_011_),
    .Q(\mem[5][0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\mem[5][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[5][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[5][3] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[5][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[5][5] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[5][6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[5][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net3),
    .DE(_012_),
    .Q(\mem[6][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\mem[6][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[6][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[6][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[6][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[6][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[6][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[6][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net3),
    .DE(_013_),
    .Q(\mem[7][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\mem[7][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[7][2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[7][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[7][4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[7][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[7][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[7][7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net3),
    .DE(_014_),
    .Q(\mem[8][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\mem[8][1] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[8][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[8][3] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[8][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[8][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[8][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[8][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net3),
    .DE(_015_),
    .Q(\mem[9][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\mem[9][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[9][2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[9][3] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[9][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[9][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[9][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[9][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_019_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_020_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[2]$_DFFE_PN0P_  (.D(_021_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_022_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_023_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_024_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[1]$_DFFE_PN0P_  (.D(_025_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[2]$_DFFE_PN0P_  (.D(_026_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \wr_ptr[3]$_DFFE_PN0P_  (.D(_027_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_028_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_4 hold1 (.A(net30),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_135 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input2 (.A(wr_data[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input3 (.A(wr_data[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(wr_data[2]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(net31),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[5]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(wr_data[6]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input9 (.A(wr_data[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(wr_en),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(data_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(data_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(data_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(data_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(data_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(wr_data[4]),
    .X(net31));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_216 ();
endmodule
