module clock_domain_crossing_fifo (rd_almost_empty,
    rd_clk,
    rd_empty,
    rd_en,
    rd_rst_n,
    wr_almost_full,
    wr_clk,
    wr_en,
    wr_full,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output rd_almost_empty;
 input rd_clk;
 output rd_empty;
 input rd_en;
 input rd_rst_n;
 output wr_almost_full;
 input wr_clk;
 input wr_en;
 output wr_full;
 input wr_rst_n;
 output [4:0] rd_count;
 output [31:0] rd_data;
 output [4:0] wr_count;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire clknet_leaf_0_wr_clk;
 wire clknet_leaf_1_wr_clk;
 wire clknet_leaf_2_wr_clk;
 wire clknet_leaf_3_wr_clk;
 wire clknet_leaf_4_wr_clk;
 wire clknet_leaf_5_wr_clk;
 wire clknet_leaf_6_wr_clk;
 wire clknet_leaf_7_wr_clk;
 wire clknet_leaf_8_wr_clk;
 wire clknet_leaf_9_wr_clk;
 wire clknet_leaf_10_wr_clk;
 wire clknet_leaf_11_wr_clk;
 wire clknet_leaf_12_wr_clk;
 wire clknet_leaf_13_wr_clk;
 wire clknet_leaf_14_wr_clk;
 wire clknet_leaf_15_wr_clk;
 wire clknet_leaf_16_wr_clk;
 wire clknet_leaf_17_wr_clk;
 wire clknet_leaf_18_wr_clk;
 wire clknet_leaf_19_wr_clk;
 wire clknet_leaf_20_wr_clk;
 wire clknet_leaf_21_wr_clk;
 wire clknet_leaf_22_wr_clk;
 wire clknet_leaf_23_wr_clk;
 wire clknet_leaf_24_wr_clk;
 wire clknet_leaf_25_wr_clk;
 wire clknet_leaf_26_wr_clk;
 wire clknet_leaf_27_wr_clk;
 wire clknet_leaf_28_wr_clk;
 wire clknet_leaf_29_wr_clk;
 wire clknet_leaf_30_wr_clk;
 wire clknet_leaf_31_wr_clk;
 wire clknet_leaf_32_wr_clk;
 wire clknet_leaf_33_wr_clk;
 wire clknet_leaf_34_wr_clk;
 wire clknet_leaf_35_wr_clk;
 wire clknet_leaf_36_wr_clk;
 wire clknet_leaf_37_wr_clk;
 wire clknet_leaf_38_wr_clk;
 wire clknet_leaf_39_wr_clk;
 wire clknet_leaf_40_wr_clk;
 wire clknet_leaf_41_wr_clk;
 wire clknet_leaf_42_wr_clk;
 wire clknet_leaf_43_wr_clk;
 wire clknet_leaf_44_wr_clk;
 wire clknet_leaf_45_wr_clk;
 wire clknet_leaf_46_wr_clk;
 wire clknet_leaf_47_wr_clk;
 wire clknet_leaf_48_wr_clk;
 wire clknet_leaf_49_wr_clk;
 wire clknet_leaf_50_wr_clk;
 wire clknet_leaf_51_wr_clk;
 wire clknet_leaf_52_wr_clk;
 wire clknet_leaf_53_wr_clk;
 wire clknet_leaf_54_wr_clk;
 wire clknet_leaf_55_wr_clk;
 wire clknet_leaf_56_wr_clk;
 wire clknet_leaf_57_wr_clk;
 wire clknet_leaf_58_wr_clk;
 wire clknet_leaf_59_wr_clk;
 wire clknet_leaf_60_wr_clk;
 wire clknet_leaf_61_wr_clk;
 wire clknet_leaf_62_wr_clk;
 wire clknet_leaf_63_wr_clk;
 wire clknet_leaf_64_wr_clk;
 wire clknet_leaf_65_wr_clk;
 wire clknet_leaf_66_wr_clk;
 wire clknet_leaf_67_wr_clk;
 wire clknet_leaf_68_wr_clk;
 wire clknet_leaf_69_wr_clk;
 wire clknet_leaf_70_wr_clk;
 wire clknet_leaf_71_wr_clk;
 wire clknet_leaf_72_wr_clk;
 wire clknet_leaf_73_wr_clk;
 wire clknet_0_wr_clk;
 wire clknet_3_0__leaf_wr_clk;
 wire clknet_3_1__leaf_wr_clk;
 wire clknet_3_2__leaf_wr_clk;
 wire clknet_3_3__leaf_wr_clk;
 wire clknet_3_4__leaf_wr_clk;
 wire clknet_3_5__leaf_wr_clk;
 wire clknet_3_6__leaf_wr_clk;
 wire clknet_3_7__leaf_wr_clk;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;

 XNOR2_X2 _2012_ (.A(\rd_ptr_gray_sync2[3] ),
    .B(\rd_ptr_gray_sync2[4] ),
    .ZN(_1979_));
 XNOR2_X2 _2013_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_1979_),
    .ZN(_0568_));
 XNOR2_X2 _2014_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_0568_),
    .ZN(_1969_));
 INV_X1 _2015_ (.A(_2011_),
    .ZN(net46));
 INV_X1 _2016_ (.A(_0568_),
    .ZN(_1976_));
 BUF_X2 _2017_ (.A(_1978_),
    .Z(_0569_));
 XOR2_X2 _2018_ (.A(\rd_ptr_gray_sync2[4] ),
    .B(\wr_ptr_bin[4] ),
    .Z(_0570_));
 AND2_X1 _2019_ (.A1(_1975_),
    .A2(_2011_),
    .ZN(_0571_));
 NAND4_X4 _2020_ (.A1(_1981_),
    .A2(_0569_),
    .A3(_0570_),
    .A4(_0571_),
    .ZN(_0572_));
 INV_X1 _2021_ (.A(_0572_),
    .ZN(net51));
 INV_X1 _2022_ (.A(_1974_),
    .ZN(_0573_));
 INV_X1 _2023_ (.A(_1975_),
    .ZN(_0574_));
 OAI21_X1 _2024_ (.A(_0573_),
    .B1(_1965_),
    .B2(_0574_),
    .ZN(_0575_));
 AOI21_X1 _2025_ (.A(_1977_),
    .B1(_0569_),
    .B2(_0575_),
    .ZN(_0576_));
 XOR2_X2 _2026_ (.A(_1981_),
    .B(_0576_),
    .Z(_0577_));
 INV_X1 _2027_ (.A(_0577_),
    .ZN(net49));
 INV_X1 _2028_ (.A(_1977_),
    .ZN(_0578_));
 INV_X1 _2029_ (.A(_0569_),
    .ZN(_0579_));
 OAI21_X1 _2030_ (.A(_0578_),
    .B1(_1967_),
    .B2(_0579_),
    .ZN(_0580_));
 AOI21_X1 _2031_ (.A(_1980_),
    .B1(_0580_),
    .B2(_1981_),
    .ZN(_0581_));
 XNOR2_X1 _2032_ (.A(_0570_),
    .B(_0581_),
    .ZN(_0582_));
 INV_X1 _2033_ (.A(_0582_),
    .ZN(net50));
 XOR2_X2 _2034_ (.A(\wr_ptr_gray_sync2[3] ),
    .B(\wr_ptr_gray_sync2[4] ),
    .Z(_1987_));
 XOR2_X2 _2035_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(_1987_),
    .Z(_1991_));
 XNOR2_X2 _2036_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_1991_),
    .ZN(_1971_));
 INV_X1 _2037_ (.A(_1973_),
    .ZN(net8));
 XNOR2_X1 _2038_ (.A(_1972_),
    .B(_1993_),
    .ZN(net9));
 INV_X1 _2039_ (.A(_1992_),
    .ZN(_0583_));
 INV_X1 _2040_ (.A(_1970_),
    .ZN(_0584_));
 AOI21_X1 _2041_ (.A(_1984_),
    .B1(_0584_),
    .B2(_1985_),
    .ZN(_0585_));
 INV_X1 _2042_ (.A(_1993_),
    .ZN(_0586_));
 OAI21_X1 _2043_ (.A(_0583_),
    .B1(_0585_),
    .B2(_0586_),
    .ZN(_0587_));
 XOR2_X1 _2044_ (.A(_1989_),
    .B(_0587_),
    .Z(net10));
 XNOR2_X2 _2045_ (.A(\wr_ptr_gray_sync2[4] ),
    .B(\rd_ptr_bin[4] ),
    .ZN(_0588_));
 OAI21_X1 _2046_ (.A(_0583_),
    .B1(_0586_),
    .B2(_1972_),
    .ZN(_0589_));
 AOI21_X1 _2047_ (.A(_1988_),
    .B1(_0589_),
    .B2(_1989_),
    .ZN(_0590_));
 XNOR2_X1 _2048_ (.A(_0588_),
    .B(_0590_),
    .ZN(net11));
 INV_X1 _2049_ (.A(_0588_),
    .ZN(_0591_));
 XNOR2_X1 _2050_ (.A(\wr_ptr_gray_sync2[3] ),
    .B(\rd_ptr_gray[3] ),
    .ZN(_0592_));
 XNOR2_X1 _2051_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(\rd_ptr_gray[0] ),
    .ZN(_0593_));
 XNOR2_X1 _2052_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(\rd_ptr_gray[1] ),
    .ZN(_0594_));
 XNOR2_X1 _2053_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(\rd_ptr_gray[2] ),
    .ZN(_0595_));
 NAND4_X2 _2054_ (.A1(_0592_),
    .A2(_0593_),
    .A3(_0594_),
    .A4(_0595_),
    .ZN(_0596_));
 NOR2_X1 _2055_ (.A1(_0591_),
    .A2(_0596_),
    .ZN(net44));
 INV_X1 _2056_ (.A(_1969_),
    .ZN(_1966_));
 INV_X1 _2057_ (.A(_1971_),
    .ZN(_1983_));
 XOR2_X2 _2058_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_1971_),
    .Z(_2008_));
 XNOR2_X1 _2059_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_1969_),
    .ZN(_2010_));
 INV_X1 _2060_ (.A(_2009_),
    .ZN(net7));
 CLKBUF_X2 _2061_ (.A(wr_data[0]),
    .Z(_0597_));
 BUF_X2 _2062_ (.A(_0597_),
    .Z(_0598_));
 BUF_X2 _2063_ (.A(\wr_ptr_bin[2] ),
    .Z(_0599_));
 NOR2_X4 _2064_ (.A1(\wr_ptr_bin[3] ),
    .A2(_0599_),
    .ZN(_0600_));
 AND2_X4 _2065_ (.A1(net4),
    .A2(net5),
    .ZN(_0601_));
 AND3_X2 _2066_ (.A1(_1994_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0602_));
 NAND2_X4 _2067_ (.A1(_0600_),
    .A2(_0602_),
    .ZN(_0603_));
 BUF_X4 _2068_ (.A(_0603_),
    .Z(_0604_));
 MUX2_X1 _2069_ (.A(_0598_),
    .B(\mem[0][0] ),
    .S(_0604_),
    .Z(_0006_));
 CLKBUF_X2 _2070_ (.A(wr_data[10]),
    .Z(_0605_));
 BUF_X2 _2071_ (.A(_0605_),
    .Z(_0606_));
 MUX2_X1 _2072_ (.A(_0606_),
    .B(\mem[0][10] ),
    .S(_0604_),
    .Z(_0007_));
 CLKBUF_X2 _2073_ (.A(wr_data[11]),
    .Z(_0607_));
 BUF_X2 _2074_ (.A(_0607_),
    .Z(_0608_));
 MUX2_X1 _2075_ (.A(_0608_),
    .B(\mem[0][11] ),
    .S(_0604_),
    .Z(_0008_));
 BUF_X1 _2076_ (.A(wr_data[12]),
    .Z(_0609_));
 CLKBUF_X2 _2077_ (.A(_0609_),
    .Z(_0610_));
 MUX2_X1 _2078_ (.A(_0610_),
    .B(\mem[0][12] ),
    .S(_0604_),
    .Z(_0009_));
 CLKBUF_X2 _2079_ (.A(wr_data[13]),
    .Z(_0611_));
 BUF_X2 _2080_ (.A(_0611_),
    .Z(_0612_));
 MUX2_X1 _2081_ (.A(_0612_),
    .B(\mem[0][13] ),
    .S(_0604_),
    .Z(_0010_));
 CLKBUF_X2 _2082_ (.A(wr_data[14]),
    .Z(_0613_));
 BUF_X2 _2083_ (.A(_0613_),
    .Z(_0614_));
 MUX2_X1 _2084_ (.A(_0614_),
    .B(\mem[0][14] ),
    .S(_0604_),
    .Z(_0011_));
 CLKBUF_X2 _2085_ (.A(wr_data[15]),
    .Z(_0615_));
 BUF_X2 _2086_ (.A(_0615_),
    .Z(_0616_));
 MUX2_X1 _2087_ (.A(_0616_),
    .B(\mem[0][15] ),
    .S(_0604_),
    .Z(_0012_));
 BUF_X1 _2088_ (.A(wr_data[16]),
    .Z(_0617_));
 BUF_X2 _2089_ (.A(_0617_),
    .Z(_0618_));
 MUX2_X1 _2090_ (.A(_0618_),
    .B(\mem[0][16] ),
    .S(_0604_),
    .Z(_0013_));
 BUF_X1 _2091_ (.A(wr_data[17]),
    .Z(_0619_));
 BUF_X2 _2092_ (.A(_0619_),
    .Z(_0620_));
 MUX2_X1 _2093_ (.A(_0620_),
    .B(\mem[0][17] ),
    .S(_0604_),
    .Z(_0014_));
 CLKBUF_X2 _2094_ (.A(wr_data[18]),
    .Z(_0621_));
 BUF_X2 _2095_ (.A(_0621_),
    .Z(_0622_));
 MUX2_X1 _2096_ (.A(_0622_),
    .B(\mem[0][18] ),
    .S(_0604_),
    .Z(_0015_));
 BUF_X1 _2097_ (.A(wr_data[19]),
    .Z(_0623_));
 BUF_X2 _2098_ (.A(_0623_),
    .Z(_0624_));
 BUF_X4 _2099_ (.A(_0603_),
    .Z(_0625_));
 MUX2_X1 _2100_ (.A(_0624_),
    .B(\mem[0][19] ),
    .S(_0625_),
    .Z(_0016_));
 BUF_X1 _2101_ (.A(wr_data[1]),
    .Z(_0626_));
 CLKBUF_X2 _2102_ (.A(_0626_),
    .Z(_0627_));
 MUX2_X1 _2103_ (.A(_0627_),
    .B(\mem[0][1] ),
    .S(_0625_),
    .Z(_0017_));
 CLKBUF_X2 _2104_ (.A(wr_data[20]),
    .Z(_0628_));
 CLKBUF_X2 _2105_ (.A(_0628_),
    .Z(_0629_));
 MUX2_X1 _2106_ (.A(_0629_),
    .B(\mem[0][20] ),
    .S(_0625_),
    .Z(_0018_));
 BUF_X1 _2107_ (.A(wr_data[21]),
    .Z(_0630_));
 BUF_X2 _2108_ (.A(_0630_),
    .Z(_0631_));
 MUX2_X1 _2109_ (.A(_0631_),
    .B(\mem[0][21] ),
    .S(_0625_),
    .Z(_0019_));
 CLKBUF_X2 _2110_ (.A(wr_data[22]),
    .Z(_0632_));
 BUF_X2 _2111_ (.A(_0632_),
    .Z(_0633_));
 MUX2_X1 _2112_ (.A(_0633_),
    .B(\mem[0][22] ),
    .S(_0625_),
    .Z(_0020_));
 CLKBUF_X2 _2113_ (.A(wr_data[23]),
    .Z(_0634_));
 BUF_X2 _2114_ (.A(_0634_),
    .Z(_0635_));
 MUX2_X1 _2115_ (.A(_0635_),
    .B(\mem[0][23] ),
    .S(_0625_),
    .Z(_0021_));
 BUF_X1 _2116_ (.A(wr_data[24]),
    .Z(_0636_));
 CLKBUF_X2 _2117_ (.A(_0636_),
    .Z(_0637_));
 MUX2_X1 _2118_ (.A(_0637_),
    .B(\mem[0][24] ),
    .S(_0625_),
    .Z(_0022_));
 CLKBUF_X2 _2119_ (.A(wr_data[25]),
    .Z(_0638_));
 BUF_X2 _2120_ (.A(_0638_),
    .Z(_0639_));
 MUX2_X1 _2121_ (.A(_0639_),
    .B(\mem[0][25] ),
    .S(_0625_),
    .Z(_0023_));
 BUF_X1 _2122_ (.A(wr_data[26]),
    .Z(_0640_));
 CLKBUF_X2 _2123_ (.A(_0640_),
    .Z(_0641_));
 MUX2_X1 _2124_ (.A(_0641_),
    .B(\mem[0][26] ),
    .S(_0625_),
    .Z(_0024_));
 CLKBUF_X2 _2125_ (.A(wr_data[27]),
    .Z(_0642_));
 BUF_X2 _2126_ (.A(_0642_),
    .Z(_0643_));
 MUX2_X1 _2127_ (.A(_0643_),
    .B(\mem[0][27] ),
    .S(_0625_),
    .Z(_0025_));
 BUF_X1 _2128_ (.A(wr_data[28]),
    .Z(_0644_));
 BUF_X2 _2129_ (.A(_0644_),
    .Z(_0645_));
 BUF_X4 _2130_ (.A(_0603_),
    .Z(_0646_));
 MUX2_X1 _2131_ (.A(_0645_),
    .B(\mem[0][28] ),
    .S(_0646_),
    .Z(_0026_));
 CLKBUF_X2 _2132_ (.A(wr_data[29]),
    .Z(_0647_));
 BUF_X2 _2133_ (.A(_0647_),
    .Z(_0648_));
 MUX2_X1 _2134_ (.A(_0648_),
    .B(\mem[0][29] ),
    .S(_0646_),
    .Z(_0027_));
 BUF_X1 _2135_ (.A(wr_data[2]),
    .Z(_0649_));
 BUF_X2 _2136_ (.A(_0649_),
    .Z(_0650_));
 MUX2_X1 _2137_ (.A(_0650_),
    .B(\mem[0][2] ),
    .S(_0646_),
    .Z(_0028_));
 BUF_X1 _2138_ (.A(wr_data[30]),
    .Z(_0651_));
 BUF_X2 _2139_ (.A(_0651_),
    .Z(_0652_));
 MUX2_X1 _2140_ (.A(_0652_),
    .B(\mem[0][30] ),
    .S(_0646_),
    .Z(_0029_));
 BUF_X2 _2141_ (.A(wr_data[31]),
    .Z(_0653_));
 BUF_X2 _2142_ (.A(_0653_),
    .Z(_0654_));
 MUX2_X1 _2143_ (.A(_0654_),
    .B(\mem[0][31] ),
    .S(_0646_),
    .Z(_0030_));
 BUF_X1 _2144_ (.A(wr_data[3]),
    .Z(_0655_));
 BUF_X2 _2145_ (.A(_0655_),
    .Z(_0656_));
 MUX2_X1 _2146_ (.A(_0656_),
    .B(\mem[0][3] ),
    .S(_0646_),
    .Z(_0031_));
 BUF_X1 _2147_ (.A(wr_data[4]),
    .Z(_0657_));
 BUF_X2 _2148_ (.A(_0657_),
    .Z(_0658_));
 MUX2_X1 _2149_ (.A(_0658_),
    .B(\mem[0][4] ),
    .S(_0646_),
    .Z(_0032_));
 CLKBUF_X2 _2150_ (.A(wr_data[5]),
    .Z(_0659_));
 BUF_X2 _2151_ (.A(_0659_),
    .Z(_0660_));
 MUX2_X1 _2152_ (.A(_0660_),
    .B(\mem[0][5] ),
    .S(_0646_),
    .Z(_0033_));
 BUF_X1 _2153_ (.A(wr_data[6]),
    .Z(_0661_));
 BUF_X2 _2154_ (.A(_0661_),
    .Z(_0662_));
 MUX2_X1 _2155_ (.A(_0662_),
    .B(\mem[0][6] ),
    .S(_0646_),
    .Z(_0034_));
 BUF_X1 _2156_ (.A(wr_data[7]),
    .Z(_0663_));
 BUF_X2 _2157_ (.A(_0663_),
    .Z(_0664_));
 MUX2_X1 _2158_ (.A(_0664_),
    .B(\mem[0][7] ),
    .S(_0646_),
    .Z(_0035_));
 BUF_X1 _2159_ (.A(wr_data[8]),
    .Z(_0665_));
 BUF_X2 _2160_ (.A(_0665_),
    .Z(_0666_));
 MUX2_X1 _2161_ (.A(_0666_),
    .B(\mem[0][8] ),
    .S(_0603_),
    .Z(_0036_));
 CLKBUF_X2 _2162_ (.A(wr_data[9]),
    .Z(_0667_));
 BUF_X2 _2163_ (.A(_0667_),
    .Z(_0668_));
 MUX2_X1 _2164_ (.A(_0668_),
    .B(\mem[0][9] ),
    .S(_0603_),
    .Z(_0037_));
 INV_X1 _2165_ (.A(_0599_),
    .ZN(_0669_));
 NAND2_X4 _2166_ (.A1(\wr_ptr_bin[3] ),
    .A2(_0669_),
    .ZN(_0670_));
 NAND3_X4 _2167_ (.A1(_1995_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0671_));
 NOR2_X4 _2168_ (.A1(_0670_),
    .A2(_0671_),
    .ZN(_0672_));
 BUF_X4 _2169_ (.A(_0672_),
    .Z(_0673_));
 MUX2_X1 _2170_ (.A(\mem[10][0] ),
    .B(_0598_),
    .S(_0673_),
    .Z(_0038_));
 MUX2_X1 _2171_ (.A(\mem[10][10] ),
    .B(_0606_),
    .S(_0673_),
    .Z(_0039_));
 MUX2_X1 _2172_ (.A(\mem[10][11] ),
    .B(_0608_),
    .S(_0673_),
    .Z(_0040_));
 MUX2_X1 _2173_ (.A(\mem[10][12] ),
    .B(_0610_),
    .S(_0673_),
    .Z(_0041_));
 MUX2_X1 _2174_ (.A(\mem[10][13] ),
    .B(_0612_),
    .S(_0673_),
    .Z(_0042_));
 MUX2_X1 _2175_ (.A(\mem[10][14] ),
    .B(_0614_),
    .S(_0673_),
    .Z(_0043_));
 MUX2_X1 _2176_ (.A(\mem[10][15] ),
    .B(_0616_),
    .S(_0673_),
    .Z(_0044_));
 MUX2_X1 _2177_ (.A(\mem[10][16] ),
    .B(_0618_),
    .S(_0673_),
    .Z(_0045_));
 MUX2_X1 _2178_ (.A(\mem[10][17] ),
    .B(_0620_),
    .S(_0673_),
    .Z(_0046_));
 MUX2_X1 _2179_ (.A(\mem[10][18] ),
    .B(_0622_),
    .S(_0673_),
    .Z(_0047_));
 BUF_X4 _2180_ (.A(_0672_),
    .Z(_0674_));
 MUX2_X1 _2181_ (.A(\mem[10][19] ),
    .B(_0624_),
    .S(_0674_),
    .Z(_0048_));
 MUX2_X1 _2182_ (.A(\mem[10][1] ),
    .B(_0627_),
    .S(_0674_),
    .Z(_0049_));
 MUX2_X1 _2183_ (.A(\mem[10][20] ),
    .B(_0629_),
    .S(_0674_),
    .Z(_0050_));
 MUX2_X1 _2184_ (.A(\mem[10][21] ),
    .B(_0631_),
    .S(_0674_),
    .Z(_0051_));
 MUX2_X1 _2185_ (.A(\mem[10][22] ),
    .B(_0633_),
    .S(_0674_),
    .Z(_0052_));
 MUX2_X1 _2186_ (.A(\mem[10][23] ),
    .B(_0635_),
    .S(_0674_),
    .Z(_0053_));
 MUX2_X1 _2187_ (.A(\mem[10][24] ),
    .B(_0637_),
    .S(_0674_),
    .Z(_0054_));
 MUX2_X1 _2188_ (.A(\mem[10][25] ),
    .B(_0639_),
    .S(_0674_),
    .Z(_0055_));
 MUX2_X1 _2189_ (.A(\mem[10][26] ),
    .B(_0641_),
    .S(_0674_),
    .Z(_0056_));
 MUX2_X1 _2190_ (.A(\mem[10][27] ),
    .B(_0643_),
    .S(_0674_),
    .Z(_0057_));
 BUF_X4 _2191_ (.A(_0672_),
    .Z(_0675_));
 MUX2_X1 _2192_ (.A(\mem[10][28] ),
    .B(_0645_),
    .S(_0675_),
    .Z(_0058_));
 MUX2_X1 _2193_ (.A(\mem[10][29] ),
    .B(_0648_),
    .S(_0675_),
    .Z(_0059_));
 MUX2_X1 _2194_ (.A(\mem[10][2] ),
    .B(_0650_),
    .S(_0675_),
    .Z(_0060_));
 MUX2_X1 _2195_ (.A(\mem[10][30] ),
    .B(_0652_),
    .S(_0675_),
    .Z(_0061_));
 MUX2_X1 _2196_ (.A(\mem[10][31] ),
    .B(_0654_),
    .S(_0675_),
    .Z(_0062_));
 MUX2_X1 _2197_ (.A(\mem[10][3] ),
    .B(_0656_),
    .S(_0675_),
    .Z(_0063_));
 MUX2_X1 _2198_ (.A(\mem[10][4] ),
    .B(_0658_),
    .S(_0675_),
    .Z(_0064_));
 MUX2_X1 _2199_ (.A(\mem[10][5] ),
    .B(_0660_),
    .S(_0675_),
    .Z(_0065_));
 MUX2_X1 _2200_ (.A(\mem[10][6] ),
    .B(_0662_),
    .S(_0675_),
    .Z(_0066_));
 MUX2_X1 _2201_ (.A(\mem[10][7] ),
    .B(_0664_),
    .S(_0675_),
    .Z(_0067_));
 MUX2_X1 _2202_ (.A(\mem[10][8] ),
    .B(_0666_),
    .S(_0672_),
    .Z(_0068_));
 MUX2_X1 _2203_ (.A(\mem[10][9] ),
    .B(_0668_),
    .S(_0672_),
    .Z(_0069_));
 NAND3_X4 _2204_ (.A1(_1999_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0676_));
 NOR2_X4 _2205_ (.A1(_0670_),
    .A2(_0676_),
    .ZN(_0677_));
 BUF_X4 _2206_ (.A(_0677_),
    .Z(_0678_));
 MUX2_X1 _2207_ (.A(\mem[11][0] ),
    .B(_0598_),
    .S(_0678_),
    .Z(_0070_));
 MUX2_X1 _2208_ (.A(\mem[11][10] ),
    .B(_0606_),
    .S(_0678_),
    .Z(_0071_));
 MUX2_X1 _2209_ (.A(\mem[11][11] ),
    .B(_0608_),
    .S(_0678_),
    .Z(_0072_));
 MUX2_X1 _2210_ (.A(\mem[11][12] ),
    .B(_0610_),
    .S(_0678_),
    .Z(_0073_));
 MUX2_X1 _2211_ (.A(\mem[11][13] ),
    .B(_0612_),
    .S(_0678_),
    .Z(_0074_));
 MUX2_X1 _2212_ (.A(\mem[11][14] ),
    .B(_0614_),
    .S(_0678_),
    .Z(_0075_));
 MUX2_X1 _2213_ (.A(\mem[11][15] ),
    .B(_0616_),
    .S(_0678_),
    .Z(_0076_));
 MUX2_X1 _2214_ (.A(\mem[11][16] ),
    .B(_0618_),
    .S(_0678_),
    .Z(_0077_));
 MUX2_X1 _2215_ (.A(\mem[11][17] ),
    .B(_0620_),
    .S(_0678_),
    .Z(_0078_));
 MUX2_X1 _2216_ (.A(\mem[11][18] ),
    .B(_0622_),
    .S(_0678_),
    .Z(_0079_));
 BUF_X4 _2217_ (.A(_0677_),
    .Z(_0679_));
 MUX2_X1 _2218_ (.A(\mem[11][19] ),
    .B(_0624_),
    .S(_0679_),
    .Z(_0080_));
 MUX2_X1 _2219_ (.A(\mem[11][1] ),
    .B(_0627_),
    .S(_0679_),
    .Z(_0081_));
 MUX2_X1 _2220_ (.A(\mem[11][20] ),
    .B(_0629_),
    .S(_0679_),
    .Z(_0082_));
 MUX2_X1 _2221_ (.A(\mem[11][21] ),
    .B(_0631_),
    .S(_0679_),
    .Z(_0083_));
 MUX2_X1 _2222_ (.A(\mem[11][22] ),
    .B(_0633_),
    .S(_0679_),
    .Z(_0084_));
 MUX2_X1 _2223_ (.A(\mem[11][23] ),
    .B(_0635_),
    .S(_0679_),
    .Z(_0085_));
 MUX2_X1 _2224_ (.A(\mem[11][24] ),
    .B(_0637_),
    .S(_0679_),
    .Z(_0086_));
 MUX2_X1 _2225_ (.A(\mem[11][25] ),
    .B(_0639_),
    .S(_0679_),
    .Z(_0087_));
 MUX2_X1 _2226_ (.A(\mem[11][26] ),
    .B(_0641_),
    .S(_0679_),
    .Z(_0088_));
 MUX2_X1 _2227_ (.A(\mem[11][27] ),
    .B(_0643_),
    .S(_0679_),
    .Z(_0089_));
 BUF_X4 _2228_ (.A(_0677_),
    .Z(_0680_));
 MUX2_X1 _2229_ (.A(\mem[11][28] ),
    .B(_0645_),
    .S(_0680_),
    .Z(_0090_));
 MUX2_X1 _2230_ (.A(\mem[11][29] ),
    .B(_0648_),
    .S(_0680_),
    .Z(_0091_));
 MUX2_X1 _2231_ (.A(\mem[11][2] ),
    .B(_0650_),
    .S(_0680_),
    .Z(_0092_));
 MUX2_X1 _2232_ (.A(\mem[11][30] ),
    .B(_0652_),
    .S(_0680_),
    .Z(_0093_));
 MUX2_X1 _2233_ (.A(\mem[11][31] ),
    .B(_0654_),
    .S(_0680_),
    .Z(_0094_));
 MUX2_X1 _2234_ (.A(\mem[11][3] ),
    .B(_0656_),
    .S(_0680_),
    .Z(_0095_));
 MUX2_X1 _2235_ (.A(\mem[11][4] ),
    .B(_0658_),
    .S(_0680_),
    .Z(_0096_));
 MUX2_X1 _2236_ (.A(\mem[11][5] ),
    .B(_0660_),
    .S(_0680_),
    .Z(_0097_));
 MUX2_X1 _2237_ (.A(\mem[11][6] ),
    .B(_0662_),
    .S(_0680_),
    .Z(_0098_));
 MUX2_X1 _2238_ (.A(\mem[11][7] ),
    .B(_0664_),
    .S(_0680_),
    .Z(_0099_));
 MUX2_X1 _2239_ (.A(\mem[11][8] ),
    .B(_0666_),
    .S(_0677_),
    .Z(_0100_));
 MUX2_X1 _2240_ (.A(\mem[11][9] ),
    .B(_0668_),
    .S(_0677_),
    .Z(_0101_));
 AND2_X1 _2241_ (.A1(\wr_ptr_bin[3] ),
    .A2(_0599_),
    .ZN(_0681_));
 BUF_X4 _2242_ (.A(_0681_),
    .Z(_0682_));
 NAND2_X4 _2243_ (.A1(_0602_),
    .A2(_0682_),
    .ZN(_0683_));
 BUF_X4 _2244_ (.A(_0683_),
    .Z(_0684_));
 MUX2_X1 _2245_ (.A(_0598_),
    .B(\mem[12][0] ),
    .S(_0684_),
    .Z(_0102_));
 MUX2_X1 _2246_ (.A(_0606_),
    .B(\mem[12][10] ),
    .S(_0684_),
    .Z(_0103_));
 MUX2_X1 _2247_ (.A(_0608_),
    .B(\mem[12][11] ),
    .S(_0684_),
    .Z(_0104_));
 MUX2_X1 _2248_ (.A(_0610_),
    .B(\mem[12][12] ),
    .S(_0684_),
    .Z(_0105_));
 MUX2_X1 _2249_ (.A(_0612_),
    .B(\mem[12][13] ),
    .S(_0684_),
    .Z(_0106_));
 MUX2_X1 _2250_ (.A(_0614_),
    .B(\mem[12][14] ),
    .S(_0684_),
    .Z(_0107_));
 MUX2_X1 _2251_ (.A(_0616_),
    .B(\mem[12][15] ),
    .S(_0684_),
    .Z(_0108_));
 MUX2_X1 _2252_ (.A(_0618_),
    .B(\mem[12][16] ),
    .S(_0684_),
    .Z(_0109_));
 MUX2_X1 _2253_ (.A(_0620_),
    .B(\mem[12][17] ),
    .S(_0684_),
    .Z(_0110_));
 MUX2_X1 _2254_ (.A(_0622_),
    .B(\mem[12][18] ),
    .S(_0684_),
    .Z(_0111_));
 BUF_X4 _2255_ (.A(_0683_),
    .Z(_0685_));
 MUX2_X1 _2256_ (.A(_0624_),
    .B(\mem[12][19] ),
    .S(_0685_),
    .Z(_0112_));
 MUX2_X1 _2257_ (.A(_0627_),
    .B(\mem[12][1] ),
    .S(_0685_),
    .Z(_0113_));
 MUX2_X1 _2258_ (.A(_0629_),
    .B(\mem[12][20] ),
    .S(_0685_),
    .Z(_0114_));
 MUX2_X1 _2259_ (.A(_0631_),
    .B(\mem[12][21] ),
    .S(_0685_),
    .Z(_0115_));
 MUX2_X1 _2260_ (.A(_0633_),
    .B(\mem[12][22] ),
    .S(_0685_),
    .Z(_0116_));
 MUX2_X1 _2261_ (.A(_0635_),
    .B(\mem[12][23] ),
    .S(_0685_),
    .Z(_0117_));
 MUX2_X1 _2262_ (.A(_0637_),
    .B(\mem[12][24] ),
    .S(_0685_),
    .Z(_0118_));
 MUX2_X1 _2263_ (.A(_0639_),
    .B(\mem[12][25] ),
    .S(_0685_),
    .Z(_0119_));
 MUX2_X1 _2264_ (.A(_0641_),
    .B(\mem[12][26] ),
    .S(_0685_),
    .Z(_0120_));
 MUX2_X1 _2265_ (.A(_0643_),
    .B(\mem[12][27] ),
    .S(_0685_),
    .Z(_0121_));
 BUF_X4 _2266_ (.A(_0683_),
    .Z(_0686_));
 MUX2_X1 _2267_ (.A(_0645_),
    .B(\mem[12][28] ),
    .S(_0686_),
    .Z(_0122_));
 MUX2_X1 _2268_ (.A(_0648_),
    .B(\mem[12][29] ),
    .S(_0686_),
    .Z(_0123_));
 MUX2_X1 _2269_ (.A(_0650_),
    .B(\mem[12][2] ),
    .S(_0686_),
    .Z(_0124_));
 MUX2_X1 _2270_ (.A(_0652_),
    .B(\mem[12][30] ),
    .S(_0686_),
    .Z(_0125_));
 MUX2_X1 _2271_ (.A(_0654_),
    .B(\mem[12][31] ),
    .S(_0686_),
    .Z(_0126_));
 MUX2_X1 _2272_ (.A(_0656_),
    .B(\mem[12][3] ),
    .S(_0686_),
    .Z(_0127_));
 MUX2_X1 _2273_ (.A(_0658_),
    .B(\mem[12][4] ),
    .S(_0686_),
    .Z(_0128_));
 MUX2_X1 _2274_ (.A(_0660_),
    .B(\mem[12][5] ),
    .S(_0686_),
    .Z(_0129_));
 MUX2_X1 _2275_ (.A(_0662_),
    .B(\mem[12][6] ),
    .S(_0686_),
    .Z(_0130_));
 MUX2_X1 _2276_ (.A(_0664_),
    .B(\mem[12][7] ),
    .S(_0686_),
    .Z(_0131_));
 MUX2_X1 _2277_ (.A(_0666_),
    .B(\mem[12][8] ),
    .S(_0683_),
    .Z(_0132_));
 MUX2_X1 _2278_ (.A(_0668_),
    .B(\mem[12][9] ),
    .S(_0683_),
    .Z(_0133_));
 AND3_X2 _2279_ (.A1(_1997_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0687_));
 NAND2_X4 _2280_ (.A1(_0682_),
    .A2(_0687_),
    .ZN(_0688_));
 BUF_X4 _2281_ (.A(_0688_),
    .Z(_0689_));
 MUX2_X1 _2282_ (.A(_0597_),
    .B(\mem[13][0] ),
    .S(_0689_),
    .Z(_0134_));
 MUX2_X1 _2283_ (.A(_0605_),
    .B(\mem[13][10] ),
    .S(_0689_),
    .Z(_0135_));
 MUX2_X1 _2284_ (.A(_0607_),
    .B(\mem[13][11] ),
    .S(_0689_),
    .Z(_0136_));
 MUX2_X1 _2285_ (.A(_0609_),
    .B(\mem[13][12] ),
    .S(_0689_),
    .Z(_0137_));
 MUX2_X1 _2286_ (.A(_0611_),
    .B(\mem[13][13] ),
    .S(_0689_),
    .Z(_0138_));
 MUX2_X1 _2287_ (.A(_0613_),
    .B(\mem[13][14] ),
    .S(_0689_),
    .Z(_0139_));
 MUX2_X1 _2288_ (.A(_0615_),
    .B(\mem[13][15] ),
    .S(_0689_),
    .Z(_0140_));
 MUX2_X1 _2289_ (.A(_0617_),
    .B(\mem[13][16] ),
    .S(_0689_),
    .Z(_0141_));
 MUX2_X1 _2290_ (.A(_0619_),
    .B(\mem[13][17] ),
    .S(_0689_),
    .Z(_0142_));
 MUX2_X1 _2291_ (.A(_0621_),
    .B(\mem[13][18] ),
    .S(_0689_),
    .Z(_0143_));
 BUF_X4 _2292_ (.A(_0688_),
    .Z(_0690_));
 MUX2_X1 _2293_ (.A(_0623_),
    .B(\mem[13][19] ),
    .S(_0690_),
    .Z(_0144_));
 MUX2_X1 _2294_ (.A(_0626_),
    .B(\mem[13][1] ),
    .S(_0690_),
    .Z(_0145_));
 MUX2_X1 _2295_ (.A(_0628_),
    .B(\mem[13][20] ),
    .S(_0690_),
    .Z(_0146_));
 MUX2_X1 _2296_ (.A(_0630_),
    .B(\mem[13][21] ),
    .S(_0690_),
    .Z(_0147_));
 MUX2_X1 _2297_ (.A(_0632_),
    .B(\mem[13][22] ),
    .S(_0690_),
    .Z(_0148_));
 MUX2_X1 _2298_ (.A(_0634_),
    .B(\mem[13][23] ),
    .S(_0690_),
    .Z(_0149_));
 MUX2_X1 _2299_ (.A(_0636_),
    .B(\mem[13][24] ),
    .S(_0690_),
    .Z(_0150_));
 MUX2_X1 _2300_ (.A(_0638_),
    .B(\mem[13][25] ),
    .S(_0690_),
    .Z(_0151_));
 MUX2_X1 _2301_ (.A(_0640_),
    .B(\mem[13][26] ),
    .S(_0690_),
    .Z(_0152_));
 MUX2_X1 _2302_ (.A(_0642_),
    .B(\mem[13][27] ),
    .S(_0690_),
    .Z(_0153_));
 BUF_X4 _2303_ (.A(_0688_),
    .Z(_0691_));
 MUX2_X1 _2304_ (.A(_0644_),
    .B(\mem[13][28] ),
    .S(_0691_),
    .Z(_0154_));
 MUX2_X1 _2305_ (.A(_0647_),
    .B(\mem[13][29] ),
    .S(_0691_),
    .Z(_0155_));
 MUX2_X1 _2306_ (.A(_0649_),
    .B(\mem[13][2] ),
    .S(_0691_),
    .Z(_0156_));
 MUX2_X1 _2307_ (.A(_0651_),
    .B(\mem[13][30] ),
    .S(_0691_),
    .Z(_0157_));
 MUX2_X1 _2308_ (.A(_0653_),
    .B(\mem[13][31] ),
    .S(_0691_),
    .Z(_0158_));
 MUX2_X1 _2309_ (.A(_0655_),
    .B(\mem[13][3] ),
    .S(_0691_),
    .Z(_0159_));
 MUX2_X1 _2310_ (.A(_0657_),
    .B(\mem[13][4] ),
    .S(_0691_),
    .Z(_0160_));
 MUX2_X1 _2311_ (.A(_0659_),
    .B(\mem[13][5] ),
    .S(_0691_),
    .Z(_0161_));
 MUX2_X1 _2312_ (.A(_0661_),
    .B(\mem[13][6] ),
    .S(_0691_),
    .Z(_0162_));
 MUX2_X1 _2313_ (.A(_0663_),
    .B(\mem[13][7] ),
    .S(_0691_),
    .Z(_0163_));
 MUX2_X1 _2314_ (.A(_0665_),
    .B(\mem[13][8] ),
    .S(_0688_),
    .Z(_0164_));
 MUX2_X1 _2315_ (.A(_0667_),
    .B(\mem[13][9] ),
    .S(_0688_),
    .Z(_0165_));
 AND3_X2 _2316_ (.A1(_1995_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0692_));
 NAND2_X4 _2317_ (.A1(_0692_),
    .A2(_0682_),
    .ZN(_0693_));
 BUF_X4 _2318_ (.A(_0693_),
    .Z(_0694_));
 MUX2_X1 _2319_ (.A(_0597_),
    .B(\mem[14][0] ),
    .S(_0694_),
    .Z(_0166_));
 MUX2_X1 _2320_ (.A(_0605_),
    .B(\mem[14][10] ),
    .S(_0694_),
    .Z(_0167_));
 MUX2_X1 _2321_ (.A(_0607_),
    .B(\mem[14][11] ),
    .S(_0694_),
    .Z(_0168_));
 MUX2_X1 _2322_ (.A(_0609_),
    .B(\mem[14][12] ),
    .S(_0694_),
    .Z(_0169_));
 MUX2_X1 _2323_ (.A(_0611_),
    .B(\mem[14][13] ),
    .S(_0694_),
    .Z(_0170_));
 MUX2_X1 _2324_ (.A(_0613_),
    .B(\mem[14][14] ),
    .S(_0694_),
    .Z(_0171_));
 MUX2_X1 _2325_ (.A(_0615_),
    .B(\mem[14][15] ),
    .S(_0694_),
    .Z(_0172_));
 MUX2_X1 _2326_ (.A(_0617_),
    .B(\mem[14][16] ),
    .S(_0694_),
    .Z(_0173_));
 MUX2_X1 _2327_ (.A(_0619_),
    .B(\mem[14][17] ),
    .S(_0694_),
    .Z(_0174_));
 MUX2_X1 _2328_ (.A(_0621_),
    .B(\mem[14][18] ),
    .S(_0694_),
    .Z(_0175_));
 BUF_X4 _2329_ (.A(_0693_),
    .Z(_0695_));
 MUX2_X1 _2330_ (.A(_0623_),
    .B(\mem[14][19] ),
    .S(_0695_),
    .Z(_0176_));
 MUX2_X1 _2331_ (.A(_0626_),
    .B(\mem[14][1] ),
    .S(_0695_),
    .Z(_0177_));
 MUX2_X1 _2332_ (.A(_0628_),
    .B(\mem[14][20] ),
    .S(_0695_),
    .Z(_0178_));
 MUX2_X1 _2333_ (.A(_0630_),
    .B(\mem[14][21] ),
    .S(_0695_),
    .Z(_0179_));
 MUX2_X1 _2334_ (.A(_0632_),
    .B(\mem[14][22] ),
    .S(_0695_),
    .Z(_0180_));
 MUX2_X1 _2335_ (.A(_0634_),
    .B(\mem[14][23] ),
    .S(_0695_),
    .Z(_0181_));
 MUX2_X1 _2336_ (.A(_0636_),
    .B(\mem[14][24] ),
    .S(_0695_),
    .Z(_0182_));
 MUX2_X1 _2337_ (.A(_0638_),
    .B(\mem[14][25] ),
    .S(_0695_),
    .Z(_0183_));
 MUX2_X1 _2338_ (.A(_0640_),
    .B(\mem[14][26] ),
    .S(_0695_),
    .Z(_0184_));
 MUX2_X1 _2339_ (.A(_0642_),
    .B(\mem[14][27] ),
    .S(_0695_),
    .Z(_0185_));
 BUF_X4 _2340_ (.A(_0693_),
    .Z(_0696_));
 MUX2_X1 _2341_ (.A(_0644_),
    .B(\mem[14][28] ),
    .S(_0696_),
    .Z(_0186_));
 MUX2_X1 _2342_ (.A(_0647_),
    .B(\mem[14][29] ),
    .S(_0696_),
    .Z(_0187_));
 MUX2_X1 _2343_ (.A(_0649_),
    .B(\mem[14][2] ),
    .S(_0696_),
    .Z(_0188_));
 MUX2_X1 _2344_ (.A(_0651_),
    .B(\mem[14][30] ),
    .S(_0696_),
    .Z(_0189_));
 MUX2_X1 _2345_ (.A(_0653_),
    .B(\mem[14][31] ),
    .S(_0696_),
    .Z(_0190_));
 MUX2_X1 _2346_ (.A(_0655_),
    .B(\mem[14][3] ),
    .S(_0696_),
    .Z(_0191_));
 MUX2_X1 _2347_ (.A(_0657_),
    .B(\mem[14][4] ),
    .S(_0696_),
    .Z(_0192_));
 MUX2_X1 _2348_ (.A(_0659_),
    .B(\mem[14][5] ),
    .S(_0696_),
    .Z(_0193_));
 MUX2_X1 _2349_ (.A(_0661_),
    .B(\mem[14][6] ),
    .S(_0696_),
    .Z(_0194_));
 MUX2_X1 _2350_ (.A(_0663_),
    .B(\mem[14][7] ),
    .S(_0696_),
    .Z(_0195_));
 MUX2_X1 _2351_ (.A(_0665_),
    .B(\mem[14][8] ),
    .S(_0693_),
    .Z(_0196_));
 MUX2_X1 _2352_ (.A(_0667_),
    .B(\mem[14][9] ),
    .S(_0693_),
    .Z(_0197_));
 AND3_X2 _2353_ (.A1(_1999_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0697_));
 NAND2_X4 _2354_ (.A1(_0697_),
    .A2(_0682_),
    .ZN(_0698_));
 BUF_X4 _2355_ (.A(_0698_),
    .Z(_0699_));
 MUX2_X1 _2356_ (.A(_0597_),
    .B(\mem[15][0] ),
    .S(_0699_),
    .Z(_0198_));
 MUX2_X1 _2357_ (.A(_0605_),
    .B(\mem[15][10] ),
    .S(_0699_),
    .Z(_0199_));
 MUX2_X1 _2358_ (.A(_0607_),
    .B(\mem[15][11] ),
    .S(_0699_),
    .Z(_0200_));
 MUX2_X1 _2359_ (.A(_0609_),
    .B(\mem[15][12] ),
    .S(_0699_),
    .Z(_0201_));
 MUX2_X1 _2360_ (.A(_0611_),
    .B(\mem[15][13] ),
    .S(_0699_),
    .Z(_0202_));
 MUX2_X1 _2361_ (.A(_0613_),
    .B(\mem[15][14] ),
    .S(_0699_),
    .Z(_0203_));
 MUX2_X1 _2362_ (.A(_0615_),
    .B(\mem[15][15] ),
    .S(_0699_),
    .Z(_0204_));
 MUX2_X1 _2363_ (.A(_0617_),
    .B(\mem[15][16] ),
    .S(_0699_),
    .Z(_0205_));
 MUX2_X1 _2364_ (.A(_0619_),
    .B(\mem[15][17] ),
    .S(_0699_),
    .Z(_0206_));
 MUX2_X1 _2365_ (.A(_0621_),
    .B(\mem[15][18] ),
    .S(_0699_),
    .Z(_0207_));
 BUF_X4 _2366_ (.A(_0698_),
    .Z(_0700_));
 MUX2_X1 _2367_ (.A(_0623_),
    .B(\mem[15][19] ),
    .S(_0700_),
    .Z(_0208_));
 MUX2_X1 _2368_ (.A(_0626_),
    .B(\mem[15][1] ),
    .S(_0700_),
    .Z(_0209_));
 MUX2_X1 _2369_ (.A(_0628_),
    .B(\mem[15][20] ),
    .S(_0700_),
    .Z(_0210_));
 MUX2_X1 _2370_ (.A(_0630_),
    .B(\mem[15][21] ),
    .S(_0700_),
    .Z(_0211_));
 MUX2_X1 _2371_ (.A(_0632_),
    .B(\mem[15][22] ),
    .S(_0700_),
    .Z(_0212_));
 MUX2_X1 _2372_ (.A(_0634_),
    .B(\mem[15][23] ),
    .S(_0700_),
    .Z(_0213_));
 MUX2_X1 _2373_ (.A(_0636_),
    .B(\mem[15][24] ),
    .S(_0700_),
    .Z(_0214_));
 MUX2_X1 _2374_ (.A(_0638_),
    .B(\mem[15][25] ),
    .S(_0700_),
    .Z(_0215_));
 MUX2_X1 _2375_ (.A(_0640_),
    .B(\mem[15][26] ),
    .S(_0700_),
    .Z(_0216_));
 MUX2_X1 _2376_ (.A(_0642_),
    .B(\mem[15][27] ),
    .S(_0700_),
    .Z(_0217_));
 BUF_X4 _2377_ (.A(_0698_),
    .Z(_0701_));
 MUX2_X1 _2378_ (.A(_0644_),
    .B(\mem[15][28] ),
    .S(_0701_),
    .Z(_0218_));
 MUX2_X1 _2379_ (.A(_0647_),
    .B(\mem[15][29] ),
    .S(_0701_),
    .Z(_0219_));
 MUX2_X1 _2380_ (.A(_0649_),
    .B(\mem[15][2] ),
    .S(_0701_),
    .Z(_0220_));
 MUX2_X1 _2381_ (.A(_0651_),
    .B(\mem[15][30] ),
    .S(_0701_),
    .Z(_0221_));
 MUX2_X1 _2382_ (.A(_0653_),
    .B(\mem[15][31] ),
    .S(_0701_),
    .Z(_0222_));
 MUX2_X1 _2383_ (.A(_0655_),
    .B(\mem[15][3] ),
    .S(_0701_),
    .Z(_0223_));
 MUX2_X1 _2384_ (.A(_0657_),
    .B(\mem[15][4] ),
    .S(_0701_),
    .Z(_0224_));
 MUX2_X1 _2385_ (.A(_0659_),
    .B(\mem[15][5] ),
    .S(_0701_),
    .Z(_0225_));
 MUX2_X1 _2386_ (.A(_0661_),
    .B(\mem[15][6] ),
    .S(_0701_),
    .Z(_0226_));
 MUX2_X1 _2387_ (.A(_0663_),
    .B(\mem[15][7] ),
    .S(_0701_),
    .Z(_0227_));
 MUX2_X1 _2388_ (.A(_0665_),
    .B(\mem[15][8] ),
    .S(_0698_),
    .Z(_0228_));
 MUX2_X1 _2389_ (.A(_0667_),
    .B(\mem[15][9] ),
    .S(_0698_),
    .Z(_0229_));
 NAND2_X4 _2390_ (.A1(_0600_),
    .A2(_0687_),
    .ZN(_0702_));
 BUF_X4 _2391_ (.A(_0702_),
    .Z(_0703_));
 MUX2_X1 _2392_ (.A(_0597_),
    .B(\mem[1][0] ),
    .S(_0703_),
    .Z(_0230_));
 MUX2_X1 _2393_ (.A(_0605_),
    .B(\mem[1][10] ),
    .S(_0703_),
    .Z(_0231_));
 MUX2_X1 _2394_ (.A(_0607_),
    .B(\mem[1][11] ),
    .S(_0703_),
    .Z(_0232_));
 MUX2_X1 _2395_ (.A(_0609_),
    .B(\mem[1][12] ),
    .S(_0703_),
    .Z(_0233_));
 MUX2_X1 _2396_ (.A(_0611_),
    .B(\mem[1][13] ),
    .S(_0703_),
    .Z(_0234_));
 MUX2_X1 _2397_ (.A(_0613_),
    .B(\mem[1][14] ),
    .S(_0703_),
    .Z(_0235_));
 MUX2_X1 _2398_ (.A(_0615_),
    .B(\mem[1][15] ),
    .S(_0703_),
    .Z(_0236_));
 MUX2_X1 _2399_ (.A(_0617_),
    .B(\mem[1][16] ),
    .S(_0703_),
    .Z(_0237_));
 MUX2_X1 _2400_ (.A(_0619_),
    .B(\mem[1][17] ),
    .S(_0703_),
    .Z(_0238_));
 MUX2_X1 _2401_ (.A(_0621_),
    .B(\mem[1][18] ),
    .S(_0703_),
    .Z(_0239_));
 BUF_X4 _2402_ (.A(_0702_),
    .Z(_0704_));
 MUX2_X1 _2403_ (.A(_0623_),
    .B(\mem[1][19] ),
    .S(_0704_),
    .Z(_0240_));
 MUX2_X1 _2404_ (.A(_0626_),
    .B(\mem[1][1] ),
    .S(_0704_),
    .Z(_0241_));
 MUX2_X1 _2405_ (.A(_0628_),
    .B(\mem[1][20] ),
    .S(_0704_),
    .Z(_0242_));
 MUX2_X1 _2406_ (.A(_0630_),
    .B(\mem[1][21] ),
    .S(_0704_),
    .Z(_0243_));
 MUX2_X1 _2407_ (.A(_0632_),
    .B(\mem[1][22] ),
    .S(_0704_),
    .Z(_0244_));
 MUX2_X1 _2408_ (.A(_0634_),
    .B(\mem[1][23] ),
    .S(_0704_),
    .Z(_0245_));
 MUX2_X1 _2409_ (.A(_0636_),
    .B(\mem[1][24] ),
    .S(_0704_),
    .Z(_0246_));
 MUX2_X1 _2410_ (.A(_0638_),
    .B(\mem[1][25] ),
    .S(_0704_),
    .Z(_0247_));
 MUX2_X1 _2411_ (.A(_0640_),
    .B(\mem[1][26] ),
    .S(_0704_),
    .Z(_0248_));
 MUX2_X1 _2412_ (.A(_0642_),
    .B(\mem[1][27] ),
    .S(_0704_),
    .Z(_0249_));
 BUF_X4 _2413_ (.A(_0702_),
    .Z(_0705_));
 MUX2_X1 _2414_ (.A(_0644_),
    .B(\mem[1][28] ),
    .S(_0705_),
    .Z(_0250_));
 MUX2_X1 _2415_ (.A(_0647_),
    .B(\mem[1][29] ),
    .S(_0705_),
    .Z(_0251_));
 MUX2_X1 _2416_ (.A(_0649_),
    .B(\mem[1][2] ),
    .S(_0705_),
    .Z(_0252_));
 MUX2_X1 _2417_ (.A(_0651_),
    .B(\mem[1][30] ),
    .S(_0705_),
    .Z(_0253_));
 MUX2_X1 _2418_ (.A(_0653_),
    .B(\mem[1][31] ),
    .S(_0705_),
    .Z(_0254_));
 MUX2_X1 _2419_ (.A(_0655_),
    .B(\mem[1][3] ),
    .S(_0705_),
    .Z(_0255_));
 MUX2_X1 _2420_ (.A(_0657_),
    .B(\mem[1][4] ),
    .S(_0705_),
    .Z(_0256_));
 MUX2_X1 _2421_ (.A(_0659_),
    .B(\mem[1][5] ),
    .S(_0705_),
    .Z(_0257_));
 MUX2_X1 _2422_ (.A(_0661_),
    .B(\mem[1][6] ),
    .S(_0705_),
    .Z(_0258_));
 MUX2_X1 _2423_ (.A(_0663_),
    .B(\mem[1][7] ),
    .S(_0705_),
    .Z(_0259_));
 MUX2_X1 _2424_ (.A(_0665_),
    .B(\mem[1][8] ),
    .S(_0702_),
    .Z(_0260_));
 MUX2_X1 _2425_ (.A(_0667_),
    .B(\mem[1][9] ),
    .S(_0702_),
    .Z(_0261_));
 NAND2_X4 _2426_ (.A1(_0600_),
    .A2(_0692_),
    .ZN(_0706_));
 BUF_X4 _2427_ (.A(_0706_),
    .Z(_0707_));
 MUX2_X1 _2428_ (.A(_0597_),
    .B(\mem[2][0] ),
    .S(_0707_),
    .Z(_0262_));
 MUX2_X1 _2429_ (.A(_0605_),
    .B(\mem[2][10] ),
    .S(_0707_),
    .Z(_0263_));
 MUX2_X1 _2430_ (.A(_0607_),
    .B(\mem[2][11] ),
    .S(_0707_),
    .Z(_0264_));
 MUX2_X1 _2431_ (.A(_0609_),
    .B(\mem[2][12] ),
    .S(_0707_),
    .Z(_0265_));
 MUX2_X1 _2432_ (.A(_0611_),
    .B(\mem[2][13] ),
    .S(_0707_),
    .Z(_0266_));
 MUX2_X1 _2433_ (.A(_0613_),
    .B(\mem[2][14] ),
    .S(_0707_),
    .Z(_0267_));
 MUX2_X1 _2434_ (.A(_0615_),
    .B(\mem[2][15] ),
    .S(_0707_),
    .Z(_0268_));
 MUX2_X1 _2435_ (.A(_0617_),
    .B(\mem[2][16] ),
    .S(_0707_),
    .Z(_0269_));
 MUX2_X1 _2436_ (.A(_0619_),
    .B(\mem[2][17] ),
    .S(_0707_),
    .Z(_0270_));
 MUX2_X1 _2437_ (.A(_0621_),
    .B(\mem[2][18] ),
    .S(_0707_),
    .Z(_0271_));
 BUF_X4 _2438_ (.A(_0706_),
    .Z(_0708_));
 MUX2_X1 _2439_ (.A(_0623_),
    .B(\mem[2][19] ),
    .S(_0708_),
    .Z(_0272_));
 MUX2_X1 _2440_ (.A(_0626_),
    .B(\mem[2][1] ),
    .S(_0708_),
    .Z(_0273_));
 MUX2_X1 _2441_ (.A(_0628_),
    .B(\mem[2][20] ),
    .S(_0708_),
    .Z(_0274_));
 MUX2_X1 _2442_ (.A(_0630_),
    .B(\mem[2][21] ),
    .S(_0708_),
    .Z(_0275_));
 MUX2_X1 _2443_ (.A(_0632_),
    .B(\mem[2][22] ),
    .S(_0708_),
    .Z(_0276_));
 MUX2_X1 _2444_ (.A(_0634_),
    .B(\mem[2][23] ),
    .S(_0708_),
    .Z(_0277_));
 MUX2_X1 _2445_ (.A(_0636_),
    .B(\mem[2][24] ),
    .S(_0708_),
    .Z(_0278_));
 MUX2_X1 _2446_ (.A(_0638_),
    .B(\mem[2][25] ),
    .S(_0708_),
    .Z(_0279_));
 MUX2_X1 _2447_ (.A(_0640_),
    .B(\mem[2][26] ),
    .S(_0708_),
    .Z(_0280_));
 MUX2_X1 _2448_ (.A(_0642_),
    .B(\mem[2][27] ),
    .S(_0708_),
    .Z(_0281_));
 BUF_X4 _2449_ (.A(_0706_),
    .Z(_0709_));
 MUX2_X1 _2450_ (.A(_0644_),
    .B(\mem[2][28] ),
    .S(_0709_),
    .Z(_0282_));
 MUX2_X1 _2451_ (.A(_0647_),
    .B(\mem[2][29] ),
    .S(_0709_),
    .Z(_0283_));
 MUX2_X1 _2452_ (.A(_0649_),
    .B(\mem[2][2] ),
    .S(_0709_),
    .Z(_0284_));
 MUX2_X1 _2453_ (.A(_0651_),
    .B(\mem[2][30] ),
    .S(_0709_),
    .Z(_0285_));
 MUX2_X1 _2454_ (.A(_0653_),
    .B(\mem[2][31] ),
    .S(_0709_),
    .Z(_0286_));
 MUX2_X1 _2455_ (.A(_0655_),
    .B(\mem[2][3] ),
    .S(_0709_),
    .Z(_0287_));
 MUX2_X1 _2456_ (.A(_0657_),
    .B(\mem[2][4] ),
    .S(_0709_),
    .Z(_0288_));
 MUX2_X1 _2457_ (.A(_0659_),
    .B(\mem[2][5] ),
    .S(_0709_),
    .Z(_0289_));
 MUX2_X1 _2458_ (.A(_0661_),
    .B(\mem[2][6] ),
    .S(_0709_),
    .Z(_0290_));
 MUX2_X1 _2459_ (.A(_0663_),
    .B(\mem[2][7] ),
    .S(_0709_),
    .Z(_0291_));
 MUX2_X1 _2460_ (.A(_0665_),
    .B(\mem[2][8] ),
    .S(_0706_),
    .Z(_0292_));
 MUX2_X1 _2461_ (.A(_0667_),
    .B(\mem[2][9] ),
    .S(_0706_),
    .Z(_0293_));
 NAND2_X4 _2462_ (.A1(_0600_),
    .A2(_0697_),
    .ZN(_0710_));
 BUF_X4 _2463_ (.A(_0710_),
    .Z(_0711_));
 MUX2_X1 _2464_ (.A(_0597_),
    .B(\mem[3][0] ),
    .S(_0711_),
    .Z(_0294_));
 MUX2_X1 _2465_ (.A(_0605_),
    .B(\mem[3][10] ),
    .S(_0711_),
    .Z(_0295_));
 MUX2_X1 _2466_ (.A(_0607_),
    .B(\mem[3][11] ),
    .S(_0711_),
    .Z(_0296_));
 MUX2_X1 _2467_ (.A(_0609_),
    .B(\mem[3][12] ),
    .S(_0711_),
    .Z(_0297_));
 MUX2_X1 _2468_ (.A(_0611_),
    .B(\mem[3][13] ),
    .S(_0711_),
    .Z(_0298_));
 MUX2_X1 _2469_ (.A(_0613_),
    .B(\mem[3][14] ),
    .S(_0711_),
    .Z(_0299_));
 MUX2_X1 _2470_ (.A(_0615_),
    .B(\mem[3][15] ),
    .S(_0711_),
    .Z(_0300_));
 MUX2_X1 _2471_ (.A(_0617_),
    .B(\mem[3][16] ),
    .S(_0711_),
    .Z(_0301_));
 MUX2_X1 _2472_ (.A(_0619_),
    .B(\mem[3][17] ),
    .S(_0711_),
    .Z(_0302_));
 MUX2_X1 _2473_ (.A(_0621_),
    .B(\mem[3][18] ),
    .S(_0711_),
    .Z(_0303_));
 BUF_X4 _2474_ (.A(_0710_),
    .Z(_0712_));
 MUX2_X1 _2475_ (.A(_0623_),
    .B(\mem[3][19] ),
    .S(_0712_),
    .Z(_0304_));
 MUX2_X1 _2476_ (.A(_0626_),
    .B(\mem[3][1] ),
    .S(_0712_),
    .Z(_0305_));
 MUX2_X1 _2477_ (.A(_0628_),
    .B(\mem[3][20] ),
    .S(_0712_),
    .Z(_0306_));
 MUX2_X1 _2478_ (.A(_0630_),
    .B(\mem[3][21] ),
    .S(_0712_),
    .Z(_0307_));
 MUX2_X1 _2479_ (.A(_0632_),
    .B(\mem[3][22] ),
    .S(_0712_),
    .Z(_0308_));
 MUX2_X1 _2480_ (.A(_0634_),
    .B(\mem[3][23] ),
    .S(_0712_),
    .Z(_0309_));
 MUX2_X1 _2481_ (.A(_0636_),
    .B(\mem[3][24] ),
    .S(_0712_),
    .Z(_0310_));
 MUX2_X1 _2482_ (.A(_0638_),
    .B(\mem[3][25] ),
    .S(_0712_),
    .Z(_0311_));
 MUX2_X1 _2483_ (.A(_0640_),
    .B(\mem[3][26] ),
    .S(_0712_),
    .Z(_0312_));
 MUX2_X1 _2484_ (.A(_0642_),
    .B(\mem[3][27] ),
    .S(_0712_),
    .Z(_0313_));
 BUF_X4 _2485_ (.A(_0710_),
    .Z(_0713_));
 MUX2_X1 _2486_ (.A(_0644_),
    .B(\mem[3][28] ),
    .S(_0713_),
    .Z(_0314_));
 MUX2_X1 _2487_ (.A(_0647_),
    .B(\mem[3][29] ),
    .S(_0713_),
    .Z(_0315_));
 MUX2_X1 _2488_ (.A(_0649_),
    .B(\mem[3][2] ),
    .S(_0713_),
    .Z(_0316_));
 MUX2_X1 _2489_ (.A(_0651_),
    .B(\mem[3][30] ),
    .S(_0713_),
    .Z(_0317_));
 MUX2_X1 _2490_ (.A(_0653_),
    .B(\mem[3][31] ),
    .S(_0713_),
    .Z(_0318_));
 MUX2_X1 _2491_ (.A(_0655_),
    .B(\mem[3][3] ),
    .S(_0713_),
    .Z(_0319_));
 MUX2_X1 _2492_ (.A(_0657_),
    .B(\mem[3][4] ),
    .S(_0713_),
    .Z(_0320_));
 MUX2_X1 _2493_ (.A(_0659_),
    .B(\mem[3][5] ),
    .S(_0713_),
    .Z(_0321_));
 MUX2_X1 _2494_ (.A(_0661_),
    .B(\mem[3][6] ),
    .S(_0713_),
    .Z(_0322_));
 MUX2_X1 _2495_ (.A(_0663_),
    .B(\mem[3][7] ),
    .S(_0713_),
    .Z(_0323_));
 MUX2_X1 _2496_ (.A(_0665_),
    .B(\mem[3][8] ),
    .S(_0710_),
    .Z(_0324_));
 MUX2_X1 _2497_ (.A(_0667_),
    .B(\mem[3][9] ),
    .S(_0710_),
    .Z(_0325_));
 NAND3_X4 _2498_ (.A1(_1994_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0714_));
 OR2_X1 _2499_ (.A1(\wr_ptr_bin[3] ),
    .A2(_0669_),
    .ZN(_0715_));
 BUF_X4 _2500_ (.A(_0715_),
    .Z(_0716_));
 NOR2_X4 _2501_ (.A1(_0714_),
    .A2(_0716_),
    .ZN(_0717_));
 BUF_X4 _2502_ (.A(_0717_),
    .Z(_0718_));
 MUX2_X1 _2503_ (.A(\mem[4][0] ),
    .B(_0598_),
    .S(_0718_),
    .Z(_0326_));
 MUX2_X1 _2504_ (.A(\mem[4][10] ),
    .B(_0606_),
    .S(_0718_),
    .Z(_0327_));
 MUX2_X1 _2505_ (.A(\mem[4][11] ),
    .B(_0608_),
    .S(_0718_),
    .Z(_0328_));
 MUX2_X1 _2506_ (.A(\mem[4][12] ),
    .B(_0610_),
    .S(_0718_),
    .Z(_0329_));
 MUX2_X1 _2507_ (.A(\mem[4][13] ),
    .B(_0612_),
    .S(_0718_),
    .Z(_0330_));
 MUX2_X1 _2508_ (.A(\mem[4][14] ),
    .B(_0614_),
    .S(_0718_),
    .Z(_0331_));
 MUX2_X1 _2509_ (.A(\mem[4][15] ),
    .B(_0616_),
    .S(_0718_),
    .Z(_0332_));
 MUX2_X1 _2510_ (.A(\mem[4][16] ),
    .B(_0618_),
    .S(_0718_),
    .Z(_0333_));
 MUX2_X1 _2511_ (.A(\mem[4][17] ),
    .B(_0620_),
    .S(_0718_),
    .Z(_0334_));
 MUX2_X1 _2512_ (.A(\mem[4][18] ),
    .B(_0622_),
    .S(_0718_),
    .Z(_0335_));
 BUF_X4 _2513_ (.A(_0717_),
    .Z(_0719_));
 MUX2_X1 _2514_ (.A(\mem[4][19] ),
    .B(_0624_),
    .S(_0719_),
    .Z(_0336_));
 MUX2_X1 _2515_ (.A(\mem[4][1] ),
    .B(_0627_),
    .S(_0719_),
    .Z(_0337_));
 MUX2_X1 _2516_ (.A(\mem[4][20] ),
    .B(_0629_),
    .S(_0719_),
    .Z(_0338_));
 MUX2_X1 _2517_ (.A(\mem[4][21] ),
    .B(_0631_),
    .S(_0719_),
    .Z(_0339_));
 MUX2_X1 _2518_ (.A(\mem[4][22] ),
    .B(_0633_),
    .S(_0719_),
    .Z(_0340_));
 MUX2_X1 _2519_ (.A(\mem[4][23] ),
    .B(_0635_),
    .S(_0719_),
    .Z(_0341_));
 MUX2_X1 _2520_ (.A(\mem[4][24] ),
    .B(_0637_),
    .S(_0719_),
    .Z(_0342_));
 MUX2_X1 _2521_ (.A(\mem[4][25] ),
    .B(_0639_),
    .S(_0719_),
    .Z(_0343_));
 MUX2_X1 _2522_ (.A(\mem[4][26] ),
    .B(_0641_),
    .S(_0719_),
    .Z(_0344_));
 MUX2_X1 _2523_ (.A(\mem[4][27] ),
    .B(_0643_),
    .S(_0719_),
    .Z(_0345_));
 BUF_X4 _2524_ (.A(_0717_),
    .Z(_0720_));
 MUX2_X1 _2525_ (.A(\mem[4][28] ),
    .B(_0645_),
    .S(_0720_),
    .Z(_0346_));
 MUX2_X1 _2526_ (.A(\mem[4][29] ),
    .B(_0648_),
    .S(_0720_),
    .Z(_0347_));
 MUX2_X1 _2527_ (.A(\mem[4][2] ),
    .B(_0650_),
    .S(_0720_),
    .Z(_0348_));
 MUX2_X1 _2528_ (.A(\mem[4][30] ),
    .B(_0652_),
    .S(_0720_),
    .Z(_0349_));
 MUX2_X1 _2529_ (.A(\mem[4][31] ),
    .B(_0654_),
    .S(_0720_),
    .Z(_0350_));
 MUX2_X1 _2530_ (.A(\mem[4][3] ),
    .B(_0656_),
    .S(_0720_),
    .Z(_0351_));
 MUX2_X1 _2531_ (.A(\mem[4][4] ),
    .B(_0658_),
    .S(_0720_),
    .Z(_0352_));
 MUX2_X1 _2532_ (.A(\mem[4][5] ),
    .B(_0660_),
    .S(_0720_),
    .Z(_0353_));
 MUX2_X1 _2533_ (.A(\mem[4][6] ),
    .B(_0662_),
    .S(_0720_),
    .Z(_0354_));
 MUX2_X1 _2534_ (.A(\mem[4][7] ),
    .B(_0664_),
    .S(_0720_),
    .Z(_0355_));
 MUX2_X1 _2535_ (.A(\mem[4][8] ),
    .B(_0666_),
    .S(_0717_),
    .Z(_0356_));
 MUX2_X1 _2536_ (.A(\mem[4][9] ),
    .B(_0668_),
    .S(_0717_),
    .Z(_0357_));
 NAND3_X4 _2537_ (.A1(_1997_),
    .A2(_0572_),
    .A3(_0601_),
    .ZN(_0721_));
 NOR2_X4 _2538_ (.A1(_0721_),
    .A2(_0716_),
    .ZN(_0722_));
 BUF_X4 _2539_ (.A(_0722_),
    .Z(_0723_));
 MUX2_X1 _2540_ (.A(\mem[5][0] ),
    .B(_0598_),
    .S(_0723_),
    .Z(_0358_));
 MUX2_X1 _2541_ (.A(\mem[5][10] ),
    .B(_0606_),
    .S(_0723_),
    .Z(_0359_));
 MUX2_X1 _2542_ (.A(\mem[5][11] ),
    .B(_0608_),
    .S(_0723_),
    .Z(_0360_));
 MUX2_X1 _2543_ (.A(\mem[5][12] ),
    .B(_0610_),
    .S(_0723_),
    .Z(_0361_));
 MUX2_X1 _2544_ (.A(\mem[5][13] ),
    .B(_0612_),
    .S(_0723_),
    .Z(_0362_));
 MUX2_X1 _2545_ (.A(\mem[5][14] ),
    .B(_0614_),
    .S(_0723_),
    .Z(_0363_));
 MUX2_X1 _2546_ (.A(\mem[5][15] ),
    .B(_0616_),
    .S(_0723_),
    .Z(_0364_));
 MUX2_X1 _2547_ (.A(\mem[5][16] ),
    .B(_0618_),
    .S(_0723_),
    .Z(_0365_));
 MUX2_X1 _2548_ (.A(\mem[5][17] ),
    .B(_0620_),
    .S(_0723_),
    .Z(_0366_));
 MUX2_X1 _2549_ (.A(\mem[5][18] ),
    .B(_0622_),
    .S(_0723_),
    .Z(_0367_));
 BUF_X4 _2550_ (.A(_0722_),
    .Z(_0724_));
 MUX2_X1 _2551_ (.A(\mem[5][19] ),
    .B(_0624_),
    .S(_0724_),
    .Z(_0368_));
 MUX2_X1 _2552_ (.A(\mem[5][1] ),
    .B(_0627_),
    .S(_0724_),
    .Z(_0369_));
 MUX2_X1 _2553_ (.A(\mem[5][20] ),
    .B(_0629_),
    .S(_0724_),
    .Z(_0370_));
 MUX2_X1 _2554_ (.A(\mem[5][21] ),
    .B(_0631_),
    .S(_0724_),
    .Z(_0371_));
 MUX2_X1 _2555_ (.A(\mem[5][22] ),
    .B(_0633_),
    .S(_0724_),
    .Z(_0372_));
 MUX2_X1 _2556_ (.A(\mem[5][23] ),
    .B(_0635_),
    .S(_0724_),
    .Z(_0373_));
 MUX2_X1 _2557_ (.A(\mem[5][24] ),
    .B(_0637_),
    .S(_0724_),
    .Z(_0374_));
 MUX2_X1 _2558_ (.A(\mem[5][25] ),
    .B(_0639_),
    .S(_0724_),
    .Z(_0375_));
 MUX2_X1 _2559_ (.A(\mem[5][26] ),
    .B(_0641_),
    .S(_0724_),
    .Z(_0376_));
 MUX2_X1 _2560_ (.A(\mem[5][27] ),
    .B(_0643_),
    .S(_0724_),
    .Z(_0377_));
 BUF_X4 _2561_ (.A(_0722_),
    .Z(_0725_));
 MUX2_X1 _2562_ (.A(\mem[5][28] ),
    .B(_0645_),
    .S(_0725_),
    .Z(_0378_));
 MUX2_X1 _2563_ (.A(\mem[5][29] ),
    .B(_0648_),
    .S(_0725_),
    .Z(_0379_));
 MUX2_X1 _2564_ (.A(\mem[5][2] ),
    .B(_0650_),
    .S(_0725_),
    .Z(_0380_));
 MUX2_X1 _2565_ (.A(\mem[5][30] ),
    .B(_0652_),
    .S(_0725_),
    .Z(_0381_));
 MUX2_X1 _2566_ (.A(\mem[5][31] ),
    .B(_0654_),
    .S(_0725_),
    .Z(_0382_));
 MUX2_X1 _2567_ (.A(\mem[5][3] ),
    .B(_0656_),
    .S(_0725_),
    .Z(_0383_));
 MUX2_X1 _2568_ (.A(\mem[5][4] ),
    .B(_0658_),
    .S(_0725_),
    .Z(_0384_));
 MUX2_X1 _2569_ (.A(\mem[5][5] ),
    .B(_0660_),
    .S(_0725_),
    .Z(_0385_));
 MUX2_X1 _2570_ (.A(\mem[5][6] ),
    .B(_0662_),
    .S(_0725_),
    .Z(_0386_));
 MUX2_X1 _2571_ (.A(\mem[5][7] ),
    .B(_0664_),
    .S(_0725_),
    .Z(_0387_));
 MUX2_X1 _2572_ (.A(\mem[5][8] ),
    .B(_0666_),
    .S(_0722_),
    .Z(_0388_));
 MUX2_X1 _2573_ (.A(\mem[5][9] ),
    .B(_0668_),
    .S(_0722_),
    .Z(_0389_));
 NOR2_X4 _2574_ (.A1(_0671_),
    .A2(_0716_),
    .ZN(_0726_));
 BUF_X4 _2575_ (.A(_0726_),
    .Z(_0727_));
 MUX2_X1 _2576_ (.A(\mem[6][0] ),
    .B(_0598_),
    .S(_0727_),
    .Z(_0390_));
 MUX2_X1 _2577_ (.A(\mem[6][10] ),
    .B(_0606_),
    .S(_0727_),
    .Z(_0391_));
 MUX2_X1 _2578_ (.A(\mem[6][11] ),
    .B(_0608_),
    .S(_0727_),
    .Z(_0392_));
 MUX2_X1 _2579_ (.A(\mem[6][12] ),
    .B(_0610_),
    .S(_0727_),
    .Z(_0393_));
 MUX2_X1 _2580_ (.A(\mem[6][13] ),
    .B(_0612_),
    .S(_0727_),
    .Z(_0394_));
 MUX2_X1 _2581_ (.A(\mem[6][14] ),
    .B(_0614_),
    .S(_0727_),
    .Z(_0395_));
 MUX2_X1 _2582_ (.A(\mem[6][15] ),
    .B(_0616_),
    .S(_0727_),
    .Z(_0396_));
 MUX2_X1 _2583_ (.A(\mem[6][16] ),
    .B(_0618_),
    .S(_0727_),
    .Z(_0397_));
 MUX2_X1 _2584_ (.A(\mem[6][17] ),
    .B(_0620_),
    .S(_0727_),
    .Z(_0398_));
 MUX2_X1 _2585_ (.A(\mem[6][18] ),
    .B(_0622_),
    .S(_0727_),
    .Z(_0399_));
 BUF_X4 _2586_ (.A(_0726_),
    .Z(_0728_));
 MUX2_X1 _2587_ (.A(\mem[6][19] ),
    .B(_0624_),
    .S(_0728_),
    .Z(_0400_));
 MUX2_X1 _2588_ (.A(\mem[6][1] ),
    .B(_0627_),
    .S(_0728_),
    .Z(_0401_));
 MUX2_X1 _2589_ (.A(\mem[6][20] ),
    .B(_0629_),
    .S(_0728_),
    .Z(_0402_));
 MUX2_X1 _2590_ (.A(\mem[6][21] ),
    .B(_0631_),
    .S(_0728_),
    .Z(_0403_));
 MUX2_X1 _2591_ (.A(\mem[6][22] ),
    .B(_0633_),
    .S(_0728_),
    .Z(_0404_));
 MUX2_X1 _2592_ (.A(\mem[6][23] ),
    .B(_0635_),
    .S(_0728_),
    .Z(_0405_));
 MUX2_X1 _2593_ (.A(\mem[6][24] ),
    .B(_0637_),
    .S(_0728_),
    .Z(_0406_));
 MUX2_X1 _2594_ (.A(\mem[6][25] ),
    .B(_0639_),
    .S(_0728_),
    .Z(_0407_));
 MUX2_X1 _2595_ (.A(\mem[6][26] ),
    .B(_0641_),
    .S(_0728_),
    .Z(_0408_));
 MUX2_X1 _2596_ (.A(\mem[6][27] ),
    .B(_0643_),
    .S(_0728_),
    .Z(_0409_));
 BUF_X4 _2597_ (.A(_0726_),
    .Z(_0729_));
 MUX2_X1 _2598_ (.A(\mem[6][28] ),
    .B(_0645_),
    .S(_0729_),
    .Z(_0410_));
 MUX2_X1 _2599_ (.A(\mem[6][29] ),
    .B(_0648_),
    .S(_0729_),
    .Z(_0411_));
 MUX2_X1 _2600_ (.A(\mem[6][2] ),
    .B(_0650_),
    .S(_0729_),
    .Z(_0412_));
 MUX2_X1 _2601_ (.A(\mem[6][30] ),
    .B(_0652_),
    .S(_0729_),
    .Z(_0413_));
 MUX2_X1 _2602_ (.A(\mem[6][31] ),
    .B(_0654_),
    .S(_0729_),
    .Z(_0414_));
 MUX2_X1 _2603_ (.A(\mem[6][3] ),
    .B(_0656_),
    .S(_0729_),
    .Z(_0415_));
 MUX2_X1 _2604_ (.A(\mem[6][4] ),
    .B(_0658_),
    .S(_0729_),
    .Z(_0416_));
 MUX2_X1 _2605_ (.A(\mem[6][5] ),
    .B(_0660_),
    .S(_0729_),
    .Z(_0417_));
 MUX2_X1 _2606_ (.A(\mem[6][6] ),
    .B(_0662_),
    .S(_0729_),
    .Z(_0418_));
 MUX2_X1 _2607_ (.A(\mem[6][7] ),
    .B(_0664_),
    .S(_0729_),
    .Z(_0419_));
 MUX2_X1 _2608_ (.A(\mem[6][8] ),
    .B(_0666_),
    .S(_0726_),
    .Z(_0420_));
 MUX2_X1 _2609_ (.A(\mem[6][9] ),
    .B(_0668_),
    .S(_0726_),
    .Z(_0421_));
 NOR2_X4 _2610_ (.A1(_0676_),
    .A2(_0716_),
    .ZN(_0730_));
 BUF_X4 _2611_ (.A(_0730_),
    .Z(_0731_));
 MUX2_X1 _2612_ (.A(\mem[7][0] ),
    .B(_0598_),
    .S(_0731_),
    .Z(_0422_));
 MUX2_X1 _2613_ (.A(\mem[7][10] ),
    .B(_0606_),
    .S(_0731_),
    .Z(_0423_));
 MUX2_X1 _2614_ (.A(\mem[7][11] ),
    .B(_0608_),
    .S(_0731_),
    .Z(_0424_));
 MUX2_X1 _2615_ (.A(\mem[7][12] ),
    .B(_0610_),
    .S(_0731_),
    .Z(_0425_));
 MUX2_X1 _2616_ (.A(\mem[7][13] ),
    .B(_0612_),
    .S(_0731_),
    .Z(_0426_));
 MUX2_X1 _2617_ (.A(\mem[7][14] ),
    .B(_0614_),
    .S(_0731_),
    .Z(_0427_));
 MUX2_X1 _2618_ (.A(\mem[7][15] ),
    .B(_0616_),
    .S(_0731_),
    .Z(_0428_));
 MUX2_X1 _2619_ (.A(\mem[7][16] ),
    .B(_0618_),
    .S(_0731_),
    .Z(_0429_));
 MUX2_X1 _2620_ (.A(\mem[7][17] ),
    .B(_0620_),
    .S(_0731_),
    .Z(_0430_));
 MUX2_X1 _2621_ (.A(\mem[7][18] ),
    .B(_0622_),
    .S(_0731_),
    .Z(_0431_));
 BUF_X4 _2622_ (.A(_0730_),
    .Z(_0732_));
 MUX2_X1 _2623_ (.A(\mem[7][19] ),
    .B(_0624_),
    .S(_0732_),
    .Z(_0432_));
 MUX2_X1 _2624_ (.A(\mem[7][1] ),
    .B(_0627_),
    .S(_0732_),
    .Z(_0433_));
 MUX2_X1 _2625_ (.A(\mem[7][20] ),
    .B(_0629_),
    .S(_0732_),
    .Z(_0434_));
 MUX2_X1 _2626_ (.A(\mem[7][21] ),
    .B(_0631_),
    .S(_0732_),
    .Z(_0435_));
 MUX2_X1 _2627_ (.A(\mem[7][22] ),
    .B(_0633_),
    .S(_0732_),
    .Z(_0436_));
 MUX2_X1 _2628_ (.A(\mem[7][23] ),
    .B(_0635_),
    .S(_0732_),
    .Z(_0437_));
 MUX2_X1 _2629_ (.A(\mem[7][24] ),
    .B(_0637_),
    .S(_0732_),
    .Z(_0438_));
 MUX2_X1 _2630_ (.A(\mem[7][25] ),
    .B(_0639_),
    .S(_0732_),
    .Z(_0439_));
 MUX2_X1 _2631_ (.A(\mem[7][26] ),
    .B(_0641_),
    .S(_0732_),
    .Z(_0440_));
 MUX2_X1 _2632_ (.A(\mem[7][27] ),
    .B(_0643_),
    .S(_0732_),
    .Z(_0441_));
 BUF_X4 _2633_ (.A(_0730_),
    .Z(_0733_));
 MUX2_X1 _2634_ (.A(\mem[7][28] ),
    .B(_0645_),
    .S(_0733_),
    .Z(_0442_));
 MUX2_X1 _2635_ (.A(\mem[7][29] ),
    .B(_0648_),
    .S(_0733_),
    .Z(_0443_));
 MUX2_X1 _2636_ (.A(\mem[7][2] ),
    .B(_0650_),
    .S(_0733_),
    .Z(_0444_));
 MUX2_X1 _2637_ (.A(\mem[7][30] ),
    .B(_0652_),
    .S(_0733_),
    .Z(_0445_));
 MUX2_X1 _2638_ (.A(\mem[7][31] ),
    .B(_0654_),
    .S(_0733_),
    .Z(_0446_));
 MUX2_X1 _2639_ (.A(\mem[7][3] ),
    .B(_0656_),
    .S(_0733_),
    .Z(_0447_));
 MUX2_X1 _2640_ (.A(\mem[7][4] ),
    .B(_0658_),
    .S(_0733_),
    .Z(_0448_));
 MUX2_X1 _2641_ (.A(\mem[7][5] ),
    .B(_0660_),
    .S(_0733_),
    .Z(_0449_));
 MUX2_X1 _2642_ (.A(\mem[7][6] ),
    .B(_0662_),
    .S(_0733_),
    .Z(_0450_));
 MUX2_X1 _2643_ (.A(\mem[7][7] ),
    .B(_0664_),
    .S(_0733_),
    .Z(_0451_));
 MUX2_X1 _2644_ (.A(\mem[7][8] ),
    .B(_0666_),
    .S(_0730_),
    .Z(_0452_));
 MUX2_X1 _2645_ (.A(\mem[7][9] ),
    .B(_0668_),
    .S(_0730_),
    .Z(_0453_));
 NOR2_X4 _2646_ (.A1(_0714_),
    .A2(_0670_),
    .ZN(_0734_));
 BUF_X4 _2647_ (.A(_0734_),
    .Z(_0735_));
 MUX2_X1 _2648_ (.A(\mem[8][0] ),
    .B(_0598_),
    .S(_0735_),
    .Z(_0454_));
 MUX2_X1 _2649_ (.A(\mem[8][10] ),
    .B(_0606_),
    .S(_0735_),
    .Z(_0455_));
 MUX2_X1 _2650_ (.A(\mem[8][11] ),
    .B(_0608_),
    .S(_0735_),
    .Z(_0456_));
 MUX2_X1 _2651_ (.A(\mem[8][12] ),
    .B(_0610_),
    .S(_0735_),
    .Z(_0457_));
 MUX2_X1 _2652_ (.A(\mem[8][13] ),
    .B(_0612_),
    .S(_0735_),
    .Z(_0458_));
 MUX2_X1 _2653_ (.A(\mem[8][14] ),
    .B(_0614_),
    .S(_0735_),
    .Z(_0459_));
 MUX2_X1 _2654_ (.A(\mem[8][15] ),
    .B(_0616_),
    .S(_0735_),
    .Z(_0460_));
 MUX2_X1 _2655_ (.A(\mem[8][16] ),
    .B(_0618_),
    .S(_0735_),
    .Z(_0461_));
 MUX2_X1 _2656_ (.A(\mem[8][17] ),
    .B(_0620_),
    .S(_0735_),
    .Z(_0462_));
 MUX2_X1 _2657_ (.A(\mem[8][18] ),
    .B(_0622_),
    .S(_0735_),
    .Z(_0463_));
 BUF_X4 _2658_ (.A(_0734_),
    .Z(_0736_));
 MUX2_X1 _2659_ (.A(\mem[8][19] ),
    .B(_0624_),
    .S(_0736_),
    .Z(_0464_));
 MUX2_X1 _2660_ (.A(\mem[8][1] ),
    .B(_0627_),
    .S(_0736_),
    .Z(_0465_));
 MUX2_X1 _2661_ (.A(\mem[8][20] ),
    .B(_0629_),
    .S(_0736_),
    .Z(_0466_));
 MUX2_X1 _2662_ (.A(\mem[8][21] ),
    .B(_0631_),
    .S(_0736_),
    .Z(_0467_));
 MUX2_X1 _2663_ (.A(\mem[8][22] ),
    .B(_0633_),
    .S(_0736_),
    .Z(_0468_));
 MUX2_X1 _2664_ (.A(\mem[8][23] ),
    .B(_0635_),
    .S(_0736_),
    .Z(_0469_));
 MUX2_X1 _2665_ (.A(\mem[8][24] ),
    .B(_0637_),
    .S(_0736_),
    .Z(_0470_));
 MUX2_X1 _2666_ (.A(\mem[8][25] ),
    .B(_0639_),
    .S(_0736_),
    .Z(_0471_));
 MUX2_X1 _2667_ (.A(\mem[8][26] ),
    .B(_0641_),
    .S(_0736_),
    .Z(_0472_));
 MUX2_X1 _2668_ (.A(\mem[8][27] ),
    .B(_0643_),
    .S(_0736_),
    .Z(_0473_));
 BUF_X4 _2669_ (.A(_0734_),
    .Z(_0737_));
 MUX2_X1 _2670_ (.A(\mem[8][28] ),
    .B(_0645_),
    .S(_0737_),
    .Z(_0474_));
 MUX2_X1 _2671_ (.A(\mem[8][29] ),
    .B(_0648_),
    .S(_0737_),
    .Z(_0475_));
 MUX2_X1 _2672_ (.A(\mem[8][2] ),
    .B(_0650_),
    .S(_0737_),
    .Z(_0476_));
 MUX2_X1 _2673_ (.A(\mem[8][30] ),
    .B(_0652_),
    .S(_0737_),
    .Z(_0477_));
 MUX2_X1 _2674_ (.A(\mem[8][31] ),
    .B(_0654_),
    .S(_0737_),
    .Z(_0478_));
 MUX2_X1 _2675_ (.A(\mem[8][3] ),
    .B(_0656_),
    .S(_0737_),
    .Z(_0479_));
 MUX2_X1 _2676_ (.A(\mem[8][4] ),
    .B(_0658_),
    .S(_0737_),
    .Z(_0480_));
 MUX2_X1 _2677_ (.A(\mem[8][5] ),
    .B(_0660_),
    .S(_0737_),
    .Z(_0481_));
 MUX2_X1 _2678_ (.A(\mem[8][6] ),
    .B(_0662_),
    .S(_0737_),
    .Z(_0482_));
 MUX2_X1 _2679_ (.A(\mem[8][7] ),
    .B(_0664_),
    .S(_0737_),
    .Z(_0483_));
 MUX2_X1 _2680_ (.A(\mem[8][8] ),
    .B(_0666_),
    .S(_0734_),
    .Z(_0484_));
 MUX2_X1 _2681_ (.A(\mem[8][9] ),
    .B(_0668_),
    .S(_0734_),
    .Z(_0485_));
 NOR2_X4 _2682_ (.A1(_0670_),
    .A2(_0721_),
    .ZN(_0738_));
 BUF_X4 _2683_ (.A(_0738_),
    .Z(_0739_));
 MUX2_X1 _2684_ (.A(\mem[9][0] ),
    .B(_0598_),
    .S(_0739_),
    .Z(_0486_));
 MUX2_X1 _2685_ (.A(\mem[9][10] ),
    .B(_0606_),
    .S(_0739_),
    .Z(_0487_));
 MUX2_X1 _2686_ (.A(\mem[9][11] ),
    .B(_0608_),
    .S(_0739_),
    .Z(_0488_));
 MUX2_X1 _2687_ (.A(\mem[9][12] ),
    .B(_0610_),
    .S(_0739_),
    .Z(_0489_));
 MUX2_X1 _2688_ (.A(\mem[9][13] ),
    .B(_0612_),
    .S(_0739_),
    .Z(_0490_));
 MUX2_X1 _2689_ (.A(\mem[9][14] ),
    .B(_0614_),
    .S(_0739_),
    .Z(_0491_));
 MUX2_X1 _2690_ (.A(\mem[9][15] ),
    .B(_0616_),
    .S(_0739_),
    .Z(_0492_));
 MUX2_X1 _2691_ (.A(\mem[9][16] ),
    .B(_0618_),
    .S(_0739_),
    .Z(_0493_));
 MUX2_X1 _2692_ (.A(\mem[9][17] ),
    .B(_0620_),
    .S(_0739_),
    .Z(_0494_));
 MUX2_X1 _2693_ (.A(\mem[9][18] ),
    .B(_0622_),
    .S(_0739_),
    .Z(_0495_));
 BUF_X4 _2694_ (.A(_0738_),
    .Z(_0740_));
 MUX2_X1 _2695_ (.A(\mem[9][19] ),
    .B(_0624_),
    .S(_0740_),
    .Z(_0496_));
 MUX2_X1 _2696_ (.A(\mem[9][1] ),
    .B(_0627_),
    .S(_0740_),
    .Z(_0497_));
 MUX2_X1 _2697_ (.A(\mem[9][20] ),
    .B(_0629_),
    .S(_0740_),
    .Z(_0498_));
 MUX2_X1 _2698_ (.A(\mem[9][21] ),
    .B(_0631_),
    .S(_0740_),
    .Z(_0499_));
 MUX2_X1 _2699_ (.A(\mem[9][22] ),
    .B(_0633_),
    .S(_0740_),
    .Z(_0500_));
 MUX2_X1 _2700_ (.A(\mem[9][23] ),
    .B(_0635_),
    .S(_0740_),
    .Z(_0501_));
 MUX2_X1 _2701_ (.A(\mem[9][24] ),
    .B(_0637_),
    .S(_0740_),
    .Z(_0502_));
 MUX2_X1 _2702_ (.A(\mem[9][25] ),
    .B(_0639_),
    .S(_0740_),
    .Z(_0503_));
 MUX2_X1 _2703_ (.A(\mem[9][26] ),
    .B(_0641_),
    .S(_0740_),
    .Z(_0504_));
 MUX2_X1 _2704_ (.A(\mem[9][27] ),
    .B(_0643_),
    .S(_0740_),
    .Z(_0505_));
 BUF_X4 _2705_ (.A(_0738_),
    .Z(_0741_));
 MUX2_X1 _2706_ (.A(\mem[9][28] ),
    .B(_0645_),
    .S(_0741_),
    .Z(_0506_));
 MUX2_X1 _2707_ (.A(\mem[9][29] ),
    .B(_0648_),
    .S(_0741_),
    .Z(_0507_));
 MUX2_X1 _2708_ (.A(\mem[9][2] ),
    .B(_0650_),
    .S(_0741_),
    .Z(_0508_));
 MUX2_X1 _2709_ (.A(\mem[9][30] ),
    .B(_0652_),
    .S(_0741_),
    .Z(_0509_));
 MUX2_X1 _2710_ (.A(\mem[9][31] ),
    .B(_0654_),
    .S(_0741_),
    .Z(_0510_));
 MUX2_X1 _2711_ (.A(\mem[9][3] ),
    .B(_0656_),
    .S(_0741_),
    .Z(_0511_));
 MUX2_X1 _2712_ (.A(\mem[9][4] ),
    .B(_0658_),
    .S(_0741_),
    .Z(_0512_));
 MUX2_X1 _2713_ (.A(\mem[9][5] ),
    .B(_0660_),
    .S(_0741_),
    .Z(_0513_));
 MUX2_X1 _2714_ (.A(\mem[9][6] ),
    .B(_0662_),
    .S(_0741_),
    .Z(_0514_));
 MUX2_X1 _2715_ (.A(\mem[9][7] ),
    .B(_0664_),
    .S(_0741_),
    .Z(_0515_));
 MUX2_X1 _2716_ (.A(\mem[9][8] ),
    .B(_0666_),
    .S(_0738_),
    .Z(_0516_));
 MUX2_X1 _2717_ (.A(\mem[9][9] ),
    .B(_0668_),
    .S(_0738_),
    .Z(_0517_));
 OAI21_X4 _2718_ (.A(net2),
    .B1(_0591_),
    .B2(_0596_),
    .ZN(_0742_));
 BUF_X4 _2719_ (.A(_0742_),
    .Z(_0743_));
 NAND2_X1 _2720_ (.A1(net12),
    .A2(_0743_),
    .ZN(_0744_));
 BUF_X4 _2721_ (.A(_2001_),
    .Z(_0745_));
 BUF_X4 _2722_ (.A(_0745_),
    .Z(_0746_));
 INV_X2 _2723_ (.A(_0746_),
    .ZN(_0747_));
 BUF_X4 _2724_ (.A(\rd_ptr_bin[3] ),
    .Z(_0748_));
 BUF_X4 _2725_ (.A(\rd_ptr_bin[2] ),
    .Z(_0749_));
 NOR2_X4 _2726_ (.A1(_0748_),
    .A2(_0749_),
    .ZN(_0750_));
 NOR2_X2 _2727_ (.A1(_0747_),
    .A2(_0750_),
    .ZN(_0751_));
 BUF_X4 _2728_ (.A(_0751_),
    .Z(_0752_));
 BUF_X2 _2729_ (.A(_2006_),
    .Z(_0753_));
 BUF_X4 _2730_ (.A(_0753_),
    .Z(_0754_));
 BUF_X4 _2731_ (.A(_0754_),
    .Z(_0755_));
 BUF_X4 _2732_ (.A(_2002_),
    .Z(_0756_));
 BUF_X4 _2733_ (.A(_0756_),
    .Z(_0757_));
 BUF_X4 _2734_ (.A(_0757_),
    .Z(_0758_));
 CLKBUF_X3 _2735_ (.A(_2004_),
    .Z(_0759_));
 BUF_X4 _2736_ (.A(_0759_),
    .Z(_0760_));
 BUF_X4 _2737_ (.A(_0760_),
    .Z(_0761_));
 OR3_X2 _2738_ (.A1(_0755_),
    .A2(_0758_),
    .A3(_0761_),
    .ZN(_0762_));
 BUF_X4 _2739_ (.A(_0762_),
    .Z(_0763_));
 BUF_X4 _2740_ (.A(_0754_),
    .Z(_0764_));
 BUF_X4 _2741_ (.A(_0764_),
    .Z(_0765_));
 AND2_X1 _2742_ (.A1(_0748_),
    .A2(_0749_),
    .ZN(_0766_));
 BUF_X4 _2743_ (.A(_0766_),
    .Z(_0767_));
 BUF_X4 _2744_ (.A(_0767_),
    .Z(_0768_));
 NAND3_X1 _2745_ (.A1(_0765_),
    .A2(\mem[15][0] ),
    .A3(_0768_),
    .ZN(_0769_));
 NOR3_X2 _2746_ (.A1(_0753_),
    .A2(_0757_),
    .A3(_0760_),
    .ZN(_0770_));
 OAI21_X4 _2747_ (.A(_0770_),
    .B1(_0750_),
    .B2(_0747_),
    .ZN(_0771_));
 BUF_X4 _2748_ (.A(_0771_),
    .Z(_0772_));
 INV_X2 _2749_ (.A(_0748_),
    .ZN(_0773_));
 BUF_X4 _2750_ (.A(_0773_),
    .Z(_0774_));
 BUF_X4 _2751_ (.A(_0774_),
    .Z(_0775_));
 BUF_X4 _2752_ (.A(_0749_),
    .Z(_0776_));
 BUF_X4 _2753_ (.A(_0776_),
    .Z(_0777_));
 BUF_X4 _2754_ (.A(_0757_),
    .Z(_0778_));
 BUF_X4 _2755_ (.A(_0778_),
    .Z(_0779_));
 NAND4_X1 _2756_ (.A1(_0775_),
    .A2(_0777_),
    .A3(\mem[6][0] ),
    .A4(_0779_),
    .ZN(_0780_));
 BUF_X4 _2757_ (.A(_0748_),
    .Z(_0781_));
 BUF_X4 _2758_ (.A(_0781_),
    .Z(_0782_));
 INV_X4 _2759_ (.A(_0749_),
    .ZN(_0783_));
 BUF_X4 _2760_ (.A(_0783_),
    .Z(_0784_));
 BUF_X4 _2761_ (.A(_0759_),
    .Z(_0785_));
 BUF_X4 _2762_ (.A(_0785_),
    .Z(_0786_));
 BUF_X4 _2763_ (.A(_0786_),
    .Z(_0787_));
 NAND4_X1 _2764_ (.A1(_0782_),
    .A2(_0784_),
    .A3(\mem[9][0] ),
    .A4(_0787_),
    .ZN(_0788_));
 NAND4_X1 _2765_ (.A1(_0769_),
    .A2(_0772_),
    .A3(_0780_),
    .A4(_0788_),
    .ZN(_0789_));
 AOI222_X2 _2766_ (.A1(_0754_),
    .A2(\mem[3][0] ),
    .B1(\mem[2][0] ),
    .B2(_0757_),
    .C1(_0759_),
    .C2(\mem[1][0] ),
    .ZN(_0790_));
 OR3_X1 _2767_ (.A1(_0781_),
    .A2(_0776_),
    .A3(_0790_),
    .ZN(_0791_));
 BUF_X4 _2768_ (.A(_0749_),
    .Z(_0792_));
 BUF_X4 _2769_ (.A(_0757_),
    .Z(_0793_));
 AOI221_X1 _2770_ (.A(_0792_),
    .B1(\mem[8][0] ),
    .B2(_0746_),
    .C1(_0793_),
    .C2(\mem[10][0] ),
    .ZN(_0794_));
 BUF_X4 _2771_ (.A(_0783_),
    .Z(_0795_));
 AND2_X1 _2772_ (.A1(\mem[14][0] ),
    .A2(_0793_),
    .ZN(_0796_));
 OAI21_X1 _2773_ (.A(_0781_),
    .B1(_0795_),
    .B2(_0796_),
    .ZN(_0797_));
 MUX2_X1 _2774_ (.A(\mem[5][0] ),
    .B(\mem[13][0] ),
    .S(_0781_),
    .Z(_0798_));
 MUX2_X1 _2775_ (.A(\mem[4][0] ),
    .B(\mem[12][0] ),
    .S(_0781_),
    .Z(_0799_));
 BUF_X4 _2776_ (.A(_0745_),
    .Z(_0800_));
 BUF_X4 _2777_ (.A(_0800_),
    .Z(_0801_));
 AOI22_X1 _2778_ (.A1(_0786_),
    .A2(_0798_),
    .B1(_0799_),
    .B2(_0801_),
    .ZN(_0802_));
 OAI221_X1 _2779_ (.A(_0791_),
    .B1(_0794_),
    .B2(_0797_),
    .C1(_0802_),
    .C2(_0784_),
    .ZN(_0803_));
 BUF_X4 _2780_ (.A(_0754_),
    .Z(_0804_));
 INV_X4 _2781_ (.A(_0804_),
    .ZN(_0805_));
 NAND3_X1 _2782_ (.A1(_0775_),
    .A2(_0777_),
    .A3(\mem[7][0] ),
    .ZN(_0806_));
 NAND3_X1 _2783_ (.A1(_0782_),
    .A2(_0784_),
    .A3(\mem[11][0] ),
    .ZN(_0807_));
 AOI21_X1 _2784_ (.A(_0805_),
    .B1(_0806_),
    .B2(_0807_),
    .ZN(_0808_));
 OAI33_X1 _2785_ (.A1(\mem[0][0] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0789_),
    .B2(_0803_),
    .B3(_0808_),
    .ZN(_0809_));
 CLKBUF_X3 _2786_ (.A(_0742_),
    .Z(_0810_));
 OAI21_X1 _2787_ (.A(_0744_),
    .B1(_0809_),
    .B2(_0810_),
    .ZN(_0518_));
 NAND2_X1 _2788_ (.A1(net13),
    .A2(_0743_),
    .ZN(_0811_));
 INV_X1 _2789_ (.A(net2),
    .ZN(_0812_));
 AND4_X1 _2790_ (.A1(_0592_),
    .A2(_0593_),
    .A3(_0594_),
    .A4(_0595_),
    .ZN(_0813_));
 AOI21_X2 _2791_ (.A(_0812_),
    .B1(_0588_),
    .B2(_0813_),
    .ZN(_0814_));
 BUF_X4 _2792_ (.A(_0814_),
    .Z(_0815_));
 BUF_X4 _2793_ (.A(_0771_),
    .Z(_0816_));
 BUF_X4 _2794_ (.A(_0816_),
    .Z(_0817_));
 OAI21_X1 _2795_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][10] ),
    .ZN(_0818_));
 MUX2_X1 _2796_ (.A(\mem[7][10] ),
    .B(\mem[15][10] ),
    .S(_0748_),
    .Z(_0819_));
 NAND3_X1 _2797_ (.A1(_0777_),
    .A2(_0804_),
    .A3(_0819_),
    .ZN(_0820_));
 NAND2_X1 _2798_ (.A1(_0771_),
    .A2(_0820_),
    .ZN(_0821_));
 AOI221_X2 _2799_ (.A(_0749_),
    .B1(\mem[10][10] ),
    .B2(_0756_),
    .C1(_0785_),
    .C2(\mem[9][10] ),
    .ZN(_0822_));
 BUF_X4 _2800_ (.A(_0757_),
    .Z(_0823_));
 AOI22_X1 _2801_ (.A1(\mem[12][10] ),
    .A2(_0801_),
    .B1(_0823_),
    .B2(\mem[14][10] ),
    .ZN(_0824_));
 AOI21_X1 _2802_ (.A(_0822_),
    .B1(_0824_),
    .B2(_0777_),
    .ZN(_0825_));
 INV_X1 _2803_ (.A(_0786_),
    .ZN(_0826_));
 MUX2_X1 _2804_ (.A(\mem[5][10] ),
    .B(\mem[13][10] ),
    .S(_0748_),
    .Z(_0827_));
 INV_X1 _2805_ (.A(_0827_),
    .ZN(_0828_));
 AOI22_X1 _2806_ (.A1(\mem[4][10] ),
    .A2(_0801_),
    .B1(_0778_),
    .B2(\mem[6][10] ),
    .ZN(_0829_));
 OAI221_X2 _2807_ (.A(_0777_),
    .B1(_0826_),
    .B2(_0828_),
    .C1(_0829_),
    .C2(_0782_),
    .ZN(_0830_));
 AOI22_X1 _2808_ (.A1(_0754_),
    .A2(\mem[11][10] ),
    .B1(\mem[8][10] ),
    .B2(_0800_),
    .ZN(_0831_));
 BUF_X4 _2809_ (.A(_0756_),
    .Z(_0832_));
 AOI22_X1 _2810_ (.A1(\mem[2][10] ),
    .A2(_0832_),
    .B1(_0785_),
    .B2(\mem[1][10] ),
    .ZN(_0833_));
 AOI21_X1 _2811_ (.A(_0748_),
    .B1(_0754_),
    .B2(\mem[3][10] ),
    .ZN(_0834_));
 AOI22_X1 _2812_ (.A1(_0781_),
    .A2(_0831_),
    .B1(_0833_),
    .B2(_0834_),
    .ZN(_0835_));
 OR2_X1 _2813_ (.A1(_0777_),
    .A2(_0835_),
    .ZN(_0836_));
 AOI221_X2 _2814_ (.A(_0821_),
    .B1(_0825_),
    .B2(_0782_),
    .C1(_0830_),
    .C2(_0836_),
    .ZN(_0837_));
 OAI21_X1 _2815_ (.A(_0811_),
    .B1(_0818_),
    .B2(_0837_),
    .ZN(_0519_));
 NAND2_X1 _2816_ (.A1(net14),
    .A2(_0743_),
    .ZN(_0838_));
 BUF_X4 _2817_ (.A(_0805_),
    .Z(_0839_));
 BUF_X4 _2818_ (.A(_0749_),
    .Z(_0840_));
 MUX2_X1 _2819_ (.A(\mem[3][11] ),
    .B(\mem[7][11] ),
    .S(_0840_),
    .Z(_0841_));
 AOI22_X1 _2820_ (.A1(\mem[15][11] ),
    .A2(_0768_),
    .B1(_0841_),
    .B2(_0775_),
    .ZN(_0842_));
 NOR2_X1 _2821_ (.A1(_0839_),
    .A2(_0842_),
    .ZN(_0843_));
 NAND2_X4 _2822_ (.A1(_0748_),
    .A2(_0749_),
    .ZN(_0844_));
 CLKBUF_X3 _2823_ (.A(_0844_),
    .Z(_0845_));
 BUF_X4 _2824_ (.A(_0800_),
    .Z(_0846_));
 AOI22_X1 _2825_ (.A1(\mem[12][11] ),
    .A2(_0846_),
    .B1(_0758_),
    .B2(\mem[14][11] ),
    .ZN(_0847_));
 OR2_X1 _2826_ (.A1(_0845_),
    .A2(_0847_),
    .ZN(_0848_));
 CLKBUF_X3 _2827_ (.A(_0750_),
    .Z(_0849_));
 NAND3_X1 _2828_ (.A1(\mem[2][11] ),
    .A2(_0779_),
    .A3(_0849_),
    .ZN(_0850_));
 AND2_X1 _2829_ (.A1(_0748_),
    .A2(_0759_),
    .ZN(_0851_));
 CLKBUF_X3 _2830_ (.A(_0851_),
    .Z(_0852_));
 CLKBUF_X3 _2831_ (.A(_0852_),
    .Z(_0853_));
 MUX2_X1 _2832_ (.A(\mem[9][11] ),
    .B(\mem[13][11] ),
    .S(_0776_),
    .Z(_0854_));
 NAND2_X1 _2833_ (.A1(_0853_),
    .A2(_0854_),
    .ZN(_0855_));
 NAND4_X1 _2834_ (.A1(_0772_),
    .A2(_0848_),
    .A3(_0850_),
    .A4(_0855_),
    .ZN(_0856_));
 NAND2_X2 _2835_ (.A1(_0781_),
    .A2(_0783_),
    .ZN(_0857_));
 BUF_X4 _2836_ (.A(_0857_),
    .Z(_0858_));
 BUF_X4 _2837_ (.A(_0754_),
    .Z(_0859_));
 AOI222_X2 _2838_ (.A1(_0859_),
    .A2(\mem[11][11] ),
    .B1(\mem[8][11] ),
    .B2(_0801_),
    .C1(_0778_),
    .C2(\mem[10][11] ),
    .ZN(_0860_));
 BUF_X4 _2839_ (.A(_0756_),
    .Z(_0861_));
 BUF_X4 _2840_ (.A(_0759_),
    .Z(_0862_));
 AOI222_X2 _2841_ (.A1(\mem[6][11] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][11] ),
    .C1(\mem[4][11] ),
    .C2(_0746_),
    .ZN(_0863_));
 NAND2_X1 _2842_ (.A1(\mem[1][11] ),
    .A2(_0761_),
    .ZN(_0864_));
 BUF_X4 _2843_ (.A(_0783_),
    .Z(_0865_));
 MUX2_X1 _2844_ (.A(_0863_),
    .B(_0864_),
    .S(_0865_),
    .Z(_0866_));
 BUF_X4 _2845_ (.A(_0781_),
    .Z(_0867_));
 OAI22_X1 _2846_ (.A1(_0858_),
    .A2(_0860_),
    .B1(_0866_),
    .B2(_0867_),
    .ZN(_0868_));
 OAI33_X1 _2847_ (.A1(\mem[0][11] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0843_),
    .B2(_0856_),
    .B3(_0868_),
    .ZN(_0869_));
 OAI21_X1 _2848_ (.A(_0838_),
    .B1(_0869_),
    .B2(_0810_),
    .ZN(_0520_));
 NAND2_X1 _2849_ (.A1(net15),
    .A2(_0743_),
    .ZN(_0870_));
 BUF_X4 _2850_ (.A(_0857_),
    .Z(_0871_));
 BUF_X4 _2851_ (.A(_0778_),
    .Z(_0872_));
 AOI22_X1 _2852_ (.A1(\mem[10][12] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][12] ),
    .ZN(_0873_));
 BUF_X4 _2853_ (.A(_0846_),
    .Z(_0874_));
 AOI22_X1 _2854_ (.A1(_0765_),
    .A2(\mem[11][12] ),
    .B1(\mem[8][12] ),
    .B2(_0874_),
    .ZN(_0875_));
 AOI21_X1 _2855_ (.A(_0871_),
    .B1(_0873_),
    .B2(_0875_),
    .ZN(_0876_));
 MUX2_X1 _2856_ (.A(\mem[7][12] ),
    .B(\mem[15][12] ),
    .S(_0781_),
    .Z(_0877_));
 NAND3_X1 _2857_ (.A1(_0777_),
    .A2(_0859_),
    .A3(_0877_),
    .ZN(_0878_));
 BUF_X4 _2858_ (.A(_0745_),
    .Z(_0879_));
 AOI222_X2 _2859_ (.A1(\mem[14][12] ),
    .A2(_0778_),
    .B1(_0786_),
    .B2(\mem[13][12] ),
    .C1(\mem[12][12] ),
    .C2(_0879_),
    .ZN(_0880_));
 OAI221_X1 _2860_ (.A(_0878_),
    .B1(_0762_),
    .B2(_0751_),
    .C1(_0845_),
    .C2(_0880_),
    .ZN(_0881_));
 AOI222_X2 _2861_ (.A1(\mem[6][12] ),
    .A2(_0793_),
    .B1(_0785_),
    .B2(\mem[5][12] ),
    .C1(\mem[4][12] ),
    .C2(_0746_),
    .ZN(_0882_));
 AOI222_X2 _2862_ (.A1(_0754_),
    .A2(\mem[3][12] ),
    .B1(\mem[2][12] ),
    .B2(_0757_),
    .C1(_0785_),
    .C2(\mem[1][12] ),
    .ZN(_0883_));
 MUX2_X1 _2863_ (.A(_0882_),
    .B(_0883_),
    .S(_0865_),
    .Z(_0884_));
 NOR2_X1 _2864_ (.A1(_0867_),
    .A2(_0884_),
    .ZN(_0885_));
 OAI33_X1 _2865_ (.A1(\mem[0][12] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0876_),
    .B2(_0881_),
    .B3(_0885_),
    .ZN(_0886_));
 OAI21_X1 _2866_ (.A(_0870_),
    .B1(_0886_),
    .B2(_0810_),
    .ZN(_0521_));
 NAND2_X1 _2867_ (.A1(net16),
    .A2(_0743_),
    .ZN(_0887_));
 MUX2_X1 _2868_ (.A(\mem[3][13] ),
    .B(\mem[7][13] ),
    .S(_0840_),
    .Z(_0888_));
 AOI22_X1 _2869_ (.A1(\mem[15][13] ),
    .A2(_0768_),
    .B1(_0888_),
    .B2(_0775_),
    .ZN(_0889_));
 NOR2_X1 _2870_ (.A1(_0839_),
    .A2(_0889_),
    .ZN(_0890_));
 BUF_X4 _2871_ (.A(_0757_),
    .Z(_0891_));
 AOI22_X1 _2872_ (.A1(\mem[12][13] ),
    .A2(_0846_),
    .B1(_0891_),
    .B2(\mem[14][13] ),
    .ZN(_0892_));
 OR2_X1 _2873_ (.A1(_0845_),
    .A2(_0892_),
    .ZN(_0893_));
 NAND3_X1 _2874_ (.A1(\mem[2][13] ),
    .A2(_0779_),
    .A3(_0849_),
    .ZN(_0894_));
 MUX2_X1 _2875_ (.A(\mem[9][13] ),
    .B(\mem[13][13] ),
    .S(_0776_),
    .Z(_0895_));
 NAND2_X1 _2876_ (.A1(_0853_),
    .A2(_0895_),
    .ZN(_0896_));
 NAND4_X1 _2877_ (.A1(_0772_),
    .A2(_0893_),
    .A3(_0894_),
    .A4(_0896_),
    .ZN(_0897_));
 AOI222_X2 _2878_ (.A1(_0859_),
    .A2(\mem[11][13] ),
    .B1(\mem[8][13] ),
    .B2(_0801_),
    .C1(_0778_),
    .C2(\mem[10][13] ),
    .ZN(_0898_));
 AOI222_X2 _2879_ (.A1(\mem[6][13] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][13] ),
    .C1(\mem[4][13] ),
    .C2(_0746_),
    .ZN(_0899_));
 NAND2_X1 _2880_ (.A1(\mem[1][13] ),
    .A2(_0761_),
    .ZN(_0900_));
 BUF_X4 _2881_ (.A(_0783_),
    .Z(_0901_));
 MUX2_X1 _2882_ (.A(_0899_),
    .B(_0900_),
    .S(_0901_),
    .Z(_0902_));
 OAI22_X1 _2883_ (.A1(_0858_),
    .A2(_0898_),
    .B1(_0902_),
    .B2(_0867_),
    .ZN(_0903_));
 OAI33_X1 _2884_ (.A1(\mem[0][13] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0890_),
    .B2(_0897_),
    .B3(_0903_),
    .ZN(_0904_));
 OAI21_X1 _2885_ (.A(_0887_),
    .B1(_0904_),
    .B2(_0810_),
    .ZN(_0522_));
 NAND2_X1 _2886_ (.A1(net17),
    .A2(_0743_),
    .ZN(_0905_));
 OAI21_X1 _2887_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][14] ),
    .ZN(_0906_));
 BUF_X4 _2888_ (.A(_0867_),
    .Z(_0907_));
 BUF_X4 _2889_ (.A(_0760_),
    .Z(_0908_));
 AOI222_X2 _2890_ (.A1(\mem[6][14] ),
    .A2(_0823_),
    .B1(_0908_),
    .B2(\mem[5][14] ),
    .C1(\mem[4][14] ),
    .C2(_0879_),
    .ZN(_0909_));
 BUF_X4 _2891_ (.A(_0757_),
    .Z(_0910_));
 BUF_X4 _2892_ (.A(_0759_),
    .Z(_0911_));
 AOI222_X2 _2893_ (.A1(_0764_),
    .A2(\mem[3][14] ),
    .B1(\mem[2][14] ),
    .B2(_0910_),
    .C1(_0911_),
    .C2(\mem[1][14] ),
    .ZN(_0912_));
 MUX2_X1 _2894_ (.A(_0909_),
    .B(_0912_),
    .S(_0784_),
    .Z(_0913_));
 NOR2_X1 _2895_ (.A1(_0907_),
    .A2(_0913_),
    .ZN(_0914_));
 BUF_X4 _2896_ (.A(_0753_),
    .Z(_0915_));
 BUF_X4 _2897_ (.A(_0745_),
    .Z(_0916_));
 AOI22_X2 _2898_ (.A1(_0915_),
    .A2(\mem[15][14] ),
    .B1(\mem[12][14] ),
    .B2(_0916_),
    .ZN(_0917_));
 BUF_X4 _2899_ (.A(_0757_),
    .Z(_0918_));
 AOI21_X1 _2900_ (.A(_0774_),
    .B1(\mem[14][14] ),
    .B2(_0918_),
    .ZN(_0919_));
 NAND2_X1 _2901_ (.A1(_0804_),
    .A2(\mem[7][14] ),
    .ZN(_0920_));
 BUF_X4 _2902_ (.A(_0774_),
    .Z(_0921_));
 AOI221_X2 _2903_ (.A(_0795_),
    .B1(_0917_),
    .B2(_0919_),
    .C1(_0920_),
    .C2(_0921_),
    .ZN(_0922_));
 NAND2_X1 _2904_ (.A1(_0786_),
    .A2(_0766_),
    .ZN(_0923_));
 BUF_X4 _2905_ (.A(_0923_),
    .Z(_0924_));
 INV_X1 _2906_ (.A(\mem[13][14] ),
    .ZN(_0925_));
 OAI21_X1 _2907_ (.A(_0816_),
    .B1(_0924_),
    .B2(_0925_),
    .ZN(_0926_));
 AOI22_X1 _2908_ (.A1(\mem[10][14] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][14] ),
    .ZN(_0927_));
 AOI22_X1 _2909_ (.A1(_0765_),
    .A2(\mem[11][14] ),
    .B1(\mem[8][14] ),
    .B2(_0874_),
    .ZN(_0928_));
 AOI21_X1 _2910_ (.A(_0871_),
    .B1(_0927_),
    .B2(_0928_),
    .ZN(_0929_));
 NOR4_X2 _2911_ (.A1(_0914_),
    .A2(_0922_),
    .A3(_0926_),
    .A4(_0929_),
    .ZN(_0930_));
 OAI21_X1 _2912_ (.A(_0905_),
    .B1(_0906_),
    .B2(_0930_),
    .ZN(_0523_));
 NAND2_X1 _2913_ (.A1(net18),
    .A2(_0743_),
    .ZN(_0931_));
 MUX2_X1 _2914_ (.A(\mem[3][15] ),
    .B(\mem[7][15] ),
    .S(_0840_),
    .Z(_0932_));
 AOI22_X1 _2915_ (.A1(\mem[15][15] ),
    .A2(_0768_),
    .B1(_0932_),
    .B2(_0775_),
    .ZN(_0933_));
 NOR2_X1 _2916_ (.A1(_0839_),
    .A2(_0933_),
    .ZN(_0934_));
 AOI22_X1 _2917_ (.A1(\mem[12][15] ),
    .A2(_0846_),
    .B1(_0891_),
    .B2(\mem[14][15] ),
    .ZN(_0935_));
 OR2_X1 _2918_ (.A1(_0845_),
    .A2(_0935_),
    .ZN(_0936_));
 NAND3_X1 _2919_ (.A1(\mem[2][15] ),
    .A2(_0779_),
    .A3(_0849_),
    .ZN(_0937_));
 MUX2_X1 _2920_ (.A(\mem[9][15] ),
    .B(\mem[13][15] ),
    .S(_0776_),
    .Z(_0938_));
 NAND2_X1 _2921_ (.A1(_0853_),
    .A2(_0938_),
    .ZN(_0939_));
 NAND4_X1 _2922_ (.A1(_0772_),
    .A2(_0936_),
    .A3(_0937_),
    .A4(_0939_),
    .ZN(_0940_));
 BUF_X4 _2923_ (.A(_0861_),
    .Z(_0941_));
 AOI222_X2 _2924_ (.A1(_0859_),
    .A2(\mem[11][15] ),
    .B1(\mem[8][15] ),
    .B2(_0801_),
    .C1(_0941_),
    .C2(\mem[10][15] ),
    .ZN(_0942_));
 AOI222_X2 _2925_ (.A1(\mem[6][15] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][15] ),
    .C1(\mem[4][15] ),
    .C2(_0746_),
    .ZN(_0943_));
 NAND2_X1 _2926_ (.A1(\mem[1][15] ),
    .A2(_0761_),
    .ZN(_0944_));
 MUX2_X1 _2927_ (.A(_0943_),
    .B(_0944_),
    .S(_0901_),
    .Z(_0945_));
 OAI22_X1 _2928_ (.A1(_0858_),
    .A2(_0942_),
    .B1(_0945_),
    .B2(_0867_),
    .ZN(_0946_));
 OAI33_X1 _2929_ (.A1(\mem[0][15] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0934_),
    .B2(_0940_),
    .B3(_0946_),
    .ZN(_0947_));
 OAI21_X1 _2930_ (.A(_0931_),
    .B1(_0947_),
    .B2(_0810_),
    .ZN(_0524_));
 NAND2_X1 _2931_ (.A1(net19),
    .A2(_0743_),
    .ZN(_0948_));
 MUX2_X1 _2932_ (.A(\mem[3][16] ),
    .B(\mem[7][16] ),
    .S(_0840_),
    .Z(_0949_));
 AOI22_X1 _2933_ (.A1(\mem[15][16] ),
    .A2(_0768_),
    .B1(_0949_),
    .B2(_0775_),
    .ZN(_0950_));
 NOR2_X1 _2934_ (.A1(_0839_),
    .A2(_0950_),
    .ZN(_0951_));
 BUF_X4 _2935_ (.A(_0771_),
    .Z(_0952_));
 AOI22_X1 _2936_ (.A1(\mem[12][16] ),
    .A2(_0846_),
    .B1(_0891_),
    .B2(\mem[14][16] ),
    .ZN(_0953_));
 OR2_X1 _2937_ (.A1(_0845_),
    .A2(_0953_),
    .ZN(_0954_));
 NAND3_X1 _2938_ (.A1(\mem[2][16] ),
    .A2(_0779_),
    .A3(_0849_),
    .ZN(_0955_));
 MUX2_X1 _2939_ (.A(\mem[9][16] ),
    .B(\mem[13][16] ),
    .S(_0776_),
    .Z(_0956_));
 NAND2_X1 _2940_ (.A1(_0853_),
    .A2(_0956_),
    .ZN(_0957_));
 NAND4_X1 _2941_ (.A1(_0952_),
    .A2(_0954_),
    .A3(_0955_),
    .A4(_0957_),
    .ZN(_0958_));
 BUF_X4 _2942_ (.A(_0800_),
    .Z(_0959_));
 AOI222_X2 _2943_ (.A1(_0859_),
    .A2(\mem[11][16] ),
    .B1(\mem[8][16] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][16] ),
    .ZN(_0960_));
 AOI222_X2 _2944_ (.A1(\mem[6][16] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][16] ),
    .C1(\mem[4][16] ),
    .C2(_0746_),
    .ZN(_0961_));
 NAND2_X1 _2945_ (.A1(\mem[1][16] ),
    .A2(_0761_),
    .ZN(_0962_));
 MUX2_X1 _2946_ (.A(_0961_),
    .B(_0962_),
    .S(_0901_),
    .Z(_0963_));
 OAI22_X1 _2947_ (.A1(_0858_),
    .A2(_0960_),
    .B1(_0963_),
    .B2(_0867_),
    .ZN(_0964_));
 OAI33_X1 _2948_ (.A1(\mem[0][16] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0951_),
    .B2(_0958_),
    .B3(_0964_),
    .ZN(_0965_));
 OAI21_X1 _2949_ (.A(_0948_),
    .B1(_0965_),
    .B2(_0810_),
    .ZN(_0525_));
 NAND2_X1 _2950_ (.A1(net20),
    .A2(_0743_),
    .ZN(_0966_));
 AOI22_X1 _2951_ (.A1(_0755_),
    .A2(\mem[11][17] ),
    .B1(\mem[8][17] ),
    .B2(_0879_),
    .ZN(_0967_));
 AOI22_X1 _2952_ (.A1(\mem[10][17] ),
    .A2(_0758_),
    .B1(_0761_),
    .B2(\mem[9][17] ),
    .ZN(_0968_));
 AND2_X1 _2953_ (.A1(_0967_),
    .A2(_0968_),
    .ZN(_0969_));
 BUF_X4 _2954_ (.A(_0857_),
    .Z(_0970_));
 AOI22_X1 _2955_ (.A1(\mem[12][17] ),
    .A2(_0874_),
    .B1(_0778_),
    .B2(\mem[14][17] ),
    .ZN(_0971_));
 OAI221_X1 _2956_ (.A(_0772_),
    .B1(_0969_),
    .B2(_0970_),
    .C1(_0971_),
    .C2(_0845_),
    .ZN(_0972_));
 NAND4_X1 _2957_ (.A1(_0782_),
    .A2(_0777_),
    .A3(\mem[13][17] ),
    .A4(_0787_),
    .ZN(_0973_));
 NAND3_X1 _2958_ (.A1(_0784_),
    .A2(\mem[2][17] ),
    .A3(_0872_),
    .ZN(_0974_));
 OAI21_X1 _2959_ (.A(_0973_),
    .B1(_0974_),
    .B2(_0867_),
    .ZN(_0975_));
 MUX2_X1 _2960_ (.A(\mem[3][17] ),
    .B(\mem[7][17] ),
    .S(_0792_),
    .Z(_0976_));
 BUF_X4 _2961_ (.A(_0774_),
    .Z(_0977_));
 AOI22_X1 _2962_ (.A1(\mem[15][17] ),
    .A2(_0767_),
    .B1(_0976_),
    .B2(_0977_),
    .ZN(_0978_));
 BUF_X4 _2963_ (.A(_0760_),
    .Z(_0979_));
 NAND2_X1 _2964_ (.A1(\mem[1][17] ),
    .A2(_0979_),
    .ZN(_0980_));
 AOI222_X2 _2965_ (.A1(\mem[6][17] ),
    .A2(_0861_),
    .B1(_0785_),
    .B2(\mem[5][17] ),
    .C1(\mem[4][17] ),
    .C2(_0746_),
    .ZN(_0981_));
 MUX2_X1 _2966_ (.A(_0980_),
    .B(_0981_),
    .S(_0776_),
    .Z(_0982_));
 BUF_X4 _2967_ (.A(_0781_),
    .Z(_0983_));
 OAI22_X1 _2968_ (.A1(_0805_),
    .A2(_0978_),
    .B1(_0982_),
    .B2(_0983_),
    .ZN(_0984_));
 OAI33_X1 _2969_ (.A1(\mem[0][17] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_0972_),
    .B2(_0975_),
    .B3(_0984_),
    .ZN(_0985_));
 OAI21_X1 _2970_ (.A(_0966_),
    .B1(_0985_),
    .B2(_0810_),
    .ZN(_0526_));
 NAND2_X1 _2971_ (.A1(net21),
    .A2(_0743_),
    .ZN(_0986_));
 OAI21_X1 _2972_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][18] ),
    .ZN(_0987_));
 AOI222_X2 _2973_ (.A1(\mem[6][18] ),
    .A2(_0823_),
    .B1(_0908_),
    .B2(\mem[5][18] ),
    .C1(\mem[4][18] ),
    .C2(_0879_),
    .ZN(_0988_));
 AOI222_X2 _2974_ (.A1(_0764_),
    .A2(\mem[3][18] ),
    .B1(\mem[2][18] ),
    .B2(_0910_),
    .C1(_0911_),
    .C2(\mem[1][18] ),
    .ZN(_0989_));
 MUX2_X1 _2975_ (.A(_0988_),
    .B(_0989_),
    .S(_0784_),
    .Z(_0990_));
 NOR2_X1 _2976_ (.A1(_0907_),
    .A2(_0990_),
    .ZN(_0991_));
 AOI22_X2 _2977_ (.A1(_0915_),
    .A2(\mem[15][18] ),
    .B1(\mem[12][18] ),
    .B2(_0916_),
    .ZN(_0992_));
 AOI21_X1 _2978_ (.A(_0774_),
    .B1(\mem[14][18] ),
    .B2(_0918_),
    .ZN(_0993_));
 NAND2_X1 _2979_ (.A1(_0804_),
    .A2(\mem[7][18] ),
    .ZN(_0994_));
 AOI221_X2 _2980_ (.A(_0795_),
    .B1(_0992_),
    .B2(_0993_),
    .C1(_0994_),
    .C2(_0921_),
    .ZN(_0995_));
 INV_X1 _2981_ (.A(\mem[13][18] ),
    .ZN(_0996_));
 OAI21_X1 _2982_ (.A(_0816_),
    .B1(_0924_),
    .B2(_0996_),
    .ZN(_0997_));
 AOI22_X1 _2983_ (.A1(\mem[10][18] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][18] ),
    .ZN(_0998_));
 AOI22_X1 _2984_ (.A1(_0765_),
    .A2(\mem[11][18] ),
    .B1(\mem[8][18] ),
    .B2(_0874_),
    .ZN(_0999_));
 AOI21_X1 _2985_ (.A(_0871_),
    .B1(_0998_),
    .B2(_0999_),
    .ZN(_1000_));
 NOR4_X2 _2986_ (.A1(_0991_),
    .A2(_0995_),
    .A3(_0997_),
    .A4(_1000_),
    .ZN(_1001_));
 OAI21_X1 _2987_ (.A(_0986_),
    .B1(_0987_),
    .B2(_1001_),
    .ZN(_0527_));
 BUF_X4 _2988_ (.A(_0742_),
    .Z(_1002_));
 NAND2_X1 _2989_ (.A1(net22),
    .A2(_1002_),
    .ZN(_1003_));
 MUX2_X1 _2990_ (.A(\mem[3][19] ),
    .B(\mem[7][19] ),
    .S(_0840_),
    .Z(_1004_));
 AOI22_X1 _2991_ (.A1(\mem[15][19] ),
    .A2(_0768_),
    .B1(_1004_),
    .B2(_0775_),
    .ZN(_1005_));
 NOR2_X1 _2992_ (.A1(_0839_),
    .A2(_1005_),
    .ZN(_1006_));
 AOI22_X1 _2993_ (.A1(\mem[12][19] ),
    .A2(_0846_),
    .B1(_0891_),
    .B2(\mem[14][19] ),
    .ZN(_1007_));
 OR2_X1 _2994_ (.A1(_0845_),
    .A2(_1007_),
    .ZN(_1008_));
 NAND3_X1 _2995_ (.A1(\mem[2][19] ),
    .A2(_0779_),
    .A3(_0849_),
    .ZN(_1009_));
 MUX2_X1 _2996_ (.A(\mem[9][19] ),
    .B(\mem[13][19] ),
    .S(_0776_),
    .Z(_1010_));
 NAND2_X1 _2997_ (.A1(_0853_),
    .A2(_1010_),
    .ZN(_1011_));
 NAND4_X1 _2998_ (.A1(_0952_),
    .A2(_1008_),
    .A3(_1009_),
    .A4(_1011_),
    .ZN(_1012_));
 AOI222_X2 _2999_ (.A1(_0859_),
    .A2(\mem[11][19] ),
    .B1(\mem[8][19] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][19] ),
    .ZN(_1013_));
 AOI222_X2 _3000_ (.A1(\mem[6][19] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][19] ),
    .C1(\mem[4][19] ),
    .C2(_0746_),
    .ZN(_1014_));
 NAND2_X1 _3001_ (.A1(\mem[1][19] ),
    .A2(_0761_),
    .ZN(_1015_));
 MUX2_X1 _3002_ (.A(_1014_),
    .B(_1015_),
    .S(_0901_),
    .Z(_1016_));
 OAI22_X1 _3003_ (.A1(_0858_),
    .A2(_1013_),
    .B1(_1016_),
    .B2(_0983_),
    .ZN(_1017_));
 OAI33_X1 _3004_ (.A1(\mem[0][19] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_1006_),
    .B2(_1012_),
    .B3(_1017_),
    .ZN(_1018_));
 OAI21_X1 _3005_ (.A(_1003_),
    .B1(_1018_),
    .B2(_0810_),
    .ZN(_0528_));
 NAND2_X1 _3006_ (.A1(net23),
    .A2(_1002_),
    .ZN(_1019_));
 MUX2_X1 _3007_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(_0840_),
    .Z(_1020_));
 AOI22_X1 _3008_ (.A1(\mem[15][1] ),
    .A2(_0768_),
    .B1(_1020_),
    .B2(_0775_),
    .ZN(_1021_));
 NOR2_X1 _3009_ (.A1(_0839_),
    .A2(_1021_),
    .ZN(_1022_));
 AOI22_X1 _3010_ (.A1(\mem[12][1] ),
    .A2(_0846_),
    .B1(_0891_),
    .B2(\mem[14][1] ),
    .ZN(_1023_));
 OR2_X1 _3011_ (.A1(_0845_),
    .A2(_1023_),
    .ZN(_1024_));
 BUF_X4 _3012_ (.A(_0778_),
    .Z(_1025_));
 NAND3_X1 _3013_ (.A1(\mem[2][1] ),
    .A2(_1025_),
    .A3(_0849_),
    .ZN(_1026_));
 MUX2_X1 _3014_ (.A(\mem[9][1] ),
    .B(\mem[13][1] ),
    .S(_0776_),
    .Z(_1027_));
 NAND2_X1 _3015_ (.A1(_0853_),
    .A2(_1027_),
    .ZN(_1028_));
 NAND4_X1 _3016_ (.A1(_0952_),
    .A2(_1024_),
    .A3(_1026_),
    .A4(_1028_),
    .ZN(_1029_));
 AOI222_X2 _3017_ (.A1(_0859_),
    .A2(\mem[11][1] ),
    .B1(\mem[8][1] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][1] ),
    .ZN(_1030_));
 BUF_X4 _3018_ (.A(_0745_),
    .Z(_1031_));
 AOI222_X2 _3019_ (.A1(\mem[6][1] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][1] ),
    .C1(\mem[4][1] ),
    .C2(_1031_),
    .ZN(_1032_));
 NAND2_X1 _3020_ (.A1(\mem[1][1] ),
    .A2(_0761_),
    .ZN(_1033_));
 MUX2_X1 _3021_ (.A(_1032_),
    .B(_1033_),
    .S(_0901_),
    .Z(_1034_));
 OAI22_X1 _3022_ (.A1(_0858_),
    .A2(_1030_),
    .B1(_1034_),
    .B2(_0983_),
    .ZN(_1035_));
 OAI33_X1 _3023_ (.A1(\mem[0][1] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_1022_),
    .B2(_1029_),
    .B3(_1035_),
    .ZN(_1036_));
 OAI21_X1 _3024_ (.A(_1019_),
    .B1(_1036_),
    .B2(_0810_),
    .ZN(_0529_));
 NAND2_X1 _3025_ (.A1(net24),
    .A2(_1002_),
    .ZN(_1037_));
 OAI21_X1 _3026_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][20] ),
    .ZN(_1038_));
 AOI222_X2 _3027_ (.A1(\mem[6][20] ),
    .A2(_0823_),
    .B1(_0908_),
    .B2(\mem[5][20] ),
    .C1(\mem[4][20] ),
    .C2(_0879_),
    .ZN(_1039_));
 AOI222_X2 _3028_ (.A1(_0764_),
    .A2(\mem[3][20] ),
    .B1(\mem[2][20] ),
    .B2(_0910_),
    .C1(_0911_),
    .C2(\mem[1][20] ),
    .ZN(_1040_));
 MUX2_X1 _3029_ (.A(_1039_),
    .B(_1040_),
    .S(_0784_),
    .Z(_1041_));
 NOR2_X1 _3030_ (.A1(_0907_),
    .A2(_1041_),
    .ZN(_1042_));
 AOI22_X2 _3031_ (.A1(_0915_),
    .A2(\mem[15][20] ),
    .B1(\mem[12][20] ),
    .B2(_0916_),
    .ZN(_1043_));
 AOI21_X1 _3032_ (.A(_0774_),
    .B1(\mem[14][20] ),
    .B2(_0918_),
    .ZN(_1044_));
 NAND2_X1 _3033_ (.A1(_0804_),
    .A2(\mem[7][20] ),
    .ZN(_1045_));
 AOI221_X2 _3034_ (.A(_0795_),
    .B1(_1043_),
    .B2(_1044_),
    .C1(_1045_),
    .C2(_0977_),
    .ZN(_1046_));
 INV_X1 _3035_ (.A(\mem[13][20] ),
    .ZN(_1047_));
 OAI21_X1 _3036_ (.A(_0816_),
    .B1(_0924_),
    .B2(_1047_),
    .ZN(_1048_));
 AOI22_X1 _3037_ (.A1(\mem[10][20] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][20] ),
    .ZN(_1049_));
 AOI22_X1 _3038_ (.A1(_0765_),
    .A2(\mem[11][20] ),
    .B1(\mem[8][20] ),
    .B2(_0874_),
    .ZN(_1050_));
 AOI21_X1 _3039_ (.A(_0871_),
    .B1(_1049_),
    .B2(_1050_),
    .ZN(_1051_));
 NOR4_X1 _3040_ (.A1(_1042_),
    .A2(_1046_),
    .A3(_1048_),
    .A4(_1051_),
    .ZN(_1052_));
 OAI21_X1 _3041_ (.A(_1037_),
    .B1(_1038_),
    .B2(_1052_),
    .ZN(_0530_));
 NAND2_X1 _3042_ (.A1(net25),
    .A2(_1002_),
    .ZN(_1053_));
 MUX2_X1 _3043_ (.A(\mem[3][21] ),
    .B(\mem[7][21] ),
    .S(_0840_),
    .Z(_1054_));
 AOI22_X1 _3044_ (.A1(\mem[15][21] ),
    .A2(_0768_),
    .B1(_1054_),
    .B2(_0775_),
    .ZN(_1055_));
 NOR2_X1 _3045_ (.A1(_0839_),
    .A2(_1055_),
    .ZN(_1056_));
 BUF_X4 _3046_ (.A(_0800_),
    .Z(_1057_));
 AOI22_X1 _3047_ (.A1(\mem[12][21] ),
    .A2(_1057_),
    .B1(_0891_),
    .B2(\mem[14][21] ),
    .ZN(_1058_));
 OR2_X1 _3048_ (.A1(_0845_),
    .A2(_1058_),
    .ZN(_1059_));
 NAND3_X1 _3049_ (.A1(\mem[2][21] ),
    .A2(_1025_),
    .A3(_0849_),
    .ZN(_1060_));
 BUF_X4 _3050_ (.A(_0749_),
    .Z(_1061_));
 MUX2_X1 _3051_ (.A(\mem[9][21] ),
    .B(\mem[13][21] ),
    .S(_1061_),
    .Z(_1062_));
 NAND2_X1 _3052_ (.A1(_0853_),
    .A2(_1062_),
    .ZN(_1063_));
 NAND4_X1 _3053_ (.A1(_0952_),
    .A2(_1059_),
    .A3(_1060_),
    .A4(_1063_),
    .ZN(_1064_));
 BUF_X4 _3054_ (.A(_0754_),
    .Z(_1065_));
 AOI222_X2 _3055_ (.A1(_1065_),
    .A2(\mem[11][21] ),
    .B1(\mem[8][21] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][21] ),
    .ZN(_1066_));
 AOI222_X2 _3056_ (.A1(\mem[6][21] ),
    .A2(_0861_),
    .B1(_0862_),
    .B2(\mem[5][21] ),
    .C1(\mem[4][21] ),
    .C2(_1031_),
    .ZN(_1067_));
 NAND2_X1 _3057_ (.A1(\mem[1][21] ),
    .A2(_0761_),
    .ZN(_1068_));
 MUX2_X1 _3058_ (.A(_1067_),
    .B(_1068_),
    .S(_0901_),
    .Z(_1069_));
 OAI22_X1 _3059_ (.A1(_0858_),
    .A2(_1066_),
    .B1(_1069_),
    .B2(_0983_),
    .ZN(_1070_));
 OAI33_X1 _3060_ (.A1(\mem[0][21] ),
    .A2(_0752_),
    .A3(_0763_),
    .B1(_1056_),
    .B2(_1064_),
    .B3(_1070_),
    .ZN(_1071_));
 OAI21_X1 _3061_ (.A(_1053_),
    .B1(_1071_),
    .B2(_0810_),
    .ZN(_0531_));
 NAND2_X1 _3062_ (.A1(net26),
    .A2(_1002_),
    .ZN(_1072_));
 OAI21_X1 _3063_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][22] ),
    .ZN(_1073_));
 AOI222_X2 _3064_ (.A1(\mem[6][22] ),
    .A2(_0823_),
    .B1(_0908_),
    .B2(\mem[5][22] ),
    .C1(\mem[4][22] ),
    .C2(_0879_),
    .ZN(_1074_));
 AOI222_X2 _3065_ (.A1(_0764_),
    .A2(\mem[3][22] ),
    .B1(\mem[2][22] ),
    .B2(_0910_),
    .C1(_0911_),
    .C2(\mem[1][22] ),
    .ZN(_1075_));
 MUX2_X1 _3066_ (.A(_1074_),
    .B(_1075_),
    .S(_0784_),
    .Z(_1076_));
 NOR2_X1 _3067_ (.A1(_0907_),
    .A2(_1076_),
    .ZN(_1077_));
 AOI22_X2 _3068_ (.A1(_0915_),
    .A2(\mem[15][22] ),
    .B1(\mem[12][22] ),
    .B2(_0916_),
    .ZN(_1078_));
 AOI21_X1 _3069_ (.A(_0774_),
    .B1(\mem[14][22] ),
    .B2(_0918_),
    .ZN(_1079_));
 NAND2_X1 _3070_ (.A1(_0804_),
    .A2(\mem[7][22] ),
    .ZN(_1080_));
 AOI221_X2 _3071_ (.A(_0865_),
    .B1(_1078_),
    .B2(_1079_),
    .C1(_1080_),
    .C2(_0977_),
    .ZN(_1081_));
 INV_X1 _3072_ (.A(\mem[13][22] ),
    .ZN(_1082_));
 OAI21_X1 _3073_ (.A(_0816_),
    .B1(_0924_),
    .B2(_1082_),
    .ZN(_1083_));
 AOI22_X1 _3074_ (.A1(\mem[10][22] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][22] ),
    .ZN(_1084_));
 AOI22_X1 _3075_ (.A1(_0765_),
    .A2(\mem[11][22] ),
    .B1(\mem[8][22] ),
    .B2(_0874_),
    .ZN(_1085_));
 AOI21_X1 _3076_ (.A(_0871_),
    .B1(_1084_),
    .B2(_1085_),
    .ZN(_1086_));
 NOR4_X1 _3077_ (.A1(_1077_),
    .A2(_1081_),
    .A3(_1083_),
    .A4(_1086_),
    .ZN(_1087_));
 OAI21_X1 _3078_ (.A(_1072_),
    .B1(_1073_),
    .B2(_1087_),
    .ZN(_0532_));
 NAND2_X1 _3079_ (.A1(net27),
    .A2(_1002_),
    .ZN(_1088_));
 BUF_X4 _3080_ (.A(_0751_),
    .Z(_1089_));
 BUF_X4 _3081_ (.A(_0762_),
    .Z(_1090_));
 MUX2_X1 _3082_ (.A(\mem[3][23] ),
    .B(\mem[7][23] ),
    .S(_0840_),
    .Z(_1091_));
 AOI22_X1 _3083_ (.A1(\mem[15][23] ),
    .A2(_0768_),
    .B1(_1091_),
    .B2(_0775_),
    .ZN(_1092_));
 NOR2_X1 _3084_ (.A1(_0839_),
    .A2(_1092_),
    .ZN(_1093_));
 AOI22_X1 _3085_ (.A1(\mem[12][23] ),
    .A2(_1057_),
    .B1(_0891_),
    .B2(\mem[14][23] ),
    .ZN(_1094_));
 OR2_X1 _3086_ (.A1(_0844_),
    .A2(_1094_),
    .ZN(_1095_));
 NAND3_X1 _3087_ (.A1(\mem[2][23] ),
    .A2(_1025_),
    .A3(_0849_),
    .ZN(_1096_));
 MUX2_X1 _3088_ (.A(\mem[9][23] ),
    .B(\mem[13][23] ),
    .S(_1061_),
    .Z(_1097_));
 NAND2_X1 _3089_ (.A1(_0853_),
    .A2(_1097_),
    .ZN(_1098_));
 NAND4_X1 _3090_ (.A1(_0952_),
    .A2(_1095_),
    .A3(_1096_),
    .A4(_1098_),
    .ZN(_1099_));
 AOI222_X2 _3091_ (.A1(_1065_),
    .A2(\mem[11][23] ),
    .B1(\mem[8][23] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][23] ),
    .ZN(_1100_));
 AOI222_X2 _3092_ (.A1(\mem[6][23] ),
    .A2(_0832_),
    .B1(_0862_),
    .B2(\mem[5][23] ),
    .C1(\mem[4][23] ),
    .C2(_1031_),
    .ZN(_1101_));
 NAND2_X1 _3093_ (.A1(\mem[1][23] ),
    .A2(_0979_),
    .ZN(_1102_));
 MUX2_X1 _3094_ (.A(_1101_),
    .B(_1102_),
    .S(_0901_),
    .Z(_1103_));
 OAI22_X1 _3095_ (.A1(_0858_),
    .A2(_1100_),
    .B1(_1103_),
    .B2(_0983_),
    .ZN(_1104_));
 OAI33_X1 _3096_ (.A1(\mem[0][23] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1093_),
    .B2(_1099_),
    .B3(_1104_),
    .ZN(_1105_));
 BUF_X4 _3097_ (.A(_0742_),
    .Z(_1106_));
 OAI21_X1 _3098_ (.A(_1088_),
    .B1(_1105_),
    .B2(_1106_),
    .ZN(_0533_));
 NAND2_X1 _3099_ (.A1(net28),
    .A2(_1002_),
    .ZN(_1107_));
 OAI21_X1 _3100_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][24] ),
    .ZN(_1108_));
 AOI222_X2 _3101_ (.A1(\mem[6][24] ),
    .A2(_0823_),
    .B1(_0908_),
    .B2(\mem[5][24] ),
    .C1(\mem[4][24] ),
    .C2(_0879_),
    .ZN(_1109_));
 AOI222_X2 _3102_ (.A1(_0764_),
    .A2(\mem[3][24] ),
    .B1(\mem[2][24] ),
    .B2(_0910_),
    .C1(_0911_),
    .C2(\mem[1][24] ),
    .ZN(_1110_));
 MUX2_X1 _3103_ (.A(_1109_),
    .B(_1110_),
    .S(_0784_),
    .Z(_1111_));
 NOR2_X1 _3104_ (.A1(_0907_),
    .A2(_1111_),
    .ZN(_1112_));
 AOI22_X2 _3105_ (.A1(_0915_),
    .A2(\mem[15][24] ),
    .B1(\mem[12][24] ),
    .B2(_0916_),
    .ZN(_1113_));
 AOI21_X1 _3106_ (.A(_0774_),
    .B1(\mem[14][24] ),
    .B2(_0793_),
    .ZN(_1114_));
 NAND2_X1 _3107_ (.A1(_0804_),
    .A2(\mem[7][24] ),
    .ZN(_1115_));
 AOI221_X2 _3108_ (.A(_0865_),
    .B1(_1113_),
    .B2(_1114_),
    .C1(_1115_),
    .C2(_0977_),
    .ZN(_1116_));
 INV_X1 _3109_ (.A(\mem[13][24] ),
    .ZN(_1117_));
 OAI21_X1 _3110_ (.A(_0816_),
    .B1(_0924_),
    .B2(_1117_),
    .ZN(_1118_));
 AOI22_X1 _3111_ (.A1(\mem[10][24] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][24] ),
    .ZN(_1119_));
 AOI22_X1 _3112_ (.A1(_0765_),
    .A2(\mem[11][24] ),
    .B1(\mem[8][24] ),
    .B2(_0874_),
    .ZN(_1120_));
 AOI21_X1 _3113_ (.A(_0871_),
    .B1(_1119_),
    .B2(_1120_),
    .ZN(_1121_));
 NOR4_X1 _3114_ (.A1(_1112_),
    .A2(_1116_),
    .A3(_1118_),
    .A4(_1121_),
    .ZN(_1122_));
 OAI21_X1 _3115_ (.A(_1107_),
    .B1(_1108_),
    .B2(_1122_),
    .ZN(_0534_));
 NAND2_X1 _3116_ (.A1(net29),
    .A2(_1002_),
    .ZN(_1123_));
 MUX2_X1 _3117_ (.A(\mem[3][25] ),
    .B(\mem[7][25] ),
    .S(_0840_),
    .Z(_1124_));
 AOI22_X1 _3118_ (.A1(\mem[15][25] ),
    .A2(_0768_),
    .B1(_1124_),
    .B2(_0921_),
    .ZN(_1125_));
 NOR2_X1 _3119_ (.A1(_0839_),
    .A2(_1125_),
    .ZN(_1126_));
 AOI22_X1 _3120_ (.A1(\mem[12][25] ),
    .A2(_1057_),
    .B1(_0891_),
    .B2(\mem[14][25] ),
    .ZN(_1127_));
 OR2_X1 _3121_ (.A1(_0844_),
    .A2(_1127_),
    .ZN(_1128_));
 NAND3_X1 _3122_ (.A1(\mem[2][25] ),
    .A2(_1025_),
    .A3(_0849_),
    .ZN(_1129_));
 MUX2_X1 _3123_ (.A(\mem[9][25] ),
    .B(\mem[13][25] ),
    .S(_1061_),
    .Z(_1130_));
 NAND2_X1 _3124_ (.A1(_0853_),
    .A2(_1130_),
    .ZN(_1131_));
 NAND4_X1 _3125_ (.A1(_0952_),
    .A2(_1128_),
    .A3(_1129_),
    .A4(_1131_),
    .ZN(_1132_));
 AOI222_X2 _3126_ (.A1(_1065_),
    .A2(\mem[11][25] ),
    .B1(\mem[8][25] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][25] ),
    .ZN(_1133_));
 AOI222_X2 _3127_ (.A1(\mem[6][25] ),
    .A2(_0832_),
    .B1(_0862_),
    .B2(\mem[5][25] ),
    .C1(\mem[4][25] ),
    .C2(_1031_),
    .ZN(_1134_));
 NAND2_X1 _3128_ (.A1(\mem[1][25] ),
    .A2(_0979_),
    .ZN(_1135_));
 MUX2_X1 _3129_ (.A(_1134_),
    .B(_1135_),
    .S(_0901_),
    .Z(_1136_));
 OAI22_X1 _3130_ (.A1(_0970_),
    .A2(_1133_),
    .B1(_1136_),
    .B2(_0983_),
    .ZN(_1137_));
 OAI33_X1 _3131_ (.A1(\mem[0][25] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1126_),
    .B2(_1132_),
    .B3(_1137_),
    .ZN(_1138_));
 OAI21_X1 _3132_ (.A(_1123_),
    .B1(_1138_),
    .B2(_1106_),
    .ZN(_0535_));
 NAND2_X1 _3133_ (.A1(net30),
    .A2(_1002_),
    .ZN(_1139_));
 OAI21_X1 _3134_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][26] ),
    .ZN(_1140_));
 AOI222_X2 _3135_ (.A1(\mem[6][26] ),
    .A2(_0758_),
    .B1(_0908_),
    .B2(\mem[5][26] ),
    .C1(\mem[4][26] ),
    .C2(_0879_),
    .ZN(_1141_));
 AOI222_X2 _3136_ (.A1(_0755_),
    .A2(\mem[3][26] ),
    .B1(\mem[2][26] ),
    .B2(_0918_),
    .C1(_0911_),
    .C2(\mem[1][26] ),
    .ZN(_1142_));
 MUX2_X1 _3137_ (.A(_1141_),
    .B(_1142_),
    .S(_0795_),
    .Z(_1143_));
 NOR2_X1 _3138_ (.A1(_0907_),
    .A2(_1143_),
    .ZN(_1144_));
 AOI22_X1 _3139_ (.A1(_0915_),
    .A2(\mem[15][26] ),
    .B1(\mem[12][26] ),
    .B2(_0916_),
    .ZN(_1145_));
 AOI21_X1 _3140_ (.A(_0774_),
    .B1(\mem[14][26] ),
    .B2(_0793_),
    .ZN(_1146_));
 NAND2_X1 _3141_ (.A1(_0804_),
    .A2(\mem[7][26] ),
    .ZN(_1147_));
 AOI221_X1 _3142_ (.A(_0865_),
    .B1(_1145_),
    .B2(_1146_),
    .C1(_1147_),
    .C2(_0977_),
    .ZN(_1148_));
 INV_X1 _3143_ (.A(\mem[13][26] ),
    .ZN(_1149_));
 OAI21_X1 _3144_ (.A(_0816_),
    .B1(_0924_),
    .B2(_1149_),
    .ZN(_1150_));
 AOI22_X1 _3145_ (.A1(\mem[10][26] ),
    .A2(_0872_),
    .B1(_0787_),
    .B2(\mem[9][26] ),
    .ZN(_1151_));
 AOI22_X1 _3146_ (.A1(_0765_),
    .A2(\mem[11][26] ),
    .B1(\mem[8][26] ),
    .B2(_0874_),
    .ZN(_1152_));
 AOI21_X1 _3147_ (.A(_0871_),
    .B1(_1151_),
    .B2(_1152_),
    .ZN(_1153_));
 NOR4_X1 _3148_ (.A1(_1144_),
    .A2(_1148_),
    .A3(_1150_),
    .A4(_1153_),
    .ZN(_1154_));
 OAI21_X1 _3149_ (.A(_1139_),
    .B1(_1140_),
    .B2(_1154_),
    .ZN(_0536_));
 NAND2_X1 _3150_ (.A1(net31),
    .A2(_1002_),
    .ZN(_1155_));
 MUX2_X1 _3151_ (.A(\mem[3][27] ),
    .B(\mem[7][27] ),
    .S(_0840_),
    .Z(_1156_));
 AOI22_X1 _3152_ (.A1(\mem[15][27] ),
    .A2(_0767_),
    .B1(_1156_),
    .B2(_0921_),
    .ZN(_1157_));
 NOR2_X1 _3153_ (.A1(_0839_),
    .A2(_1157_),
    .ZN(_1158_));
 AOI22_X1 _3154_ (.A1(\mem[12][27] ),
    .A2(_1057_),
    .B1(_0891_),
    .B2(\mem[14][27] ),
    .ZN(_1159_));
 OR2_X1 _3155_ (.A1(_0844_),
    .A2(_1159_),
    .ZN(_1160_));
 NAND3_X1 _3156_ (.A1(\mem[2][27] ),
    .A2(_1025_),
    .A3(_0849_),
    .ZN(_1161_));
 MUX2_X1 _3157_ (.A(\mem[9][27] ),
    .B(\mem[13][27] ),
    .S(_1061_),
    .Z(_1162_));
 NAND2_X1 _3158_ (.A1(_0853_),
    .A2(_1162_),
    .ZN(_1163_));
 NAND4_X1 _3159_ (.A1(_0952_),
    .A2(_1160_),
    .A3(_1161_),
    .A4(_1163_),
    .ZN(_1164_));
 AOI222_X2 _3160_ (.A1(_1065_),
    .A2(\mem[11][27] ),
    .B1(\mem[8][27] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][27] ),
    .ZN(_1165_));
 AOI222_X2 _3161_ (.A1(\mem[6][27] ),
    .A2(_0832_),
    .B1(_0862_),
    .B2(\mem[5][27] ),
    .C1(\mem[4][27] ),
    .C2(_1031_),
    .ZN(_1166_));
 NAND2_X1 _3162_ (.A1(\mem[1][27] ),
    .A2(_0979_),
    .ZN(_1167_));
 MUX2_X1 _3163_ (.A(_1166_),
    .B(_1167_),
    .S(_0901_),
    .Z(_1168_));
 OAI22_X1 _3164_ (.A1(_0970_),
    .A2(_1165_),
    .B1(_1168_),
    .B2(_0983_),
    .ZN(_1169_));
 OAI33_X1 _3165_ (.A1(\mem[0][27] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1158_),
    .B2(_1164_),
    .B3(_1169_),
    .ZN(_1170_));
 OAI21_X1 _3166_ (.A(_1155_),
    .B1(_1170_),
    .B2(_1106_),
    .ZN(_0537_));
 CLKBUF_X3 _3167_ (.A(_0742_),
    .Z(_1171_));
 NAND2_X1 _3168_ (.A1(net32),
    .A2(_1171_),
    .ZN(_1172_));
 OAI21_X1 _3169_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][28] ),
    .ZN(_1173_));
 AOI222_X2 _3170_ (.A1(\mem[6][28] ),
    .A2(_0758_),
    .B1(_0908_),
    .B2(\mem[5][28] ),
    .C1(\mem[4][28] ),
    .C2(_0879_),
    .ZN(_1174_));
 AOI222_X2 _3171_ (.A1(_0755_),
    .A2(\mem[3][28] ),
    .B1(\mem[2][28] ),
    .B2(_0918_),
    .C1(_0911_),
    .C2(\mem[1][28] ),
    .ZN(_1175_));
 MUX2_X1 _3172_ (.A(_1174_),
    .B(_1175_),
    .S(_0795_),
    .Z(_1176_));
 NOR2_X1 _3173_ (.A1(_0907_),
    .A2(_1176_),
    .ZN(_1177_));
 AOI22_X1 _3174_ (.A1(_0915_),
    .A2(\mem[15][28] ),
    .B1(\mem[12][28] ),
    .B2(_0800_),
    .ZN(_1178_));
 AOI21_X1 _3175_ (.A(_0773_),
    .B1(\mem[14][28] ),
    .B2(_0793_),
    .ZN(_1179_));
 NAND2_X1 _3176_ (.A1(_0804_),
    .A2(\mem[7][28] ),
    .ZN(_1180_));
 AOI221_X1 _3177_ (.A(_0865_),
    .B1(_1178_),
    .B2(_1179_),
    .C1(_1180_),
    .C2(_0977_),
    .ZN(_1181_));
 INV_X1 _3178_ (.A(\mem[13][28] ),
    .ZN(_1182_));
 OAI21_X1 _3179_ (.A(_0816_),
    .B1(_0924_),
    .B2(_1182_),
    .ZN(_1183_));
 AOI22_X1 _3180_ (.A1(\mem[10][28] ),
    .A2(_0872_),
    .B1(_0786_),
    .B2(\mem[9][28] ),
    .ZN(_1184_));
 AOI22_X1 _3181_ (.A1(_0765_),
    .A2(\mem[11][28] ),
    .B1(\mem[8][28] ),
    .B2(_0874_),
    .ZN(_1185_));
 AOI21_X1 _3182_ (.A(_0871_),
    .B1(_1184_),
    .B2(_1185_),
    .ZN(_1186_));
 NOR4_X1 _3183_ (.A1(_1177_),
    .A2(_1181_),
    .A3(_1183_),
    .A4(_1186_),
    .ZN(_1187_));
 OAI21_X1 _3184_ (.A(_1172_),
    .B1(_1173_),
    .B2(_1187_),
    .ZN(_0538_));
 NAND2_X1 _3185_ (.A1(net33),
    .A2(_1171_),
    .ZN(_1188_));
 MUX2_X1 _3186_ (.A(\mem[3][29] ),
    .B(\mem[7][29] ),
    .S(_0792_),
    .Z(_1189_));
 AOI22_X1 _3187_ (.A1(\mem[15][29] ),
    .A2(_0767_),
    .B1(_1189_),
    .B2(_0921_),
    .ZN(_1190_));
 NOR2_X1 _3188_ (.A1(_0805_),
    .A2(_1190_),
    .ZN(_1191_));
 AOI22_X1 _3189_ (.A1(\mem[12][29] ),
    .A2(_1057_),
    .B1(_0891_),
    .B2(\mem[14][29] ),
    .ZN(_1192_));
 OR2_X1 _3190_ (.A1(_0844_),
    .A2(_1192_),
    .ZN(_1193_));
 NAND3_X1 _3191_ (.A1(\mem[2][29] ),
    .A2(_1025_),
    .A3(_0750_),
    .ZN(_1194_));
 MUX2_X1 _3192_ (.A(\mem[9][29] ),
    .B(\mem[13][29] ),
    .S(_1061_),
    .Z(_1195_));
 NAND2_X1 _3193_ (.A1(_0852_),
    .A2(_1195_),
    .ZN(_1196_));
 NAND4_X1 _3194_ (.A1(_0952_),
    .A2(_1193_),
    .A3(_1194_),
    .A4(_1196_),
    .ZN(_1197_));
 AOI222_X2 _3195_ (.A1(_1065_),
    .A2(\mem[11][29] ),
    .B1(\mem[8][29] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][29] ),
    .ZN(_1198_));
 AOI222_X2 _3196_ (.A1(\mem[6][29] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][29] ),
    .C1(\mem[4][29] ),
    .C2(_1031_),
    .ZN(_1199_));
 NAND2_X1 _3197_ (.A1(\mem[1][29] ),
    .A2(_0979_),
    .ZN(_1200_));
 MUX2_X1 _3198_ (.A(_1199_),
    .B(_1200_),
    .S(_0901_),
    .Z(_1201_));
 OAI22_X1 _3199_ (.A1(_0970_),
    .A2(_1198_),
    .B1(_1201_),
    .B2(_0983_),
    .ZN(_1202_));
 OAI33_X1 _3200_ (.A1(\mem[0][29] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1191_),
    .B2(_1197_),
    .B3(_1202_),
    .ZN(_1203_));
 OAI21_X1 _3201_ (.A(_1188_),
    .B1(_1203_),
    .B2(_1106_),
    .ZN(_0539_));
 NAND2_X1 _3202_ (.A1(net34),
    .A2(_1171_),
    .ZN(_1204_));
 OAI21_X1 _3203_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][2] ),
    .ZN(_1205_));
 AOI222_X2 _3204_ (.A1(\mem[6][2] ),
    .A2(_0758_),
    .B1(_0908_),
    .B2(\mem[5][2] ),
    .C1(\mem[4][2] ),
    .C2(_0916_),
    .ZN(_1206_));
 AOI222_X2 _3205_ (.A1(_0755_),
    .A2(\mem[3][2] ),
    .B1(\mem[2][2] ),
    .B2(_0918_),
    .C1(_0911_),
    .C2(\mem[1][2] ),
    .ZN(_1207_));
 MUX2_X1 _3206_ (.A(_1206_),
    .B(_1207_),
    .S(_0795_),
    .Z(_1208_));
 NOR2_X1 _3207_ (.A1(_0907_),
    .A2(_1208_),
    .ZN(_1209_));
 AOI22_X1 _3208_ (.A1(_0915_),
    .A2(\mem[15][2] ),
    .B1(\mem[12][2] ),
    .B2(_0800_),
    .ZN(_1210_));
 AOI21_X1 _3209_ (.A(_0773_),
    .B1(\mem[14][2] ),
    .B2(_0793_),
    .ZN(_1211_));
 NAND2_X1 _3210_ (.A1(_0764_),
    .A2(\mem[7][2] ),
    .ZN(_1212_));
 AOI221_X1 _3211_ (.A(_0865_),
    .B1(_1210_),
    .B2(_1211_),
    .C1(_1212_),
    .C2(_0977_),
    .ZN(_1213_));
 INV_X1 _3212_ (.A(\mem[13][2] ),
    .ZN(_1214_));
 OAI21_X1 _3213_ (.A(_0772_),
    .B1(_0924_),
    .B2(_1214_),
    .ZN(_1215_));
 AOI22_X1 _3214_ (.A1(\mem[10][2] ),
    .A2(_0779_),
    .B1(_0786_),
    .B2(\mem[9][2] ),
    .ZN(_1216_));
 AOI22_X1 _3215_ (.A1(_0765_),
    .A2(\mem[11][2] ),
    .B1(\mem[8][2] ),
    .B2(_0801_),
    .ZN(_1217_));
 AOI21_X1 _3216_ (.A(_0871_),
    .B1(_1216_),
    .B2(_1217_),
    .ZN(_1218_));
 NOR4_X1 _3217_ (.A1(_1209_),
    .A2(_1213_),
    .A3(_1215_),
    .A4(_1218_),
    .ZN(_1219_));
 OAI21_X1 _3218_ (.A(_1204_),
    .B1(_1205_),
    .B2(_1219_),
    .ZN(_0540_));
 NAND2_X1 _3219_ (.A1(net35),
    .A2(_1171_),
    .ZN(_1220_));
 MUX2_X1 _3220_ (.A(\mem[3][30] ),
    .B(\mem[7][30] ),
    .S(_0792_),
    .Z(_1221_));
 AOI22_X1 _3221_ (.A1(\mem[15][30] ),
    .A2(_0767_),
    .B1(_1221_),
    .B2(_0921_),
    .ZN(_1222_));
 NOR2_X1 _3222_ (.A1(_0805_),
    .A2(_1222_),
    .ZN(_1223_));
 AOI22_X1 _3223_ (.A1(\mem[12][30] ),
    .A2(_1057_),
    .B1(_0910_),
    .B2(\mem[14][30] ),
    .ZN(_1224_));
 OR2_X1 _3224_ (.A1(_0844_),
    .A2(_1224_),
    .ZN(_1225_));
 NAND3_X1 _3225_ (.A1(\mem[2][30] ),
    .A2(_1025_),
    .A3(_0750_),
    .ZN(_1226_));
 MUX2_X1 _3226_ (.A(\mem[9][30] ),
    .B(\mem[13][30] ),
    .S(_1061_),
    .Z(_1227_));
 NAND2_X1 _3227_ (.A1(_0852_),
    .A2(_1227_),
    .ZN(_1228_));
 NAND4_X1 _3228_ (.A1(_0952_),
    .A2(_1225_),
    .A3(_1226_),
    .A4(_1228_),
    .ZN(_1229_));
 AOI222_X2 _3229_ (.A1(_1065_),
    .A2(\mem[11][30] ),
    .B1(\mem[8][30] ),
    .B2(_0959_),
    .C1(_0941_),
    .C2(\mem[10][30] ),
    .ZN(_1230_));
 AOI222_X2 _3230_ (.A1(\mem[6][30] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][30] ),
    .C1(\mem[4][30] ),
    .C2(_1031_),
    .ZN(_1231_));
 NAND2_X1 _3231_ (.A1(\mem[1][30] ),
    .A2(_0979_),
    .ZN(_1232_));
 MUX2_X1 _3232_ (.A(_1231_),
    .B(_1232_),
    .S(_0783_),
    .Z(_1233_));
 OAI22_X1 _3233_ (.A1(_0970_),
    .A2(_1230_),
    .B1(_1233_),
    .B2(_0983_),
    .ZN(_1234_));
 OAI33_X1 _3234_ (.A1(\mem[0][30] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1223_),
    .B2(_1229_),
    .B3(_1234_),
    .ZN(_1235_));
 OAI21_X1 _3235_ (.A(_1220_),
    .B1(_1235_),
    .B2(_1106_),
    .ZN(_0541_));
 NAND2_X1 _3236_ (.A1(net36),
    .A2(_1171_),
    .ZN(_1236_));
 AOI22_X1 _3237_ (.A1(_0755_),
    .A2(\mem[11][31] ),
    .B1(\mem[8][31] ),
    .B2(_0879_),
    .ZN(_1237_));
 AOI22_X1 _3238_ (.A1(\mem[10][31] ),
    .A2(_0758_),
    .B1(_0761_),
    .B2(\mem[9][31] ),
    .ZN(_1238_));
 AND2_X1 _3239_ (.A1(_1237_),
    .A2(_1238_),
    .ZN(_1239_));
 AOI22_X1 _3240_ (.A1(\mem[12][31] ),
    .A2(_0874_),
    .B1(_0778_),
    .B2(\mem[14][31] ),
    .ZN(_1240_));
 OAI221_X1 _3241_ (.A(_0772_),
    .B1(_1239_),
    .B2(_0970_),
    .C1(_1240_),
    .C2(_0845_),
    .ZN(_1241_));
 NAND4_X1 _3242_ (.A1(_0782_),
    .A2(_0777_),
    .A3(\mem[13][31] ),
    .A4(_0787_),
    .ZN(_1242_));
 NAND3_X1 _3243_ (.A1(_0784_),
    .A2(\mem[2][31] ),
    .A3(_0872_),
    .ZN(_1243_));
 OAI21_X1 _3244_ (.A(_1242_),
    .B1(_1243_),
    .B2(_0867_),
    .ZN(_1244_));
 MUX2_X1 _3245_ (.A(\mem[3][31] ),
    .B(\mem[7][31] ),
    .S(_0792_),
    .Z(_1245_));
 AOI22_X1 _3246_ (.A1(\mem[15][31] ),
    .A2(_0767_),
    .B1(_1245_),
    .B2(_0774_),
    .ZN(_1246_));
 NAND2_X1 _3247_ (.A1(\mem[1][31] ),
    .A2(_0908_),
    .ZN(_1247_));
 AOI222_X2 _3248_ (.A1(\mem[6][31] ),
    .A2(_0861_),
    .B1(_0785_),
    .B2(\mem[5][31] ),
    .C1(\mem[4][31] ),
    .C2(_0746_),
    .ZN(_1248_));
 MUX2_X1 _3249_ (.A(_1247_),
    .B(_1248_),
    .S(_0776_),
    .Z(_1249_));
 OAI22_X1 _3250_ (.A1(_0805_),
    .A2(_1246_),
    .B1(_1249_),
    .B2(_0983_),
    .ZN(_1250_));
 OAI33_X1 _3251_ (.A1(\mem[0][31] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1241_),
    .B2(_1244_),
    .B3(_1250_),
    .ZN(_1251_));
 OAI21_X1 _3252_ (.A(_1236_),
    .B1(_1251_),
    .B2(_1106_),
    .ZN(_0542_));
 NAND2_X1 _3253_ (.A1(net37),
    .A2(_1171_),
    .ZN(_1252_));
 MUX2_X1 _3254_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(_0792_),
    .Z(_1253_));
 AOI22_X1 _3255_ (.A1(\mem[15][3] ),
    .A2(_0767_),
    .B1(_1253_),
    .B2(_0921_),
    .ZN(_1254_));
 NOR2_X1 _3256_ (.A1(_0805_),
    .A2(_1254_),
    .ZN(_1255_));
 AOI22_X1 _3257_ (.A1(\mem[12][3] ),
    .A2(_1057_),
    .B1(_0910_),
    .B2(\mem[14][3] ),
    .ZN(_1256_));
 OR2_X1 _3258_ (.A1(_0844_),
    .A2(_1256_),
    .ZN(_1257_));
 NAND3_X1 _3259_ (.A1(\mem[2][3] ),
    .A2(_1025_),
    .A3(_0750_),
    .ZN(_1258_));
 MUX2_X1 _3260_ (.A(\mem[9][3] ),
    .B(\mem[13][3] ),
    .S(_1061_),
    .Z(_1259_));
 NAND2_X1 _3261_ (.A1(_0852_),
    .A2(_1259_),
    .ZN(_1260_));
 NAND4_X1 _3262_ (.A1(_0952_),
    .A2(_1257_),
    .A3(_1258_),
    .A4(_1260_),
    .ZN(_1261_));
 AOI222_X2 _3263_ (.A1(_1065_),
    .A2(\mem[11][3] ),
    .B1(\mem[8][3] ),
    .B2(_0959_),
    .C1(_0823_),
    .C2(\mem[10][3] ),
    .ZN(_1262_));
 AOI222_X2 _3264_ (.A1(\mem[6][3] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][3] ),
    .C1(\mem[4][3] ),
    .C2(_1031_),
    .ZN(_1263_));
 NAND2_X1 _3265_ (.A1(\mem[1][3] ),
    .A2(_0979_),
    .ZN(_1264_));
 MUX2_X1 _3266_ (.A(_1263_),
    .B(_1264_),
    .S(_0783_),
    .Z(_1265_));
 OAI22_X2 _3267_ (.A1(_0970_),
    .A2(_1262_),
    .B1(_1265_),
    .B2(_0782_),
    .ZN(_1266_));
 OAI33_X1 _3268_ (.A1(\mem[0][3] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1255_),
    .B2(_1261_),
    .B3(_1266_),
    .ZN(_1267_));
 OAI21_X1 _3269_ (.A(_1252_),
    .B1(_1267_),
    .B2(_1106_),
    .ZN(_0543_));
 NAND2_X1 _3270_ (.A1(net38),
    .A2(_1171_),
    .ZN(_1268_));
 OAI21_X1 _3271_ (.A(_0815_),
    .B1(_0817_),
    .B2(\mem[0][4] ),
    .ZN(_1269_));
 AOI222_X2 _3272_ (.A1(\mem[6][4] ),
    .A2(_0758_),
    .B1(_0908_),
    .B2(\mem[5][4] ),
    .C1(\mem[4][4] ),
    .C2(_0916_),
    .ZN(_1270_));
 AOI222_X2 _3273_ (.A1(_0755_),
    .A2(\mem[3][4] ),
    .B1(\mem[2][4] ),
    .B2(_0918_),
    .C1(_0785_),
    .C2(\mem[1][4] ),
    .ZN(_1271_));
 MUX2_X1 _3274_ (.A(_1270_),
    .B(_1271_),
    .S(_0795_),
    .Z(_1272_));
 NOR2_X1 _3275_ (.A1(_0907_),
    .A2(_1272_),
    .ZN(_1273_));
 AOI22_X1 _3276_ (.A1(_0915_),
    .A2(\mem[15][4] ),
    .B1(\mem[12][4] ),
    .B2(_0800_),
    .ZN(_1274_));
 AOI21_X1 _3277_ (.A(_0773_),
    .B1(\mem[14][4] ),
    .B2(_0793_),
    .ZN(_1275_));
 NAND2_X1 _3278_ (.A1(_0764_),
    .A2(\mem[7][4] ),
    .ZN(_1276_));
 AOI221_X1 _3279_ (.A(_0865_),
    .B1(_1274_),
    .B2(_1275_),
    .C1(_1276_),
    .C2(_0977_),
    .ZN(_1277_));
 INV_X1 _3280_ (.A(\mem[13][4] ),
    .ZN(_1278_));
 OAI21_X1 _3281_ (.A(_0772_),
    .B1(_0924_),
    .B2(_1278_),
    .ZN(_1279_));
 AOI22_X1 _3282_ (.A1(\mem[10][4] ),
    .A2(_0779_),
    .B1(_0786_),
    .B2(\mem[9][4] ),
    .ZN(_1280_));
 AOI22_X1 _3283_ (.A1(_0859_),
    .A2(\mem[11][4] ),
    .B1(\mem[8][4] ),
    .B2(_0801_),
    .ZN(_1281_));
 AOI21_X1 _3284_ (.A(_0871_),
    .B1(_1280_),
    .B2(_1281_),
    .ZN(_1282_));
 NOR4_X1 _3285_ (.A1(_1273_),
    .A2(_1277_),
    .A3(_1279_),
    .A4(_1282_),
    .ZN(_1283_));
 OAI21_X1 _3286_ (.A(_1268_),
    .B1(_1269_),
    .B2(_1283_),
    .ZN(_0544_));
 NAND2_X1 _3287_ (.A1(net39),
    .A2(_1171_),
    .ZN(_1284_));
 MUX2_X1 _3288_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(_0792_),
    .Z(_1285_));
 AOI22_X1 _3289_ (.A1(\mem[15][5] ),
    .A2(_0767_),
    .B1(_1285_),
    .B2(_0921_),
    .ZN(_1286_));
 NOR2_X1 _3290_ (.A1(_0805_),
    .A2(_1286_),
    .ZN(_1287_));
 AOI22_X1 _3291_ (.A1(\mem[12][5] ),
    .A2(_1057_),
    .B1(_0910_),
    .B2(\mem[14][5] ),
    .ZN(_1288_));
 OR2_X1 _3292_ (.A1(_0844_),
    .A2(_1288_),
    .ZN(_1289_));
 NAND3_X1 _3293_ (.A1(\mem[2][5] ),
    .A2(_1025_),
    .A3(_0750_),
    .ZN(_1290_));
 MUX2_X1 _3294_ (.A(\mem[9][5] ),
    .B(\mem[13][5] ),
    .S(_1061_),
    .Z(_1291_));
 NAND2_X1 _3295_ (.A1(_0852_),
    .A2(_1291_),
    .ZN(_1292_));
 NAND4_X1 _3296_ (.A1(_0771_),
    .A2(_1289_),
    .A3(_1290_),
    .A4(_1292_),
    .ZN(_1293_));
 AOI222_X2 _3297_ (.A1(_1065_),
    .A2(\mem[11][5] ),
    .B1(\mem[8][5] ),
    .B2(_0846_),
    .C1(_0823_),
    .C2(\mem[10][5] ),
    .ZN(_1294_));
 AOI222_X2 _3298_ (.A1(\mem[6][5] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][5] ),
    .C1(\mem[4][5] ),
    .C2(_1031_),
    .ZN(_1295_));
 NAND2_X1 _3299_ (.A1(\mem[1][5] ),
    .A2(_0979_),
    .ZN(_1296_));
 MUX2_X1 _3300_ (.A(_1295_),
    .B(_1296_),
    .S(_0783_),
    .Z(_1297_));
 OAI22_X2 _3301_ (.A1(_0970_),
    .A2(_1294_),
    .B1(_1297_),
    .B2(_0782_),
    .ZN(_1298_));
 OAI33_X1 _3302_ (.A1(\mem[0][5] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1287_),
    .B2(_1293_),
    .B3(_1298_),
    .ZN(_1299_));
 OAI21_X1 _3303_ (.A(_1284_),
    .B1(_1299_),
    .B2(_1106_),
    .ZN(_0545_));
 NAND2_X1 _3304_ (.A1(net40),
    .A2(_1171_),
    .ZN(_1300_));
 CLKBUF_X3 _3305_ (.A(_0814_),
    .Z(_1301_));
 OAI21_X1 _3306_ (.A(_1301_),
    .B1(_0816_),
    .B2(\mem[0][6] ),
    .ZN(_1302_));
 AOI222_X2 _3307_ (.A1(\mem[6][6] ),
    .A2(_0758_),
    .B1(_0911_),
    .B2(\mem[5][6] ),
    .C1(\mem[4][6] ),
    .C2(_0916_),
    .ZN(_1303_));
 AOI222_X2 _3308_ (.A1(_0755_),
    .A2(\mem[3][6] ),
    .B1(\mem[2][6] ),
    .B2(_0918_),
    .C1(_0785_),
    .C2(\mem[1][6] ),
    .ZN(_1304_));
 MUX2_X1 _3309_ (.A(_1303_),
    .B(_1304_),
    .S(_0795_),
    .Z(_1305_));
 NOR2_X1 _3310_ (.A1(_0867_),
    .A2(_1305_),
    .ZN(_1306_));
 AOI22_X2 _3311_ (.A1(_0915_),
    .A2(\mem[15][6] ),
    .B1(\mem[12][6] ),
    .B2(_0800_),
    .ZN(_1307_));
 AOI21_X1 _3312_ (.A(_0773_),
    .B1(\mem[14][6] ),
    .B2(_0793_),
    .ZN(_1308_));
 NAND2_X1 _3313_ (.A1(_0764_),
    .A2(\mem[7][6] ),
    .ZN(_1309_));
 AOI221_X2 _3314_ (.A(_0865_),
    .B1(_1307_),
    .B2(_1308_),
    .C1(_1309_),
    .C2(_0977_),
    .ZN(_1310_));
 INV_X1 _3315_ (.A(\mem[13][6] ),
    .ZN(_1311_));
 OAI21_X1 _3316_ (.A(_0772_),
    .B1(_0924_),
    .B2(_1311_),
    .ZN(_1312_));
 AOI22_X1 _3317_ (.A1(\mem[10][6] ),
    .A2(_0779_),
    .B1(_0786_),
    .B2(\mem[9][6] ),
    .ZN(_1313_));
 AOI22_X1 _3318_ (.A1(_0859_),
    .A2(\mem[11][6] ),
    .B1(\mem[8][6] ),
    .B2(_0801_),
    .ZN(_1314_));
 AOI21_X1 _3319_ (.A(_0858_),
    .B1(_1313_),
    .B2(_1314_),
    .ZN(_1315_));
 NOR4_X1 _3320_ (.A1(_1306_),
    .A2(_1310_),
    .A3(_1312_),
    .A4(_1315_),
    .ZN(_1316_));
 OAI21_X1 _3321_ (.A(_1300_),
    .B1(_1302_),
    .B2(_1316_),
    .ZN(_0546_));
 NAND2_X1 _3322_ (.A1(net41),
    .A2(_1171_),
    .ZN(_1317_));
 MUX2_X1 _3323_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(_0792_),
    .Z(_1318_));
 AOI22_X1 _3324_ (.A1(\mem[15][7] ),
    .A2(_0767_),
    .B1(_1318_),
    .B2(_0921_),
    .ZN(_1319_));
 NOR2_X1 _3325_ (.A1(_0805_),
    .A2(_1319_),
    .ZN(_1320_));
 AOI22_X1 _3326_ (.A1(\mem[12][7] ),
    .A2(_1057_),
    .B1(_0910_),
    .B2(\mem[14][7] ),
    .ZN(_1321_));
 OR2_X1 _3327_ (.A1(_0844_),
    .A2(_1321_),
    .ZN(_1322_));
 NAND3_X1 _3328_ (.A1(\mem[2][7] ),
    .A2(_1025_),
    .A3(_0750_),
    .ZN(_1323_));
 MUX2_X1 _3329_ (.A(\mem[9][7] ),
    .B(\mem[13][7] ),
    .S(_1061_),
    .Z(_1324_));
 NAND2_X1 _3330_ (.A1(_0852_),
    .A2(_1324_),
    .ZN(_1325_));
 NAND4_X1 _3331_ (.A1(_0771_),
    .A2(_1322_),
    .A3(_1323_),
    .A4(_1325_),
    .ZN(_1326_));
 AOI222_X2 _3332_ (.A1(_1065_),
    .A2(\mem[11][7] ),
    .B1(\mem[8][7] ),
    .B2(_0846_),
    .C1(_0823_),
    .C2(\mem[10][7] ),
    .ZN(_1327_));
 AOI222_X2 _3333_ (.A1(\mem[6][7] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][7] ),
    .C1(\mem[4][7] ),
    .C2(_1031_),
    .ZN(_1328_));
 NAND2_X1 _3334_ (.A1(\mem[1][7] ),
    .A2(_0979_),
    .ZN(_1329_));
 MUX2_X1 _3335_ (.A(_1328_),
    .B(_1329_),
    .S(_0783_),
    .Z(_1330_));
 OAI22_X2 _3336_ (.A1(_0970_),
    .A2(_1327_),
    .B1(_1330_),
    .B2(_0782_),
    .ZN(_1331_));
 OAI33_X1 _3337_ (.A1(\mem[0][7] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1320_),
    .B2(_1326_),
    .B3(_1331_),
    .ZN(_1332_));
 OAI21_X1 _3338_ (.A(_1317_),
    .B1(_1332_),
    .B2(_1106_),
    .ZN(_0547_));
 NAND2_X1 _3339_ (.A1(net42),
    .A2(_0742_),
    .ZN(_1333_));
 OAI21_X1 _3340_ (.A(_1301_),
    .B1(_0816_),
    .B2(\mem[0][8] ),
    .ZN(_1334_));
 AOI222_X2 _3341_ (.A1(\mem[6][8] ),
    .A2(_0758_),
    .B1(_0911_),
    .B2(\mem[5][8] ),
    .C1(\mem[4][8] ),
    .C2(_0916_),
    .ZN(_1335_));
 AOI222_X2 _3342_ (.A1(_0755_),
    .A2(\mem[3][8] ),
    .B1(\mem[2][8] ),
    .B2(_0918_),
    .C1(_0785_),
    .C2(\mem[1][8] ),
    .ZN(_1336_));
 MUX2_X1 _3343_ (.A(_1335_),
    .B(_1336_),
    .S(_0795_),
    .Z(_1337_));
 NOR2_X1 _3344_ (.A1(_0867_),
    .A2(_1337_),
    .ZN(_1338_));
 AOI22_X2 _3345_ (.A1(_0754_),
    .A2(\mem[15][8] ),
    .B1(\mem[12][8] ),
    .B2(_0800_),
    .ZN(_1339_));
 AOI21_X1 _3346_ (.A(_0773_),
    .B1(\mem[14][8] ),
    .B2(_0793_),
    .ZN(_1340_));
 NAND2_X1 _3347_ (.A1(_0764_),
    .A2(\mem[7][8] ),
    .ZN(_1341_));
 AOI221_X2 _3348_ (.A(_0865_),
    .B1(_1339_),
    .B2(_1340_),
    .C1(_1341_),
    .C2(_0977_),
    .ZN(_1342_));
 INV_X1 _3349_ (.A(\mem[13][8] ),
    .ZN(_1343_));
 OAI21_X1 _3350_ (.A(_0772_),
    .B1(_0923_),
    .B2(_1343_),
    .ZN(_1344_));
 AOI22_X1 _3351_ (.A1(\mem[10][8] ),
    .A2(_0779_),
    .B1(_0786_),
    .B2(\mem[9][8] ),
    .ZN(_1345_));
 AOI22_X1 _3352_ (.A1(_0859_),
    .A2(\mem[11][8] ),
    .B1(\mem[8][8] ),
    .B2(_0801_),
    .ZN(_1346_));
 AOI21_X1 _3353_ (.A(_0858_),
    .B1(_1345_),
    .B2(_1346_),
    .ZN(_1347_));
 NOR4_X1 _3354_ (.A1(_1338_),
    .A2(_1342_),
    .A3(_1344_),
    .A4(_1347_),
    .ZN(_1348_));
 OAI21_X1 _3355_ (.A(_1333_),
    .B1(_1334_),
    .B2(_1348_),
    .ZN(_0548_));
 NAND2_X1 _3356_ (.A1(net43),
    .A2(_0742_),
    .ZN(_1349_));
 MUX2_X1 _3357_ (.A(\mem[3][9] ),
    .B(\mem[7][9] ),
    .S(_0792_),
    .Z(_1350_));
 AOI22_X1 _3358_ (.A1(\mem[15][9] ),
    .A2(_0767_),
    .B1(_1350_),
    .B2(_0921_),
    .ZN(_1351_));
 NOR2_X1 _3359_ (.A1(_0805_),
    .A2(_1351_),
    .ZN(_1352_));
 AOI22_X1 _3360_ (.A1(\mem[12][9] ),
    .A2(_1057_),
    .B1(_0910_),
    .B2(\mem[14][9] ),
    .ZN(_1353_));
 OR2_X1 _3361_ (.A1(_0844_),
    .A2(_1353_),
    .ZN(_1354_));
 NAND3_X1 _3362_ (.A1(\mem[2][9] ),
    .A2(_0778_),
    .A3(_0750_),
    .ZN(_1355_));
 MUX2_X1 _3363_ (.A(\mem[9][9] ),
    .B(\mem[13][9] ),
    .S(_1061_),
    .Z(_1356_));
 NAND2_X1 _3364_ (.A1(_0852_),
    .A2(_1356_),
    .ZN(_1357_));
 NAND4_X1 _3365_ (.A1(_0771_),
    .A2(_1354_),
    .A3(_1355_),
    .A4(_1357_),
    .ZN(_1358_));
 AOI222_X2 _3366_ (.A1(_1065_),
    .A2(\mem[11][9] ),
    .B1(\mem[8][9] ),
    .B2(_0846_),
    .C1(_0823_),
    .C2(\mem[10][9] ),
    .ZN(_1359_));
 AOI222_X2 _3367_ (.A1(\mem[6][9] ),
    .A2(_0832_),
    .B1(_0760_),
    .B2(\mem[5][9] ),
    .C1(\mem[4][9] ),
    .C2(_0745_),
    .ZN(_1360_));
 NAND2_X1 _3368_ (.A1(\mem[1][9] ),
    .A2(_0979_),
    .ZN(_1361_));
 MUX2_X1 _3369_ (.A(_1360_),
    .B(_1361_),
    .S(_0783_),
    .Z(_1362_));
 OAI22_X1 _3370_ (.A1(_0970_),
    .A2(_1359_),
    .B1(_1362_),
    .B2(_0782_),
    .ZN(_1363_));
 OAI33_X1 _3371_ (.A1(\mem[0][9] ),
    .A2(_1089_),
    .A3(_1090_),
    .B1(_1352_),
    .B2(_1358_),
    .B3(_1363_),
    .ZN(_1364_));
 OAI21_X1 _3372_ (.A(_1349_),
    .B1(_1364_),
    .B2(_1106_),
    .ZN(_0549_));
 MUX2_X1 _3373_ (.A(\rd_ptr_bin[0] ),
    .B(_0004_),
    .S(_1301_),
    .Z(_0550_));
 MUX2_X1 _3374_ (.A(\rd_ptr_bin[1] ),
    .B(_0005_),
    .S(_1301_),
    .Z(_0551_));
 XNOR2_X2 _3375_ (.A(_0804_),
    .B(_1990_),
    .ZN(_1365_));
 MUX2_X1 _3376_ (.A(_0777_),
    .B(_1365_),
    .S(_1301_),
    .Z(_0552_));
 NAND3_X1 _3377_ (.A1(_0792_),
    .A2(\rd_ptr_bin[0] ),
    .A3(\rd_ptr_bin[1] ),
    .ZN(_1366_));
 XOR2_X2 _3378_ (.A(_1986_),
    .B(_1366_),
    .Z(_1367_));
 MUX2_X1 _3379_ (.A(_0907_),
    .B(_1367_),
    .S(_1301_),
    .Z(_0553_));
 XNOR2_X1 _3380_ (.A(\rd_ptr_bin[0] ),
    .B(_0005_),
    .ZN(_1368_));
 MUX2_X1 _3381_ (.A(\rd_ptr_gray[0] ),
    .B(_1368_),
    .S(_1301_),
    .Z(_0554_));
 XOR2_X1 _3382_ (.A(_0005_),
    .B(_1365_),
    .Z(_1369_));
 MUX2_X1 _3383_ (.A(\rd_ptr_gray[1] ),
    .B(_1369_),
    .S(_1301_),
    .Z(_0555_));
 XOR2_X1 _3384_ (.A(_1365_),
    .B(_1367_),
    .Z(_1370_));
 MUX2_X1 _3385_ (.A(\rd_ptr_gray[2] ),
    .B(_1370_),
    .S(_1301_),
    .Z(_0556_));
 NAND2_X1 _3386_ (.A1(_0755_),
    .A2(_0766_),
    .ZN(_1371_));
 XOR2_X1 _3387_ (.A(\rd_ptr_bin[4] ),
    .B(_1371_),
    .Z(_1372_));
 XNOR2_X1 _3388_ (.A(_1367_),
    .B(_1372_),
    .ZN(_1373_));
 MUX2_X1 _3389_ (.A(\rd_ptr_gray[3] ),
    .B(_1373_),
    .S(_1301_),
    .Z(_0557_));
 NOR2_X1 _3390_ (.A1(_1371_),
    .A2(_0742_),
    .ZN(_1374_));
 XOR2_X1 _3391_ (.A(\rd_ptr_bin[4] ),
    .B(_1374_),
    .Z(_0558_));
 NAND2_X4 _3392_ (.A1(net4),
    .A2(_0572_),
    .ZN(_1375_));
 MUX2_X1 _3393_ (.A(_0002_),
    .B(\wr_ptr_bin[0] ),
    .S(_1375_),
    .Z(_0559_));
 MUX2_X1 _3394_ (.A(_0003_),
    .B(\wr_ptr_bin[1] ),
    .S(_1375_),
    .Z(_0560_));
 NAND2_X1 _3395_ (.A1(_0599_),
    .A2(_1375_),
    .ZN(_1376_));
 XOR2_X2 _3396_ (.A(_1999_),
    .B(_0000_),
    .Z(_1377_));
 OAI21_X1 _3397_ (.A(_1376_),
    .B1(_1377_),
    .B2(_1375_),
    .ZN(_0561_));
 NAND3_X1 _3398_ (.A1(_0599_),
    .A2(\wr_ptr_bin[0] ),
    .A3(\wr_ptr_bin[1] ),
    .ZN(_1378_));
 XOR2_X2 _3399_ (.A(_0001_),
    .B(_1378_),
    .Z(_1379_));
 MUX2_X1 _3400_ (.A(_1379_),
    .B(\wr_ptr_bin[3] ),
    .S(_1375_),
    .Z(_0562_));
 XNOR2_X1 _3401_ (.A(\wr_ptr_bin[0] ),
    .B(_0003_),
    .ZN(_1380_));
 MUX2_X1 _3402_ (.A(_1380_),
    .B(\wr_ptr_gray[0] ),
    .S(_1375_),
    .Z(_0563_));
 XNOR2_X1 _3403_ (.A(_0003_),
    .B(_1377_),
    .ZN(_1381_));
 MUX2_X1 _3404_ (.A(_1381_),
    .B(\wr_ptr_gray[1] ),
    .S(_1375_),
    .Z(_0564_));
 XNOR2_X1 _3405_ (.A(_1377_),
    .B(_1379_),
    .ZN(_1382_));
 MUX2_X1 _3406_ (.A(_1382_),
    .B(\wr_ptr_gray[2] ),
    .S(_1375_),
    .Z(_0565_));
 NAND2_X1 _3407_ (.A1(_1999_),
    .A2(_0682_),
    .ZN(_1383_));
 XOR2_X1 _3408_ (.A(\wr_ptr_bin[4] ),
    .B(_1383_),
    .Z(_1384_));
 XNOR2_X1 _3409_ (.A(_1379_),
    .B(_1384_),
    .ZN(_1385_));
 MUX2_X1 _3410_ (.A(_1385_),
    .B(\wr_ptr_gray[3] ),
    .S(_1375_),
    .Z(_0566_));
 NOR2_X1 _3411_ (.A1(_1375_),
    .A2(_1383_),
    .ZN(_1386_));
 XOR2_X1 _3412_ (.A(\wr_ptr_bin[4] ),
    .B(_1386_),
    .Z(_0567_));
 NOR2_X1 _3413_ (.A1(_2009_),
    .A2(_1973_),
    .ZN(_1387_));
 OR2_X1 _3414_ (.A1(net9),
    .A2(_1387_),
    .ZN(_1388_));
 NOR4_X1 _3415_ (.A1(net10),
    .A2(net11),
    .A3(net44),
    .A4(_1388_),
    .ZN(net6));
 INV_X1 _3416_ (.A(_1968_),
    .ZN(net47));
 XNOR2_X1 _3417_ (.A(_1967_),
    .B(_0569_),
    .ZN(net48));
 NAND2_X1 _3418_ (.A1(net47),
    .A2(net48),
    .ZN(_1389_));
 OAI21_X1 _3419_ (.A(_0582_),
    .B1(_1389_),
    .B2(_0577_),
    .ZN(net45));
 FA_X1 _3420_ (.A(_1964_),
    .B(_1965_),
    .CI(_1966_),
    .CO(_1967_),
    .S(_1968_));
 FA_X1 _3421_ (.A(\rd_ptr_bin[1] ),
    .B(_1970_),
    .CI(_1971_),
    .CO(_1972_),
    .S(_1973_));
 HA_X1 _3422_ (.A(\wr_ptr_bin[1] ),
    .B(_1969_),
    .CO(_1974_),
    .S(_1975_));
 HA_X1 _3423_ (.A(\wr_ptr_bin[2] ),
    .B(_1976_),
    .CO(_1977_),
    .S(_1978_));
 HA_X1 _3424_ (.A(\wr_ptr_bin[3] ),
    .B(_1979_),
    .CO(_1980_),
    .S(_1981_));
 HA_X1 _3425_ (.A(_1982_),
    .B(_1983_),
    .CO(_1984_),
    .S(_1985_));
 HA_X1 _3426_ (.A(_1986_),
    .B(_1987_),
    .CO(_1988_),
    .S(_1989_));
 HA_X1 _3427_ (.A(_1990_),
    .B(_1991_),
    .CO(_1992_),
    .S(_1993_));
 HA_X1 _3428_ (.A(_0002_),
    .B(_1964_),
    .CO(_1994_),
    .S(_0003_));
 HA_X1 _3429_ (.A(_0002_),
    .B(\wr_ptr_bin[1] ),
    .CO(_1995_),
    .S(_1996_));
 HA_X1 _3430_ (.A(\wr_ptr_bin[0] ),
    .B(_1964_),
    .CO(_1997_),
    .S(_1998_));
 HA_X1 _3431_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .CO(_1999_),
    .S(_2000_));
 HA_X1 _3432_ (.A(_0004_),
    .B(_1982_),
    .CO(_2001_),
    .S(_0005_));
 HA_X1 _3433_ (.A(_0004_),
    .B(\rd_ptr_bin[1] ),
    .CO(_2002_),
    .S(_2003_));
 HA_X1 _3434_ (.A(\rd_ptr_bin[0] ),
    .B(_1982_),
    .CO(_2004_),
    .S(_2005_));
 HA_X1 _3435_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .CO(_2006_),
    .S(_2007_));
 HA_X1 _3436_ (.A(\rd_ptr_bin[0] ),
    .B(_2008_),
    .CO(_1970_),
    .S(_2009_));
 HA_X1 _3437_ (.A(_0002_),
    .B(_2010_),
    .CO(_1965_),
    .S(_2011_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0006_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[0][0] ),
    .QN(_1943_));
 DFF_X1 \mem[0][10]$_DFFE_PP_  (.D(_0007_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[0][10] ),
    .QN(_1942_));
 DFF_X1 \mem[0][11]$_DFFE_PP_  (.D(_0008_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[0][11] ),
    .QN(_1941_));
 DFF_X1 \mem[0][12]$_DFFE_PP_  (.D(_0009_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[0][12] ),
    .QN(_1940_));
 DFF_X1 \mem[0][13]$_DFFE_PP_  (.D(_0010_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[0][13] ),
    .QN(_1939_));
 DFF_X1 \mem[0][14]$_DFFE_PP_  (.D(_0011_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[0][14] ),
    .QN(_1938_));
 DFF_X1 \mem[0][15]$_DFFE_PP_  (.D(_0012_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[0][15] ),
    .QN(_1937_));
 DFF_X1 \mem[0][16]$_DFFE_PP_  (.D(_0013_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[0][16] ),
    .QN(_1936_));
 DFF_X1 \mem[0][17]$_DFFE_PP_  (.D(_0014_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[0][17] ),
    .QN(_1935_));
 DFF_X1 \mem[0][18]$_DFFE_PP_  (.D(_0015_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[0][18] ),
    .QN(_1934_));
 DFF_X1 \mem[0][19]$_DFFE_PP_  (.D(_0016_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[0][19] ),
    .QN(_1933_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0017_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[0][1] ),
    .QN(_1932_));
 DFF_X1 \mem[0][20]$_DFFE_PP_  (.D(_0018_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[0][20] ),
    .QN(_1931_));
 DFF_X1 \mem[0][21]$_DFFE_PP_  (.D(_0019_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[0][21] ),
    .QN(_1930_));
 DFF_X1 \mem[0][22]$_DFFE_PP_  (.D(_0020_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[0][22] ),
    .QN(_1929_));
 DFF_X1 \mem[0][23]$_DFFE_PP_  (.D(_0021_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[0][23] ),
    .QN(_1928_));
 DFF_X1 \mem[0][24]$_DFFE_PP_  (.D(_0022_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[0][24] ),
    .QN(_1927_));
 DFF_X1 \mem[0][25]$_DFFE_PP_  (.D(_0023_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][25] ),
    .QN(_1926_));
 DFF_X1 \mem[0][26]$_DFFE_PP_  (.D(_0024_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[0][26] ),
    .QN(_1925_));
 DFF_X1 \mem[0][27]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[0][27] ),
    .QN(_1924_));
 DFF_X1 \mem[0][28]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[0][28] ),
    .QN(_1923_));
 DFF_X1 \mem[0][29]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[0][29] ),
    .QN(_1922_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0028_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[0][2] ),
    .QN(_1921_));
 DFF_X1 \mem[0][30]$_DFFE_PP_  (.D(_0029_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[0][30] ),
    .QN(_1920_));
 DFF_X1 \mem[0][31]$_DFFE_PP_  (.D(_0030_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[0][31] ),
    .QN(_1919_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0031_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[0][3] ),
    .QN(_1918_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[0][4] ),
    .QN(_1917_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[0][5] ),
    .QN(_1916_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[0][6] ),
    .QN(_1915_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[0][7] ),
    .QN(_1914_));
 DFF_X1 \mem[0][8]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\mem[0][8] ),
    .QN(_1913_));
 DFF_X1 \mem[0][9]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[0][9] ),
    .QN(_1912_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[10][0] ),
    .QN(_1911_));
 DFF_X1 \mem[10][10]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[10][10] ),
    .QN(_1910_));
 DFF_X1 \mem[10][11]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[10][11] ),
    .QN(_1909_));
 DFF_X1 \mem[10][12]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[10][12] ),
    .QN(_1908_));
 DFF_X1 \mem[10][13]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[10][13] ),
    .QN(_1907_));
 DFF_X1 \mem[10][14]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[10][14] ),
    .QN(_1906_));
 DFF_X1 \mem[10][15]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[10][15] ),
    .QN(_1905_));
 DFF_X1 \mem[10][16]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[10][16] ),
    .QN(_1904_));
 DFF_X1 \mem[10][17]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[10][17] ),
    .QN(_1903_));
 DFF_X1 \mem[10][18]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[10][18] ),
    .QN(_1902_));
 DFF_X1 \mem[10][19]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[10][19] ),
    .QN(_1901_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[10][1] ),
    .QN(_1900_));
 DFF_X1 \mem[10][20]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[10][20] ),
    .QN(_1899_));
 DFF_X1 \mem[10][21]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[10][21] ),
    .QN(_1898_));
 DFF_X1 \mem[10][22]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[10][22] ),
    .QN(_1897_));
 DFF_X1 \mem[10][23]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[10][23] ),
    .QN(_1896_));
 DFF_X1 \mem[10][24]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[10][24] ),
    .QN(_1895_));
 DFF_X1 \mem[10][25]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[10][25] ),
    .QN(_1894_));
 DFF_X1 \mem[10][26]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[10][26] ),
    .QN(_1893_));
 DFF_X1 \mem[10][27]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[10][27] ),
    .QN(_1892_));
 DFF_X1 \mem[10][28]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[10][28] ),
    .QN(_1891_));
 DFF_X1 \mem[10][29]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[10][29] ),
    .QN(_1890_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[10][2] ),
    .QN(_1889_));
 DFF_X1 \mem[10][30]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[10][30] ),
    .QN(_1888_));
 DFF_X1 \mem[10][31]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[10][31] ),
    .QN(_1887_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[10][3] ),
    .QN(_1886_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[10][4] ),
    .QN(_1885_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[10][5] ),
    .QN(_1884_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[10][6] ),
    .QN(_1883_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[10][7] ),
    .QN(_1882_));
 DFF_X1 \mem[10][8]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[10][8] ),
    .QN(_1881_));
 DFF_X1 \mem[10][9]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[10][9] ),
    .QN(_1880_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[11][0] ),
    .QN(_1879_));
 DFF_X1 \mem[11][10]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[11][10] ),
    .QN(_1878_));
 DFF_X1 \mem[11][11]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[11][11] ),
    .QN(_1877_));
 DFF_X1 \mem[11][12]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[11][12] ),
    .QN(_1876_));
 DFF_X1 \mem[11][13]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[11][13] ),
    .QN(_1875_));
 DFF_X1 \mem[11][14]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[11][14] ),
    .QN(_1874_));
 DFF_X1 \mem[11][15]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[11][15] ),
    .QN(_1873_));
 DFF_X1 \mem[11][16]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[11][16] ),
    .QN(_1872_));
 DFF_X1 \mem[11][17]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[11][17] ),
    .QN(_1871_));
 DFF_X1 \mem[11][18]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[11][18] ),
    .QN(_1870_));
 DFF_X1 \mem[11][19]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[11][19] ),
    .QN(_1869_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[11][1] ),
    .QN(_1868_));
 DFF_X1 \mem[11][20]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[11][20] ),
    .QN(_1867_));
 DFF_X1 \mem[11][21]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[11][21] ),
    .QN(_1866_));
 DFF_X1 \mem[11][22]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[11][22] ),
    .QN(_1865_));
 DFF_X1 \mem[11][23]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[11][23] ),
    .QN(_1864_));
 DFF_X1 \mem[11][24]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[11][24] ),
    .QN(_1863_));
 DFF_X1 \mem[11][25]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[11][25] ),
    .QN(_1862_));
 DFF_X1 \mem[11][26]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[11][26] ),
    .QN(_1861_));
 DFF_X1 \mem[11][27]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[11][27] ),
    .QN(_1860_));
 DFF_X1 \mem[11][28]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[11][28] ),
    .QN(_1859_));
 DFF_X1 \mem[11][29]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[11][29] ),
    .QN(_1858_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[11][2] ),
    .QN(_1857_));
 DFF_X1 \mem[11][30]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[11][30] ),
    .QN(_1856_));
 DFF_X1 \mem[11][31]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[11][31] ),
    .QN(_1855_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[11][3] ),
    .QN(_1854_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[11][4] ),
    .QN(_1853_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[11][5] ),
    .QN(_1852_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[11][6] ),
    .QN(_1851_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[11][7] ),
    .QN(_1850_));
 DFF_X1 \mem[11][8]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[11][8] ),
    .QN(_1849_));
 DFF_X1 \mem[11][9]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[11][9] ),
    .QN(_1848_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[12][0] ),
    .QN(_1847_));
 DFF_X1 \mem[12][10]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[12][10] ),
    .QN(_1846_));
 DFF_X1 \mem[12][11]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[12][11] ),
    .QN(_1845_));
 DFF_X1 \mem[12][12]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[12][12] ),
    .QN(_1844_));
 DFF_X1 \mem[12][13]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[12][13] ),
    .QN(_1843_));
 DFF_X1 \mem[12][14]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[12][14] ),
    .QN(_1842_));
 DFF_X1 \mem[12][15]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[12][15] ),
    .QN(_1841_));
 DFF_X1 \mem[12][16]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[12][16] ),
    .QN(_1840_));
 DFF_X1 \mem[12][17]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[12][17] ),
    .QN(_1839_));
 DFF_X1 \mem[12][18]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[12][18] ),
    .QN(_1838_));
 DFF_X1 \mem[12][19]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[12][19] ),
    .QN(_1837_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[12][1] ),
    .QN(_1836_));
 DFF_X1 \mem[12][20]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[12][20] ),
    .QN(_1835_));
 DFF_X1 \mem[12][21]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[12][21] ),
    .QN(_1834_));
 DFF_X1 \mem[12][22]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[12][22] ),
    .QN(_1833_));
 DFF_X1 \mem[12][23]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[12][23] ),
    .QN(_1832_));
 DFF_X1 \mem[12][24]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[12][24] ),
    .QN(_1831_));
 DFF_X1 \mem[12][25]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[12][25] ),
    .QN(_1830_));
 DFF_X1 \mem[12][26]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[12][26] ),
    .QN(_1829_));
 DFF_X1 \mem[12][27]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[12][27] ),
    .QN(_1828_));
 DFF_X1 \mem[12][28]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[12][28] ),
    .QN(_1827_));
 DFF_X1 \mem[12][29]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[12][29] ),
    .QN(_1826_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[12][2] ),
    .QN(_1825_));
 DFF_X1 \mem[12][30]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_leaf_73_wr_clk),
    .Q(\mem[12][30] ),
    .QN(_1824_));
 DFF_X1 \mem[12][31]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[12][31] ),
    .QN(_1823_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[12][3] ),
    .QN(_1822_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[12][4] ),
    .QN(_1821_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[12][5] ),
    .QN(_1820_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[12][6] ),
    .QN(_1819_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[12][7] ),
    .QN(_1818_));
 DFF_X1 \mem[12][8]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\mem[12][8] ),
    .QN(_1817_));
 DFF_X1 \mem[12][9]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[12][9] ),
    .QN(_1816_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[13][0] ),
    .QN(_1815_));
 DFF_X1 \mem[13][10]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[13][10] ),
    .QN(_1814_));
 DFF_X1 \mem[13][11]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[13][11] ),
    .QN(_1813_));
 DFF_X1 \mem[13][12]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[13][12] ),
    .QN(_1812_));
 DFF_X1 \mem[13][13]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[13][13] ),
    .QN(_1811_));
 DFF_X1 \mem[13][14]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[13][14] ),
    .QN(_1810_));
 DFF_X1 \mem[13][15]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[13][15] ),
    .QN(_1809_));
 DFF_X1 \mem[13][16]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[13][16] ),
    .QN(_1808_));
 DFF_X1 \mem[13][17]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[13][17] ),
    .QN(_1807_));
 DFF_X1 \mem[13][18]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[13][18] ),
    .QN(_1806_));
 DFF_X1 \mem[13][19]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[13][19] ),
    .QN(_1805_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[13][1] ),
    .QN(_1804_));
 DFF_X1 \mem[13][20]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[13][20] ),
    .QN(_1803_));
 DFF_X1 \mem[13][21]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[13][21] ),
    .QN(_1802_));
 DFF_X1 \mem[13][22]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[13][22] ),
    .QN(_1801_));
 DFF_X1 \mem[13][23]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[13][23] ),
    .QN(_1800_));
 DFF_X1 \mem[13][24]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[13][24] ),
    .QN(_1799_));
 DFF_X1 \mem[13][25]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[13][25] ),
    .QN(_1798_));
 DFF_X1 \mem[13][26]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[13][26] ),
    .QN(_1797_));
 DFF_X1 \mem[13][27]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[13][27] ),
    .QN(_1796_));
 DFF_X1 \mem[13][28]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[13][28] ),
    .QN(_1795_));
 DFF_X1 \mem[13][29]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[13][29] ),
    .QN(_1794_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[13][2] ),
    .QN(_1793_));
 DFF_X1 \mem[13][30]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[13][30] ),
    .QN(_1792_));
 DFF_X1 \mem[13][31]$_DFFE_PP_  (.D(_0158_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[13][31] ),
    .QN(_1791_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0159_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[13][3] ),
    .QN(_1790_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0160_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[13][4] ),
    .QN(_1789_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0161_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[13][5] ),
    .QN(_1788_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0162_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[13][6] ),
    .QN(_1787_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0163_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[13][7] ),
    .QN(_1786_));
 DFF_X1 \mem[13][8]$_DFFE_PP_  (.D(_0164_),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\mem[13][8] ),
    .QN(_1785_));
 DFF_X1 \mem[13][9]$_DFFE_PP_  (.D(_0165_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[13][9] ),
    .QN(_1784_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[14][0] ),
    .QN(_1783_));
 DFF_X1 \mem[14][10]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[14][10] ),
    .QN(_1782_));
 DFF_X1 \mem[14][11]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[14][11] ),
    .QN(_1781_));
 DFF_X1 \mem[14][12]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[14][12] ),
    .QN(_1780_));
 DFF_X1 \mem[14][13]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[14][13] ),
    .QN(_1779_));
 DFF_X1 \mem[14][14]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[14][14] ),
    .QN(_1778_));
 DFF_X1 \mem[14][15]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[14][15] ),
    .QN(_1777_));
 DFF_X1 \mem[14][16]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[14][16] ),
    .QN(_1776_));
 DFF_X1 \mem[14][17]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[14][17] ),
    .QN(_1775_));
 DFF_X1 \mem[14][18]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[14][18] ),
    .QN(_1774_));
 DFF_X1 \mem[14][19]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[14][19] ),
    .QN(_1773_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[14][1] ),
    .QN(_1772_));
 DFF_X1 \mem[14][20]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[14][20] ),
    .QN(_1771_));
 DFF_X1 \mem[14][21]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[14][21] ),
    .QN(_1770_));
 DFF_X1 \mem[14][22]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[14][22] ),
    .QN(_1769_));
 DFF_X1 \mem[14][23]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[14][23] ),
    .QN(_1768_));
 DFF_X1 \mem[14][24]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[14][24] ),
    .QN(_1767_));
 DFF_X1 \mem[14][25]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[14][25] ),
    .QN(_1766_));
 DFF_X1 \mem[14][26]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[14][26] ),
    .QN(_1765_));
 DFF_X1 \mem[14][27]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[14][27] ),
    .QN(_1764_));
 DFF_X1 \mem[14][28]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[14][28] ),
    .QN(_1763_));
 DFF_X1 \mem[14][29]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[14][29] ),
    .QN(_1762_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[14][2] ),
    .QN(_1761_));
 DFF_X1 \mem[14][30]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_leaf_73_wr_clk),
    .Q(\mem[14][30] ),
    .QN(_1760_));
 DFF_X1 \mem[14][31]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[14][31] ),
    .QN(_1759_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[14][3] ),
    .QN(_1758_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[14][4] ),
    .QN(_1757_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[14][5] ),
    .QN(_1756_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0194_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[14][6] ),
    .QN(_1755_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0195_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[14][7] ),
    .QN(_1754_));
 DFF_X1 \mem[14][8]$_DFFE_PP_  (.D(_0196_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[14][8] ),
    .QN(_1753_));
 DFF_X1 \mem[14][9]$_DFFE_PP_  (.D(_0197_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[14][9] ),
    .QN(_1752_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0198_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[15][0] ),
    .QN(_1751_));
 DFF_X1 \mem[15][10]$_DFFE_PP_  (.D(_0199_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[15][10] ),
    .QN(_1750_));
 DFF_X1 \mem[15][11]$_DFFE_PP_  (.D(_0200_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[15][11] ),
    .QN(_1749_));
 DFF_X1 \mem[15][12]$_DFFE_PP_  (.D(_0201_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[15][12] ),
    .QN(_1748_));
 DFF_X1 \mem[15][13]$_DFFE_PP_  (.D(_0202_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[15][13] ),
    .QN(_1747_));
 DFF_X1 \mem[15][14]$_DFFE_PP_  (.D(_0203_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[15][14] ),
    .QN(_1746_));
 DFF_X1 \mem[15][15]$_DFFE_PP_  (.D(_0204_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[15][15] ),
    .QN(_1745_));
 DFF_X1 \mem[15][16]$_DFFE_PP_  (.D(_0205_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[15][16] ),
    .QN(_1744_));
 DFF_X1 \mem[15][17]$_DFFE_PP_  (.D(_0206_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[15][17] ),
    .QN(_1743_));
 DFF_X1 \mem[15][18]$_DFFE_PP_  (.D(_0207_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[15][18] ),
    .QN(_1742_));
 DFF_X1 \mem[15][19]$_DFFE_PP_  (.D(_0208_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[15][19] ),
    .QN(_1741_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0209_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[15][1] ),
    .QN(_1740_));
 DFF_X1 \mem[15][20]$_DFFE_PP_  (.D(_0210_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[15][20] ),
    .QN(_1739_));
 DFF_X1 \mem[15][21]$_DFFE_PP_  (.D(_0211_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[15][21] ),
    .QN(_1738_));
 DFF_X1 \mem[15][22]$_DFFE_PP_  (.D(_0212_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[15][22] ),
    .QN(_1737_));
 DFF_X1 \mem[15][23]$_DFFE_PP_  (.D(_0213_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[15][23] ),
    .QN(_1736_));
 DFF_X1 \mem[15][24]$_DFFE_PP_  (.D(_0214_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[15][24] ),
    .QN(_1735_));
 DFF_X1 \mem[15][25]$_DFFE_PP_  (.D(_0215_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[15][25] ),
    .QN(_1734_));
 DFF_X1 \mem[15][26]$_DFFE_PP_  (.D(_0216_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[15][26] ),
    .QN(_1733_));
 DFF_X1 \mem[15][27]$_DFFE_PP_  (.D(_0217_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[15][27] ),
    .QN(_1732_));
 DFF_X1 \mem[15][28]$_DFFE_PP_  (.D(_0218_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[15][28] ),
    .QN(_1731_));
 DFF_X1 \mem[15][29]$_DFFE_PP_  (.D(_0219_),
    .CK(clknet_leaf_73_wr_clk),
    .Q(\mem[15][29] ),
    .QN(_1730_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0220_),
    .CK(clknet_leaf_68_wr_clk),
    .Q(\mem[15][2] ),
    .QN(_1729_));
 DFF_X1 \mem[15][30]$_DFFE_PP_  (.D(_0221_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[15][30] ),
    .QN(_1728_));
 DFF_X1 \mem[15][31]$_DFFE_PP_  (.D(_0222_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[15][31] ),
    .QN(_1727_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0223_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[15][3] ),
    .QN(_1726_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0224_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[15][4] ),
    .QN(_1725_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0225_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[15][5] ),
    .QN(_1724_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0226_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[15][6] ),
    .QN(_1723_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0227_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[15][7] ),
    .QN(_1722_));
 DFF_X1 \mem[15][8]$_DFFE_PP_  (.D(_0228_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[15][8] ),
    .QN(_1721_));
 DFF_X1 \mem[15][9]$_DFFE_PP_  (.D(_0229_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[15][9] ),
    .QN(_1720_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0230_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[1][0] ),
    .QN(_1719_));
 DFF_X1 \mem[1][10]$_DFFE_PP_  (.D(_0231_),
    .CK(clknet_leaf_52_wr_clk),
    .Q(\mem[1][10] ),
    .QN(_1718_));
 DFF_X1 \mem[1][11]$_DFFE_PP_  (.D(_0232_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[1][11] ),
    .QN(_1717_));
 DFF_X1 \mem[1][12]$_DFFE_PP_  (.D(_0233_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[1][12] ),
    .QN(_1716_));
 DFF_X1 \mem[1][13]$_DFFE_PP_  (.D(_0234_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[1][13] ),
    .QN(_1715_));
 DFF_X1 \mem[1][14]$_DFFE_PP_  (.D(_0235_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[1][14] ),
    .QN(_1714_));
 DFF_X1 \mem[1][15]$_DFFE_PP_  (.D(_0236_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[1][15] ),
    .QN(_1713_));
 DFF_X1 \mem[1][16]$_DFFE_PP_  (.D(_0237_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[1][16] ),
    .QN(_1712_));
 DFF_X1 \mem[1][17]$_DFFE_PP_  (.D(_0238_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[1][17] ),
    .QN(_1711_));
 DFF_X1 \mem[1][18]$_DFFE_PP_  (.D(_0239_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[1][18] ),
    .QN(_1710_));
 DFF_X1 \mem[1][19]$_DFFE_PP_  (.D(_0240_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[1][19] ),
    .QN(_1709_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0241_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[1][1] ),
    .QN(_1708_));
 DFF_X1 \mem[1][20]$_DFFE_PP_  (.D(_0242_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[1][20] ),
    .QN(_1707_));
 DFF_X1 \mem[1][21]$_DFFE_PP_  (.D(_0243_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[1][21] ),
    .QN(_1706_));
 DFF_X1 \mem[1][22]$_DFFE_PP_  (.D(_0244_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[1][22] ),
    .QN(_1705_));
 DFF_X1 \mem[1][23]$_DFFE_PP_  (.D(_0245_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[1][23] ),
    .QN(_1704_));
 DFF_X1 \mem[1][24]$_DFFE_PP_  (.D(_0246_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[1][24] ),
    .QN(_1703_));
 DFF_X1 \mem[1][25]$_DFFE_PP_  (.D(_0247_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[1][25] ),
    .QN(_1702_));
 DFF_X1 \mem[1][26]$_DFFE_PP_  (.D(_0248_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[1][26] ),
    .QN(_1701_));
 DFF_X1 \mem[1][27]$_DFFE_PP_  (.D(_0249_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[1][27] ),
    .QN(_1700_));
 DFF_X1 \mem[1][28]$_DFFE_PP_  (.D(_0250_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[1][28] ),
    .QN(_1699_));
 DFF_X1 \mem[1][29]$_DFFE_PP_  (.D(_0251_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[1][29] ),
    .QN(_1698_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0252_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[1][2] ),
    .QN(_1697_));
 DFF_X1 \mem[1][30]$_DFFE_PP_  (.D(_0253_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[1][30] ),
    .QN(_1696_));
 DFF_X1 \mem[1][31]$_DFFE_PP_  (.D(_0254_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[1][31] ),
    .QN(_1695_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0255_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[1][3] ),
    .QN(_1694_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0256_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[1][4] ),
    .QN(_1693_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0257_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[1][5] ),
    .QN(_1692_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0258_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[1][6] ),
    .QN(_1691_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0259_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[1][7] ),
    .QN(_1690_));
 DFF_X1 \mem[1][8]$_DFFE_PP_  (.D(_0260_),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\mem[1][8] ),
    .QN(_1689_));
 DFF_X1 \mem[1][9]$_DFFE_PP_  (.D(_0261_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[1][9] ),
    .QN(_1688_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0262_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[2][0] ),
    .QN(_1687_));
 DFF_X1 \mem[2][10]$_DFFE_PP_  (.D(_0263_),
    .CK(clknet_leaf_52_wr_clk),
    .Q(\mem[2][10] ),
    .QN(_1686_));
 DFF_X1 \mem[2][11]$_DFFE_PP_  (.D(_0264_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[2][11] ),
    .QN(_1685_));
 DFF_X1 \mem[2][12]$_DFFE_PP_  (.D(_0265_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[2][12] ),
    .QN(_1684_));
 DFF_X1 \mem[2][13]$_DFFE_PP_  (.D(_0266_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[2][13] ),
    .QN(_1683_));
 DFF_X1 \mem[2][14]$_DFFE_PP_  (.D(_0267_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[2][14] ),
    .QN(_1682_));
 DFF_X1 \mem[2][15]$_DFFE_PP_  (.D(_0268_),
    .CK(clknet_leaf_34_wr_clk),
    .Q(\mem[2][15] ),
    .QN(_1681_));
 DFF_X1 \mem[2][16]$_DFFE_PP_  (.D(_0269_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[2][16] ),
    .QN(_1680_));
 DFF_X1 \mem[2][17]$_DFFE_PP_  (.D(_0270_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[2][17] ),
    .QN(_1679_));
 DFF_X1 \mem[2][18]$_DFFE_PP_  (.D(_0271_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[2][18] ),
    .QN(_1678_));
 DFF_X1 \mem[2][19]$_DFFE_PP_  (.D(_0272_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[2][19] ),
    .QN(_1677_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0273_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[2][1] ),
    .QN(_1676_));
 DFF_X1 \mem[2][20]$_DFFE_PP_  (.D(_0274_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[2][20] ),
    .QN(_1675_));
 DFF_X1 \mem[2][21]$_DFFE_PP_  (.D(_0275_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[2][21] ),
    .QN(_1674_));
 DFF_X1 \mem[2][22]$_DFFE_PP_  (.D(_0276_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[2][22] ),
    .QN(_1673_));
 DFF_X1 \mem[2][23]$_DFFE_PP_  (.D(_0277_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[2][23] ),
    .QN(_1672_));
 DFF_X1 \mem[2][24]$_DFFE_PP_  (.D(_0278_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[2][24] ),
    .QN(_1671_));
 DFF_X1 \mem[2][25]$_DFFE_PP_  (.D(_0279_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[2][25] ),
    .QN(_1670_));
 DFF_X1 \mem[2][26]$_DFFE_PP_  (.D(_0280_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[2][26] ),
    .QN(_1669_));
 DFF_X1 \mem[2][27]$_DFFE_PP_  (.D(_0281_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[2][27] ),
    .QN(_1668_));
 DFF_X1 \mem[2][28]$_DFFE_PP_  (.D(_0282_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[2][28] ),
    .QN(_1667_));
 DFF_X1 \mem[2][29]$_DFFE_PP_  (.D(_0283_),
    .CK(clknet_leaf_73_wr_clk),
    .Q(\mem[2][29] ),
    .QN(_1666_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0284_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[2][2] ),
    .QN(_1665_));
 DFF_X1 \mem[2][30]$_DFFE_PP_  (.D(_0285_),
    .CK(clknet_leaf_73_wr_clk),
    .Q(\mem[2][30] ),
    .QN(_1664_));
 DFF_X1 \mem[2][31]$_DFFE_PP_  (.D(_0286_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[2][31] ),
    .QN(_1663_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0287_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[2][3] ),
    .QN(_1662_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0288_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[2][4] ),
    .QN(_1661_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0289_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[2][5] ),
    .QN(_1660_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0290_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[2][6] ),
    .QN(_1659_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0291_),
    .CK(clknet_leaf_69_wr_clk),
    .Q(\mem[2][7] ),
    .QN(_1658_));
 DFF_X1 \mem[2][8]$_DFFE_PP_  (.D(_0292_),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\mem[2][8] ),
    .QN(_1657_));
 DFF_X1 \mem[2][9]$_DFFE_PP_  (.D(_0293_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[2][9] ),
    .QN(_1656_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0294_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[3][0] ),
    .QN(_1655_));
 DFF_X1 \mem[3][10]$_DFFE_PP_  (.D(_0295_),
    .CK(clknet_leaf_52_wr_clk),
    .Q(\mem[3][10] ),
    .QN(_1654_));
 DFF_X1 \mem[3][11]$_DFFE_PP_  (.D(_0296_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[3][11] ),
    .QN(_1653_));
 DFF_X1 \mem[3][12]$_DFFE_PP_  (.D(_0297_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[3][12] ),
    .QN(_1652_));
 DFF_X1 \mem[3][13]$_DFFE_PP_  (.D(_0298_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[3][13] ),
    .QN(_1651_));
 DFF_X1 \mem[3][14]$_DFFE_PP_  (.D(_0299_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[3][14] ),
    .QN(_1650_));
 DFF_X1 \mem[3][15]$_DFFE_PP_  (.D(_0300_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[3][15] ),
    .QN(_1649_));
 DFF_X1 \mem[3][16]$_DFFE_PP_  (.D(_0301_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[3][16] ),
    .QN(_1648_));
 DFF_X1 \mem[3][17]$_DFFE_PP_  (.D(_0302_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[3][17] ),
    .QN(_1647_));
 DFF_X1 \mem[3][18]$_DFFE_PP_  (.D(_0303_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[3][18] ),
    .QN(_1646_));
 DFF_X1 \mem[3][19]$_DFFE_PP_  (.D(_0304_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[3][19] ),
    .QN(_1645_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0305_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[3][1] ),
    .QN(_1644_));
 DFF_X1 \mem[3][20]$_DFFE_PP_  (.D(_0306_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[3][20] ),
    .QN(_1643_));
 DFF_X1 \mem[3][21]$_DFFE_PP_  (.D(_0307_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[3][21] ),
    .QN(_1642_));
 DFF_X1 \mem[3][22]$_DFFE_PP_  (.D(_0308_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[3][22] ),
    .QN(_1641_));
 DFF_X1 \mem[3][23]$_DFFE_PP_  (.D(_0309_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[3][23] ),
    .QN(_1640_));
 DFF_X1 \mem[3][24]$_DFFE_PP_  (.D(_0310_),
    .CK(clknet_leaf_46_wr_clk),
    .Q(\mem[3][24] ),
    .QN(_1639_));
 DFF_X1 \mem[3][25]$_DFFE_PP_  (.D(_0311_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[3][25] ),
    .QN(_1638_));
 DFF_X1 \mem[3][26]$_DFFE_PP_  (.D(_0312_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[3][26] ),
    .QN(_1637_));
 DFF_X1 \mem[3][27]$_DFFE_PP_  (.D(_0313_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[3][27] ),
    .QN(_1636_));
 DFF_X1 \mem[3][28]$_DFFE_PP_  (.D(_0314_),
    .CK(clknet_leaf_67_wr_clk),
    .Q(\mem[3][28] ),
    .QN(_1635_));
 DFF_X1 \mem[3][29]$_DFFE_PP_  (.D(_0315_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[3][29] ),
    .QN(_1634_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0316_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[3][2] ),
    .QN(_1633_));
 DFF_X1 \mem[3][30]$_DFFE_PP_  (.D(_0317_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[3][30] ),
    .QN(_1632_));
 DFF_X1 \mem[3][31]$_DFFE_PP_  (.D(_0318_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[3][31] ),
    .QN(_1631_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0319_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[3][3] ),
    .QN(_1630_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0320_),
    .CK(clknet_leaf_66_wr_clk),
    .Q(\mem[3][4] ),
    .QN(_1629_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0321_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[3][5] ),
    .QN(_1628_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0322_),
    .CK(clknet_leaf_57_wr_clk),
    .Q(\mem[3][6] ),
    .QN(_1627_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0323_),
    .CK(clknet_leaf_70_wr_clk),
    .Q(\mem[3][7] ),
    .QN(_1626_));
 DFF_X1 \mem[3][8]$_DFFE_PP_  (.D(_0324_),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\mem[3][8] ),
    .QN(_1625_));
 DFF_X1 \mem[3][9]$_DFFE_PP_  (.D(_0325_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[3][9] ),
    .QN(_1624_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0326_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[4][0] ),
    .QN(_1623_));
 DFF_X1 \mem[4][10]$_DFFE_PP_  (.D(_0327_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[4][10] ),
    .QN(_1622_));
 DFF_X1 \mem[4][11]$_DFFE_PP_  (.D(_0328_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[4][11] ),
    .QN(_1621_));
 DFF_X1 \mem[4][12]$_DFFE_PP_  (.D(_0329_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[4][12] ),
    .QN(_1620_));
 DFF_X1 \mem[4][13]$_DFFE_PP_  (.D(_0330_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[4][13] ),
    .QN(_1619_));
 DFF_X1 \mem[4][14]$_DFFE_PP_  (.D(_0331_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[4][14] ),
    .QN(_1618_));
 DFF_X1 \mem[4][15]$_DFFE_PP_  (.D(_0332_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[4][15] ),
    .QN(_1617_));
 DFF_X1 \mem[4][16]$_DFFE_PP_  (.D(_0333_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[4][16] ),
    .QN(_1616_));
 DFF_X1 \mem[4][17]$_DFFE_PP_  (.D(_0334_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[4][17] ),
    .QN(_1615_));
 DFF_X1 \mem[4][18]$_DFFE_PP_  (.D(_0335_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[4][18] ),
    .QN(_1614_));
 DFF_X1 \mem[4][19]$_DFFE_PP_  (.D(_0336_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[4][19] ),
    .QN(_1613_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0337_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[4][1] ),
    .QN(_1612_));
 DFF_X1 \mem[4][20]$_DFFE_PP_  (.D(_0338_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[4][20] ),
    .QN(_1611_));
 DFF_X1 \mem[4][21]$_DFFE_PP_  (.D(_0339_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[4][21] ),
    .QN(_1610_));
 DFF_X1 \mem[4][22]$_DFFE_PP_  (.D(_0340_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[4][22] ),
    .QN(_1609_));
 DFF_X1 \mem[4][23]$_DFFE_PP_  (.D(_0341_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[4][23] ),
    .QN(_1608_));
 DFF_X1 \mem[4][24]$_DFFE_PP_  (.D(_0342_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[4][24] ),
    .QN(_1607_));
 DFF_X1 \mem[4][25]$_DFFE_PP_  (.D(_0343_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[4][25] ),
    .QN(_1606_));
 DFF_X1 \mem[4][26]$_DFFE_PP_  (.D(_0344_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[4][26] ),
    .QN(_1605_));
 DFF_X1 \mem[4][27]$_DFFE_PP_  (.D(_0345_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[4][27] ),
    .QN(_1604_));
 DFF_X1 \mem[4][28]$_DFFE_PP_  (.D(_0346_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[4][28] ),
    .QN(_1603_));
 DFF_X1 \mem[4][29]$_DFFE_PP_  (.D(_0347_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[4][29] ),
    .QN(_1602_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0348_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[4][2] ),
    .QN(_1601_));
 DFF_X1 \mem[4][30]$_DFFE_PP_  (.D(_0349_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[4][30] ),
    .QN(_1600_));
 DFF_X1 \mem[4][31]$_DFFE_PP_  (.D(_0350_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[4][31] ),
    .QN(_1599_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0351_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[4][3] ),
    .QN(_1598_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0352_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[4][4] ),
    .QN(_1597_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0353_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[4][5] ),
    .QN(_1596_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0354_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[4][6] ),
    .QN(_1595_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0355_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[4][7] ),
    .QN(_1594_));
 DFF_X1 \mem[4][8]$_DFFE_PP_  (.D(_0356_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[4][8] ),
    .QN(_1593_));
 DFF_X1 \mem[4][9]$_DFFE_PP_  (.D(_0357_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[4][9] ),
    .QN(_1592_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0358_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[5][0] ),
    .QN(_1591_));
 DFF_X1 \mem[5][10]$_DFFE_PP_  (.D(_0359_),
    .CK(clknet_leaf_52_wr_clk),
    .Q(\mem[5][10] ),
    .QN(_1590_));
 DFF_X1 \mem[5][11]$_DFFE_PP_  (.D(_0360_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[5][11] ),
    .QN(_1589_));
 DFF_X1 \mem[5][12]$_DFFE_PP_  (.D(_0361_),
    .CK(clknet_leaf_40_wr_clk),
    .Q(\mem[5][12] ),
    .QN(_1588_));
 DFF_X1 \mem[5][13]$_DFFE_PP_  (.D(_0362_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[5][13] ),
    .QN(_1587_));
 DFF_X1 \mem[5][14]$_DFFE_PP_  (.D(_0363_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[5][14] ),
    .QN(_1586_));
 DFF_X1 \mem[5][15]$_DFFE_PP_  (.D(_0364_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[5][15] ),
    .QN(_1585_));
 DFF_X1 \mem[5][16]$_DFFE_PP_  (.D(_0365_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[5][16] ),
    .QN(_1584_));
 DFF_X1 \mem[5][17]$_DFFE_PP_  (.D(_0366_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[5][17] ),
    .QN(_1583_));
 DFF_X1 \mem[5][18]$_DFFE_PP_  (.D(_0367_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[5][18] ),
    .QN(_1582_));
 DFF_X1 \mem[5][19]$_DFFE_PP_  (.D(_0368_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[5][19] ),
    .QN(_1581_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0369_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[5][1] ),
    .QN(_1580_));
 DFF_X1 \mem[5][20]$_DFFE_PP_  (.D(_0370_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[5][20] ),
    .QN(_1579_));
 DFF_X1 \mem[5][21]$_DFFE_PP_  (.D(_0371_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[5][21] ),
    .QN(_1578_));
 DFF_X1 \mem[5][22]$_DFFE_PP_  (.D(_0372_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[5][22] ),
    .QN(_1577_));
 DFF_X1 \mem[5][23]$_DFFE_PP_  (.D(_0373_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[5][23] ),
    .QN(_1576_));
 DFF_X1 \mem[5][24]$_DFFE_PP_  (.D(_0374_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[5][24] ),
    .QN(_1575_));
 DFF_X1 \mem[5][25]$_DFFE_PP_  (.D(_0375_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[5][25] ),
    .QN(_1574_));
 DFF_X1 \mem[5][26]$_DFFE_PP_  (.D(_0376_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[5][26] ),
    .QN(_1573_));
 DFF_X1 \mem[5][27]$_DFFE_PP_  (.D(_0377_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[5][27] ),
    .QN(_1572_));
 DFF_X1 \mem[5][28]$_DFFE_PP_  (.D(_0378_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[5][28] ),
    .QN(_1571_));
 DFF_X1 \mem[5][29]$_DFFE_PP_  (.D(_0379_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[5][29] ),
    .QN(_1570_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0380_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[5][2] ),
    .QN(_1569_));
 DFF_X1 \mem[5][30]$_DFFE_PP_  (.D(_0381_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[5][30] ),
    .QN(_1568_));
 DFF_X1 \mem[5][31]$_DFFE_PP_  (.D(_0382_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[5][31] ),
    .QN(_1567_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0383_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[5][3] ),
    .QN(_1566_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0384_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[5][4] ),
    .QN(_1565_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0385_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[5][5] ),
    .QN(_1564_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0386_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[5][6] ),
    .QN(_1563_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0387_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[5][7] ),
    .QN(_1562_));
 DFF_X1 \mem[5][8]$_DFFE_PP_  (.D(_0388_),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\mem[5][8] ),
    .QN(_1561_));
 DFF_X1 \mem[5][9]$_DFFE_PP_  (.D(_0389_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[5][9] ),
    .QN(_1560_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0390_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[6][0] ),
    .QN(_1559_));
 DFF_X1 \mem[6][10]$_DFFE_PP_  (.D(_0391_),
    .CK(clknet_leaf_52_wr_clk),
    .Q(\mem[6][10] ),
    .QN(_1558_));
 DFF_X1 \mem[6][11]$_DFFE_PP_  (.D(_0392_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[6][11] ),
    .QN(_1557_));
 DFF_X1 \mem[6][12]$_DFFE_PP_  (.D(_0393_),
    .CK(clknet_leaf_39_wr_clk),
    .Q(\mem[6][12] ),
    .QN(_1556_));
 DFF_X1 \mem[6][13]$_DFFE_PP_  (.D(_0394_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[6][13] ),
    .QN(_1555_));
 DFF_X1 \mem[6][14]$_DFFE_PP_  (.D(_0395_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[6][14] ),
    .QN(_1554_));
 DFF_X1 \mem[6][15]$_DFFE_PP_  (.D(_0396_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[6][15] ),
    .QN(_1553_));
 DFF_X1 \mem[6][16]$_DFFE_PP_  (.D(_0397_),
    .CK(clknet_leaf_33_wr_clk),
    .Q(\mem[6][16] ),
    .QN(_1552_));
 DFF_X1 \mem[6][17]$_DFFE_PP_  (.D(_0398_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[6][17] ),
    .QN(_1551_));
 DFF_X1 \mem[6][18]$_DFFE_PP_  (.D(_0399_),
    .CK(clknet_leaf_41_wr_clk),
    .Q(\mem[6][18] ),
    .QN(_1550_));
 DFF_X1 \mem[6][19]$_DFFE_PP_  (.D(_0400_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[6][19] ),
    .QN(_1549_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0401_),
    .CK(clknet_leaf_22_wr_clk),
    .Q(\mem[6][1] ),
    .QN(_1548_));
 DFF_X1 \mem[6][20]$_DFFE_PP_  (.D(_0402_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[6][20] ),
    .QN(_1547_));
 DFF_X1 \mem[6][21]$_DFFE_PP_  (.D(_0403_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[6][21] ),
    .QN(_1546_));
 DFF_X1 \mem[6][22]$_DFFE_PP_  (.D(_0404_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[6][22] ),
    .QN(_1545_));
 DFF_X1 \mem[6][23]$_DFFE_PP_  (.D(_0405_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[6][23] ),
    .QN(_1544_));
 DFF_X1 \mem[6][24]$_DFFE_PP_  (.D(_0406_),
    .CK(clknet_leaf_27_wr_clk),
    .Q(\mem[6][24] ),
    .QN(_1543_));
 DFF_X1 \mem[6][25]$_DFFE_PP_  (.D(_0407_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[6][25] ),
    .QN(_1542_));
 DFF_X1 \mem[6][26]$_DFFE_PP_  (.D(_0408_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[6][26] ),
    .QN(_1541_));
 DFF_X1 \mem[6][27]$_DFFE_PP_  (.D(_0409_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[6][27] ),
    .QN(_1540_));
 DFF_X1 \mem[6][28]$_DFFE_PP_  (.D(_0410_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[6][28] ),
    .QN(_1539_));
 DFF_X1 \mem[6][29]$_DFFE_PP_  (.D(_0411_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[6][29] ),
    .QN(_1538_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0412_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[6][2] ),
    .QN(_1537_));
 DFF_X1 \mem[6][30]$_DFFE_PP_  (.D(_0413_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[6][30] ),
    .QN(_1536_));
 DFF_X1 \mem[6][31]$_DFFE_PP_  (.D(_0414_),
    .CK(clknet_leaf_7_wr_clk),
    .Q(\mem[6][31] ),
    .QN(_1535_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0415_),
    .CK(clknet_leaf_12_wr_clk),
    .Q(\mem[6][3] ),
    .QN(_1534_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0416_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[6][4] ),
    .QN(_1533_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0417_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[6][5] ),
    .QN(_1532_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0418_),
    .CK(clknet_leaf_58_wr_clk),
    .Q(\mem[6][6] ),
    .QN(_1531_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0419_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[6][7] ),
    .QN(_1530_));
 DFF_X1 \mem[6][8]$_DFFE_PP_  (.D(_0420_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[6][8] ),
    .QN(_1529_));
 DFF_X1 \mem[6][9]$_DFFE_PP_  (.D(_0421_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[6][9] ),
    .QN(_1528_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0422_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[7][0] ),
    .QN(_1527_));
 DFF_X1 \mem[7][10]$_DFFE_PP_  (.D(_0423_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[7][10] ),
    .QN(_1526_));
 DFF_X1 \mem[7][11]$_DFFE_PP_  (.D(_0424_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[7][11] ),
    .QN(_1525_));
 DFF_X1 \mem[7][12]$_DFFE_PP_  (.D(_0425_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[7][12] ),
    .QN(_1524_));
 DFF_X1 \mem[7][13]$_DFFE_PP_  (.D(_0426_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[7][13] ),
    .QN(_1523_));
 DFF_X1 \mem[7][14]$_DFFE_PP_  (.D(_0427_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[7][14] ),
    .QN(_1522_));
 DFF_X1 \mem[7][15]$_DFFE_PP_  (.D(_0428_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[7][15] ),
    .QN(_1521_));
 DFF_X1 \mem[7][16]$_DFFE_PP_  (.D(_0429_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[7][16] ),
    .QN(_1520_));
 DFF_X1 \mem[7][17]$_DFFE_PP_  (.D(_0430_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[7][17] ),
    .QN(_1519_));
 DFF_X1 \mem[7][18]$_DFFE_PP_  (.D(_0431_),
    .CK(clknet_leaf_45_wr_clk),
    .Q(\mem[7][18] ),
    .QN(_1518_));
 DFF_X1 \mem[7][19]$_DFFE_PP_  (.D(_0432_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[7][19] ),
    .QN(_1517_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0433_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[7][1] ),
    .QN(_1516_));
 DFF_X1 \mem[7][20]$_DFFE_PP_  (.D(_0434_),
    .CK(clknet_leaf_8_wr_clk),
    .Q(\mem[7][20] ),
    .QN(_1515_));
 DFF_X1 \mem[7][21]$_DFFE_PP_  (.D(_0435_),
    .CK(clknet_leaf_19_wr_clk),
    .Q(\mem[7][21] ),
    .QN(_1514_));
 DFF_X1 \mem[7][22]$_DFFE_PP_  (.D(_0436_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[7][22] ),
    .QN(_1513_));
 DFF_X1 \mem[7][23]$_DFFE_PP_  (.D(_0437_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[7][23] ),
    .QN(_1512_));
 DFF_X1 \mem[7][24]$_DFFE_PP_  (.D(_0438_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[7][24] ),
    .QN(_1511_));
 DFF_X1 \mem[7][25]$_DFFE_PP_  (.D(_0439_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[7][25] ),
    .QN(_1510_));
 DFF_X1 \mem[7][26]$_DFFE_PP_  (.D(_0440_),
    .CK(clknet_leaf_26_wr_clk),
    .Q(\mem[7][26] ),
    .QN(_1509_));
 DFF_X1 \mem[7][27]$_DFFE_PP_  (.D(_0441_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[7][27] ),
    .QN(_1508_));
 DFF_X1 \mem[7][28]$_DFFE_PP_  (.D(_0442_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[7][28] ),
    .QN(_1507_));
 DFF_X1 \mem[7][29]$_DFFE_PP_  (.D(_0443_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[7][29] ),
    .QN(_1506_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0444_),
    .CK(clknet_leaf_64_wr_clk),
    .Q(\mem[7][2] ),
    .QN(_1505_));
 DFF_X1 \mem[7][30]$_DFFE_PP_  (.D(_0445_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[7][30] ),
    .QN(_1504_));
 DFF_X1 \mem[7][31]$_DFFE_PP_  (.D(_0446_),
    .CK(clknet_leaf_61_wr_clk),
    .Q(\mem[7][31] ),
    .QN(_1503_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0447_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[7][3] ),
    .QN(_1502_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0448_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[7][4] ),
    .QN(_1501_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0449_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[7][5] ),
    .QN(_1500_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0450_),
    .CK(clknet_leaf_65_wr_clk),
    .Q(\mem[7][6] ),
    .QN(_1499_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0451_),
    .CK(clknet_leaf_72_wr_clk),
    .Q(\mem[7][7] ),
    .QN(_1498_));
 DFF_X1 \mem[7][8]$_DFFE_PP_  (.D(_0452_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[7][8] ),
    .QN(_1497_));
 DFF_X1 \mem[7][9]$_DFFE_PP_  (.D(_0453_),
    .CK(clknet_leaf_59_wr_clk),
    .Q(\mem[7][9] ),
    .QN(_1496_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0454_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[8][0] ),
    .QN(_1495_));
 DFF_X1 \mem[8][10]$_DFFE_PP_  (.D(_0455_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[8][10] ),
    .QN(_1494_));
 DFF_X1 \mem[8][11]$_DFFE_PP_  (.D(_0456_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[8][11] ),
    .QN(_1493_));
 DFF_X1 \mem[8][12]$_DFFE_PP_  (.D(_0457_),
    .CK(clknet_leaf_38_wr_clk),
    .Q(\mem[8][12] ),
    .QN(_1492_));
 DFF_X1 \mem[8][13]$_DFFE_PP_  (.D(_0458_),
    .CK(clknet_leaf_37_wr_clk),
    .Q(\mem[8][13] ),
    .QN(_1491_));
 DFF_X1 \mem[8][14]$_DFFE_PP_  (.D(_0459_),
    .CK(clknet_leaf_50_wr_clk),
    .Q(\mem[8][14] ),
    .QN(_1490_));
 DFF_X1 \mem[8][15]$_DFFE_PP_  (.D(_0460_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[8][15] ),
    .QN(_1489_));
 DFF_X1 \mem[8][16]$_DFFE_PP_  (.D(_0461_),
    .CK(clknet_leaf_29_wr_clk),
    .Q(\mem[8][16] ),
    .QN(_1488_));
 DFF_X1 \mem[8][17]$_DFFE_PP_  (.D(_0462_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[8][17] ),
    .QN(_1487_));
 DFF_X1 \mem[8][18]$_DFFE_PP_  (.D(_0463_),
    .CK(clknet_leaf_42_wr_clk),
    .Q(\mem[8][18] ),
    .QN(_1486_));
 DFF_X1 \mem[8][19]$_DFFE_PP_  (.D(_0464_),
    .CK(clknet_leaf_30_wr_clk),
    .Q(\mem[8][19] ),
    .QN(_1485_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0465_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[8][1] ),
    .QN(_1484_));
 DFF_X1 \mem[8][20]$_DFFE_PP_  (.D(_0466_),
    .CK(clknet_leaf_9_wr_clk),
    .Q(\mem[8][20] ),
    .QN(_1483_));
 DFF_X1 \mem[8][21]$_DFFE_PP_  (.D(_0467_),
    .CK(clknet_leaf_18_wr_clk),
    .Q(\mem[8][21] ),
    .QN(_1482_));
 DFF_X1 \mem[8][22]$_DFFE_PP_  (.D(_0468_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[8][22] ),
    .QN(_1481_));
 DFF_X1 \mem[8][23]$_DFFE_PP_  (.D(_0469_),
    .CK(clknet_leaf_15_wr_clk),
    .Q(\mem[8][23] ),
    .QN(_1480_));
 DFF_X1 \mem[8][24]$_DFFE_PP_  (.D(_0470_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[8][24] ),
    .QN(_1479_));
 DFF_X1 \mem[8][25]$_DFFE_PP_  (.D(_0471_),
    .CK(clknet_leaf_14_wr_clk),
    .Q(\mem[8][25] ),
    .QN(_1478_));
 DFF_X1 \mem[8][26]$_DFFE_PP_  (.D(_0472_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[8][26] ),
    .QN(_1477_));
 DFF_X1 \mem[8][27]$_DFFE_PP_  (.D(_0473_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[8][27] ),
    .QN(_1476_));
 DFF_X1 \mem[8][28]$_DFFE_PP_  (.D(_0474_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[8][28] ),
    .QN(_1475_));
 DFF_X1 \mem[8][29]$_DFFE_PP_  (.D(_0475_),
    .CK(clknet_leaf_11_wr_clk),
    .Q(\mem[8][29] ),
    .QN(_1474_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0476_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[8][2] ),
    .QN(_1473_));
 DFF_X1 \mem[8][30]$_DFFE_PP_  (.D(_0477_),
    .CK(clknet_leaf_2_wr_clk),
    .Q(\mem[8][30] ),
    .QN(_1472_));
 DFF_X1 \mem[8][31]$_DFFE_PP_  (.D(_0478_),
    .CK(clknet_leaf_6_wr_clk),
    .Q(\mem[8][31] ),
    .QN(_1471_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0479_),
    .CK(clknet_leaf_10_wr_clk),
    .Q(\mem[8][3] ),
    .QN(_1470_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0480_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[8][4] ),
    .QN(_1469_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0481_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[8][5] ),
    .QN(_1468_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0482_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[8][6] ),
    .QN(_1467_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0483_),
    .CK(clknet_leaf_3_wr_clk),
    .Q(\mem[8][7] ),
    .QN(_1466_));
 DFF_X1 \mem[8][8]$_DFFE_PP_  (.D(_0484_),
    .CK(clknet_leaf_49_wr_clk),
    .Q(\mem[8][8] ),
    .QN(_1465_));
 DFF_X1 \mem[8][9]$_DFFE_PP_  (.D(_0485_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[8][9] ),
    .QN(_1464_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0486_),
    .CK(clknet_leaf_43_wr_clk),
    .Q(\mem[9][0] ),
    .QN(_1463_));
 DFF_X1 \mem[9][10]$_DFFE_PP_  (.D(_0487_),
    .CK(clknet_leaf_51_wr_clk),
    .Q(\mem[9][10] ),
    .QN(_1462_));
 DFF_X1 \mem[9][11]$_DFFE_PP_  (.D(_0488_),
    .CK(clknet_leaf_35_wr_clk),
    .Q(\mem[9][11] ),
    .QN(_1461_));
 DFF_X1 \mem[9][12]$_DFFE_PP_  (.D(_0489_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[9][12] ),
    .QN(_1460_));
 DFF_X1 \mem[9][13]$_DFFE_PP_  (.D(_0490_),
    .CK(clknet_leaf_36_wr_clk),
    .Q(\mem[9][13] ),
    .QN(_1459_));
 DFF_X1 \mem[9][14]$_DFFE_PP_  (.D(_0491_),
    .CK(clknet_leaf_47_wr_clk),
    .Q(\mem[9][14] ),
    .QN(_1458_));
 DFF_X1 \mem[9][15]$_DFFE_PP_  (.D(_0492_),
    .CK(clknet_leaf_32_wr_clk),
    .Q(\mem[9][15] ),
    .QN(_1457_));
 DFF_X1 \mem[9][16]$_DFFE_PP_  (.D(_0493_),
    .CK(clknet_leaf_31_wr_clk),
    .Q(\mem[9][16] ),
    .QN(_1456_));
 DFF_X1 \mem[9][17]$_DFFE_PP_  (.D(_0494_),
    .CK(clknet_leaf_28_wr_clk),
    .Q(\mem[9][17] ),
    .QN(_1455_));
 DFF_X1 \mem[9][18]$_DFFE_PP_  (.D(_0495_),
    .CK(clknet_leaf_44_wr_clk),
    .Q(\mem[9][18] ),
    .QN(_1454_));
 DFF_X1 \mem[9][19]$_DFFE_PP_  (.D(_0496_),
    .CK(clknet_leaf_21_wr_clk),
    .Q(\mem[9][19] ),
    .QN(_1453_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0497_),
    .CK(clknet_leaf_20_wr_clk),
    .Q(\mem[9][1] ),
    .QN(_1452_));
 DFF_X1 \mem[9][20]$_DFFE_PP_  (.D(_0498_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[9][20] ),
    .QN(_1451_));
 DFF_X1 \mem[9][21]$_DFFE_PP_  (.D(_0499_),
    .CK(clknet_leaf_17_wr_clk),
    .Q(\mem[9][21] ),
    .QN(_1450_));
 DFF_X1 \mem[9][22]$_DFFE_PP_  (.D(_0500_),
    .CK(clknet_leaf_23_wr_clk),
    .Q(\mem[9][22] ),
    .QN(_1449_));
 DFF_X1 \mem[9][23]$_DFFE_PP_  (.D(_0501_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][23] ),
    .QN(_1448_));
 DFF_X1 \mem[9][24]$_DFFE_PP_  (.D(_0502_),
    .CK(clknet_leaf_25_wr_clk),
    .Q(\mem[9][24] ),
    .QN(_1447_));
 DFF_X1 \mem[9][25]$_DFFE_PP_  (.D(_0503_),
    .CK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][25] ),
    .QN(_1446_));
 DFF_X1 \mem[9][26]$_DFFE_PP_  (.D(_0504_),
    .CK(clknet_leaf_24_wr_clk),
    .Q(\mem[9][26] ),
    .QN(_1445_));
 DFF_X1 \mem[9][27]$_DFFE_PP_  (.D(_0505_),
    .CK(clknet_leaf_13_wr_clk),
    .Q(\mem[9][27] ),
    .QN(_1444_));
 DFF_X1 \mem[9][28]$_DFFE_PP_  (.D(_0506_),
    .CK(clknet_leaf_4_wr_clk),
    .Q(\mem[9][28] ),
    .QN(_1443_));
 DFF_X1 \mem[9][29]$_DFFE_PP_  (.D(_0507_),
    .CK(clknet_leaf_1_wr_clk),
    .Q(\mem[9][29] ),
    .QN(_1442_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0508_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[9][2] ),
    .QN(_1441_));
 DFF_X1 \mem[9][30]$_DFFE_PP_  (.D(_0509_),
    .CK(clknet_leaf_0_wr_clk),
    .Q(\mem[9][30] ),
    .QN(_1440_));
 DFF_X1 \mem[9][31]$_DFFE_PP_  (.D(_0510_),
    .CK(clknet_leaf_5_wr_clk),
    .Q(\mem[9][31] ),
    .QN(_1439_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0511_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[9][3] ),
    .QN(_1438_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0512_),
    .CK(clknet_leaf_63_wr_clk),
    .Q(\mem[9][4] ),
    .QN(_1437_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0513_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[9][5] ),
    .QN(_1436_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0514_),
    .CK(clknet_leaf_62_wr_clk),
    .Q(\mem[9][6] ),
    .QN(_1435_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0515_),
    .CK(clknet_leaf_71_wr_clk),
    .Q(\mem[9][7] ),
    .QN(_1434_));
 DFF_X1 \mem[9][8]$_DFFE_PP_  (.D(_0516_),
    .CK(clknet_leaf_48_wr_clk),
    .Q(\mem[9][8] ),
    .QN(_1433_));
 DFF_X1 \mem[9][9]$_DFFE_PP_  (.D(_0517_),
    .CK(clknet_leaf_60_wr_clk),
    .Q(\mem[9][9] ),
    .QN(_1432_));
 DFFR_X1 \rd_data[0]$_DFFE_PN0P_  (.D(_0518_),
    .RN(net3),
    .CK(net1),
    .Q(net12),
    .QN(_1431_));
 DFFR_X1 \rd_data[10]$_DFFE_PN0P_  (.D(_0519_),
    .RN(net3),
    .CK(net1),
    .Q(net13),
    .QN(_1430_));
 DFFR_X1 \rd_data[11]$_DFFE_PN0P_  (.D(_0520_),
    .RN(net3),
    .CK(net1),
    .Q(net14),
    .QN(_1429_));
 DFFR_X1 \rd_data[12]$_DFFE_PN0P_  (.D(_0521_),
    .RN(net3),
    .CK(net1),
    .Q(net15),
    .QN(_1428_));
 DFFR_X1 \rd_data[13]$_DFFE_PN0P_  (.D(_0522_),
    .RN(net3),
    .CK(net1),
    .Q(net16),
    .QN(_1427_));
 DFFR_X1 \rd_data[14]$_DFFE_PN0P_  (.D(_0523_),
    .RN(net3),
    .CK(net1),
    .Q(net17),
    .QN(_1426_));
 DFFR_X1 \rd_data[15]$_DFFE_PN0P_  (.D(_0524_),
    .RN(net3),
    .CK(net1),
    .Q(net18),
    .QN(_1425_));
 DFFR_X1 \rd_data[16]$_DFFE_PN0P_  (.D(_0525_),
    .RN(net3),
    .CK(net1),
    .Q(net19),
    .QN(_1424_));
 DFFR_X1 \rd_data[17]$_DFFE_PN0P_  (.D(_0526_),
    .RN(net3),
    .CK(net1),
    .Q(net20),
    .QN(_1423_));
 DFFR_X1 \rd_data[18]$_DFFE_PN0P_  (.D(_0527_),
    .RN(net3),
    .CK(net1),
    .Q(net21),
    .QN(_1422_));
 DFFR_X1 \rd_data[19]$_DFFE_PN0P_  (.D(_0528_),
    .RN(net3),
    .CK(net1),
    .Q(net22),
    .QN(_1421_));
 DFFR_X1 \rd_data[1]$_DFFE_PN0P_  (.D(_0529_),
    .RN(net3),
    .CK(net1),
    .Q(net23),
    .QN(_1420_));
 DFFR_X1 \rd_data[20]$_DFFE_PN0P_  (.D(_0530_),
    .RN(net3),
    .CK(net1),
    .Q(net24),
    .QN(_1419_));
 DFFR_X1 \rd_data[21]$_DFFE_PN0P_  (.D(_0531_),
    .RN(net3),
    .CK(net1),
    .Q(net25),
    .QN(_1418_));
 DFFR_X1 \rd_data[22]$_DFFE_PN0P_  (.D(_0532_),
    .RN(net3),
    .CK(net1),
    .Q(net26),
    .QN(_1417_));
 DFFR_X1 \rd_data[23]$_DFFE_PN0P_  (.D(_0533_),
    .RN(net3),
    .CK(net1),
    .Q(net27),
    .QN(_1416_));
 DFFR_X1 \rd_data[24]$_DFFE_PN0P_  (.D(_0534_),
    .RN(net3),
    .CK(net1),
    .Q(net28),
    .QN(_1415_));
 DFFR_X1 \rd_data[25]$_DFFE_PN0P_  (.D(_0535_),
    .RN(net3),
    .CK(net1),
    .Q(net29),
    .QN(_1414_));
 DFFR_X1 \rd_data[26]$_DFFE_PN0P_  (.D(_0536_),
    .RN(net3),
    .CK(net1),
    .Q(net30),
    .QN(_1413_));
 DFFR_X1 \rd_data[27]$_DFFE_PN0P_  (.D(_0537_),
    .RN(net3),
    .CK(net1),
    .Q(net31),
    .QN(_1412_));
 DFFR_X1 \rd_data[28]$_DFFE_PN0P_  (.D(_0538_),
    .RN(net3),
    .CK(net1),
    .Q(net32),
    .QN(_1411_));
 DFFR_X1 \rd_data[29]$_DFFE_PN0P_  (.D(_0539_),
    .RN(net3),
    .CK(net1),
    .Q(net33),
    .QN(_1410_));
 DFFR_X1 \rd_data[2]$_DFFE_PN0P_  (.D(_0540_),
    .RN(net3),
    .CK(net1),
    .Q(net34),
    .QN(_1409_));
 DFFR_X1 \rd_data[30]$_DFFE_PN0P_  (.D(_0541_),
    .RN(net3),
    .CK(net1),
    .Q(net35),
    .QN(_1408_));
 DFFR_X1 \rd_data[31]$_DFFE_PN0P_  (.D(_0542_),
    .RN(net3),
    .CK(net1),
    .Q(net36),
    .QN(_1407_));
 DFFR_X1 \rd_data[3]$_DFFE_PN0P_  (.D(_0543_),
    .RN(net3),
    .CK(net1),
    .Q(net37),
    .QN(_1406_));
 DFFR_X1 \rd_data[4]$_DFFE_PN0P_  (.D(_0544_),
    .RN(net3),
    .CK(net1),
    .Q(net38),
    .QN(_1405_));
 DFFR_X1 \rd_data[5]$_DFFE_PN0P_  (.D(_0545_),
    .RN(net3),
    .CK(net1),
    .Q(net39),
    .QN(_1404_));
 DFFR_X1 \rd_data[6]$_DFFE_PN0P_  (.D(_0546_),
    .RN(net3),
    .CK(net1),
    .Q(net40),
    .QN(_1403_));
 DFFR_X1 \rd_data[7]$_DFFE_PN0P_  (.D(_0547_),
    .RN(net3),
    .CK(net1),
    .Q(net41),
    .QN(_1402_));
 DFFR_X1 \rd_data[8]$_DFFE_PN0P_  (.D(_0548_),
    .RN(net3),
    .CK(net1),
    .Q(net42),
    .QN(_1401_));
 DFFR_X1 \rd_data[9]$_DFFE_PN0P_  (.D(_0549_),
    .RN(net3),
    .CK(net1),
    .Q(net43),
    .QN(_1400_));
 DFFR_X2 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_0550_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[0] ),
    .QN(_0004_));
 DFFR_X2 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_0551_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[1] ),
    .QN(_1982_));
 DFFR_X2 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_0552_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[2] ),
    .QN(_1990_));
 DFFR_X1 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_0553_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[3] ),
    .QN(_1986_));
 DFFR_X1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_0554_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[0] ),
    .QN(_1399_));
 DFFR_X1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_0555_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[1] ),
    .QN(_1398_));
 DFFR_X1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_0556_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[2] ),
    .QN(_1397_));
 DFFR_X1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_0557_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_gray[3] ),
    .QN(_1396_));
 DFFR_X2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_0558_),
    .RN(net3),
    .CK(net1),
    .Q(\rd_ptr_bin[4] ),
    .QN(_1944_));
 DFFR_X1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync1[0] ),
    .QN(_1945_));
 DFFR_X1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync1[1] ),
    .QN(_1946_));
 DFFR_X1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync1[2] ),
    .QN(_1947_));
 DFFR_X1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\rd_ptr_gray_sync1[3] ),
    .QN(_1948_));
 DFFR_X1 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\rd_ptr_gray_sync1[4] ),
    .QN(_1949_));
 DFFR_X1 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync2[0] ),
    .QN(_1950_));
 DFFR_X1 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync2[1] ),
    .QN(_1951_));
 DFFR_X1 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .RN(net53),
    .CK(clknet_leaf_53_wr_clk),
    .Q(\rd_ptr_gray_sync2[2] ),
    .QN(_1952_));
 DFFR_X1 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\rd_ptr_gray_sync2[3] ),
    .QN(_1953_));
 DFFR_X2 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\rd_ptr_gray_sync2[4] ),
    .QN(_1395_));
 DFFR_X2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_0559_),
    .RN(net53),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\wr_ptr_bin[0] ),
    .QN(_0002_));
 DFFR_X2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_0560_),
    .RN(net53),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\wr_ptr_bin[1] ),
    .QN(_1964_));
 DFFR_X1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_0561_),
    .RN(net53),
    .CK(clknet_leaf_56_wr_clk),
    .Q(\wr_ptr_bin[2] ),
    .QN(_0000_));
 DFFR_X2 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_0562_),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\wr_ptr_bin[3] ),
    .QN(_0001_));
 DFFR_X1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_0563_),
    .RN(net53),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\wr_ptr_gray[0] ),
    .QN(_1394_));
 DFFR_X1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_0564_),
    .RN(net53),
    .CK(clknet_leaf_55_wr_clk),
    .Q(\wr_ptr_gray[1] ),
    .QN(_1393_));
 DFFR_X1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_0565_),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\wr_ptr_gray[2] ),
    .QN(_1392_));
 DFFR_X1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_0566_),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\wr_ptr_gray[3] ),
    .QN(_1391_));
 DFFR_X2 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_0567_),
    .RN(net53),
    .CK(clknet_leaf_54_wr_clk),
    .Q(\wr_ptr_bin[4] ),
    .QN(_1954_));
 DFFR_X1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[0] ),
    .QN(_1955_));
 DFFR_X1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[1] ),
    .QN(_1956_));
 DFFR_X1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[2] ),
    .QN(_1957_));
 DFFR_X1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[3] ),
    .QN(_1958_));
 DFFR_X1 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync1[4] ),
    .QN(_1959_));
 DFFR_X1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[0] ),
    .QN(_1960_));
 DFFR_X1 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[1] ),
    .QN(_1961_));
 DFFR_X1 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[2] ),
    .QN(_1962_));
 DFFR_X1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[3] ),
    .QN(_1963_));
 DFFR_X1 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .RN(net3),
    .CK(net1),
    .Q(\wr_ptr_gray_sync2[4] ),
    .QN(_1390_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_139 ();
 BUF_X8 input1 (.A(rd_clk),
    .Z(net1));
 BUF_X1 input2 (.A(rd_en),
    .Z(net2));
 BUF_X16 input3 (.A(rd_rst_n),
    .Z(net3));
 BUF_X1 input4 (.A(wr_en),
    .Z(net4));
 BUF_X4 input5 (.A(net55),
    .Z(net5));
 BUF_X1 output6 (.A(net6),
    .Z(rd_almost_empty));
 BUF_X1 output7 (.A(net7),
    .Z(rd_count[0]));
 BUF_X1 output8 (.A(net8),
    .Z(rd_count[1]));
 BUF_X1 output9 (.A(net9),
    .Z(rd_count[2]));
 BUF_X1 output10 (.A(net10),
    .Z(rd_count[3]));
 BUF_X1 output11 (.A(net11),
    .Z(rd_count[4]));
 BUF_X1 output12 (.A(net12),
    .Z(rd_data[0]));
 BUF_X1 output13 (.A(net13),
    .Z(rd_data[10]));
 BUF_X1 output14 (.A(net14),
    .Z(rd_data[11]));
 BUF_X1 output15 (.A(net15),
    .Z(rd_data[12]));
 BUF_X1 output16 (.A(net16),
    .Z(rd_data[13]));
 BUF_X1 output17 (.A(net17),
    .Z(rd_data[14]));
 BUF_X1 output18 (.A(net18),
    .Z(rd_data[15]));
 BUF_X1 output19 (.A(net19),
    .Z(rd_data[16]));
 BUF_X1 output20 (.A(net20),
    .Z(rd_data[17]));
 BUF_X1 output21 (.A(net21),
    .Z(rd_data[18]));
 BUF_X1 output22 (.A(net22),
    .Z(rd_data[19]));
 BUF_X1 output23 (.A(net23),
    .Z(rd_data[1]));
 BUF_X1 output24 (.A(net24),
    .Z(rd_data[20]));
 BUF_X1 output25 (.A(net25),
    .Z(rd_data[21]));
 BUF_X1 output26 (.A(net26),
    .Z(rd_data[22]));
 BUF_X1 output27 (.A(net27),
    .Z(rd_data[23]));
 BUF_X1 output28 (.A(net28),
    .Z(rd_data[24]));
 BUF_X1 output29 (.A(net29),
    .Z(rd_data[25]));
 BUF_X1 output30 (.A(net30),
    .Z(rd_data[26]));
 BUF_X1 output31 (.A(net31),
    .Z(rd_data[27]));
 BUF_X1 output32 (.A(net32),
    .Z(rd_data[28]));
 BUF_X1 output33 (.A(net33),
    .Z(rd_data[29]));
 BUF_X1 output34 (.A(net34),
    .Z(rd_data[2]));
 BUF_X1 output35 (.A(net35),
    .Z(rd_data[30]));
 BUF_X1 output36 (.A(net36),
    .Z(rd_data[31]));
 BUF_X1 output37 (.A(net37),
    .Z(rd_data[3]));
 BUF_X1 output38 (.A(net38),
    .Z(rd_data[4]));
 BUF_X1 output39 (.A(net39),
    .Z(rd_data[5]));
 BUF_X1 output40 (.A(net40),
    .Z(rd_data[6]));
 BUF_X1 output41 (.A(net41),
    .Z(rd_data[7]));
 BUF_X1 output42 (.A(net42),
    .Z(rd_data[8]));
 BUF_X1 output43 (.A(net43),
    .Z(rd_data[9]));
 BUF_X1 output44 (.A(net44),
    .Z(rd_empty));
 BUF_X1 output45 (.A(net45),
    .Z(wr_almost_full));
 BUF_X1 output46 (.A(net46),
    .Z(wr_count[0]));
 BUF_X1 output47 (.A(net47),
    .Z(wr_count[1]));
 BUF_X1 output48 (.A(net48),
    .Z(wr_count[2]));
 BUF_X1 output49 (.A(net49),
    .Z(wr_count[3]));
 BUF_X1 output50 (.A(net50),
    .Z(wr_count[4]));
 BUF_X1 output51 (.A(net51),
    .Z(wr_full));
 CLKBUF_X3 clkbuf_leaf_0_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_0_wr_clk));
 CLKBUF_X3 clkbuf_leaf_1_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_1_wr_clk));
 CLKBUF_X3 clkbuf_leaf_2_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_2_wr_clk));
 CLKBUF_X3 clkbuf_leaf_3_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_3_wr_clk));
 CLKBUF_X3 clkbuf_leaf_4_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_4_wr_clk));
 CLKBUF_X3 clkbuf_leaf_5_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_5_wr_clk));
 CLKBUF_X3 clkbuf_leaf_6_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_6_wr_clk));
 CLKBUF_X3 clkbuf_leaf_7_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_7_wr_clk));
 CLKBUF_X3 clkbuf_leaf_8_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_8_wr_clk));
 CLKBUF_X3 clkbuf_leaf_9_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_9_wr_clk));
 CLKBUF_X3 clkbuf_leaf_10_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_10_wr_clk));
 CLKBUF_X3 clkbuf_leaf_11_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_11_wr_clk));
 CLKBUF_X3 clkbuf_leaf_12_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_12_wr_clk));
 CLKBUF_X3 clkbuf_leaf_13_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_13_wr_clk));
 CLKBUF_X3 clkbuf_leaf_14_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_14_wr_clk));
 CLKBUF_X3 clkbuf_leaf_15_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_15_wr_clk));
 CLKBUF_X3 clkbuf_leaf_16_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_16_wr_clk));
 CLKBUF_X3 clkbuf_leaf_17_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_17_wr_clk));
 CLKBUF_X3 clkbuf_leaf_18_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_18_wr_clk));
 CLKBUF_X3 clkbuf_leaf_19_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_19_wr_clk));
 CLKBUF_X3 clkbuf_leaf_20_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_20_wr_clk));
 CLKBUF_X3 clkbuf_leaf_21_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_21_wr_clk));
 CLKBUF_X3 clkbuf_leaf_22_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_22_wr_clk));
 CLKBUF_X3 clkbuf_leaf_23_wr_clk (.A(clknet_3_5__leaf_wr_clk),
    .Z(clknet_leaf_23_wr_clk));
 CLKBUF_X3 clkbuf_leaf_24_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_24_wr_clk));
 CLKBUF_X3 clkbuf_leaf_25_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_25_wr_clk));
 CLKBUF_X3 clkbuf_leaf_26_wr_clk (.A(clknet_3_4__leaf_wr_clk),
    .Z(clknet_leaf_26_wr_clk));
 CLKBUF_X3 clkbuf_leaf_27_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_27_wr_clk));
 CLKBUF_X3 clkbuf_leaf_28_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_28_wr_clk));
 CLKBUF_X3 clkbuf_leaf_29_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_29_wr_clk));
 CLKBUF_X3 clkbuf_leaf_30_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_30_wr_clk));
 CLKBUF_X3 clkbuf_leaf_31_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_31_wr_clk));
 CLKBUF_X3 clkbuf_leaf_32_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_32_wr_clk));
 CLKBUF_X3 clkbuf_leaf_33_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_33_wr_clk));
 CLKBUF_X3 clkbuf_leaf_34_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_34_wr_clk));
 CLKBUF_X3 clkbuf_leaf_35_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_35_wr_clk));
 CLKBUF_X3 clkbuf_leaf_36_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_36_wr_clk));
 CLKBUF_X3 clkbuf_leaf_37_wr_clk (.A(clknet_3_7__leaf_wr_clk),
    .Z(clknet_leaf_37_wr_clk));
 CLKBUF_X3 clkbuf_leaf_38_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_38_wr_clk));
 CLKBUF_X3 clkbuf_leaf_39_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_39_wr_clk));
 CLKBUF_X3 clkbuf_leaf_40_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_40_wr_clk));
 CLKBUF_X3 clkbuf_leaf_41_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_41_wr_clk));
 CLKBUF_X3 clkbuf_leaf_42_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_42_wr_clk));
 CLKBUF_X3 clkbuf_leaf_43_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_43_wr_clk));
 CLKBUF_X3 clkbuf_leaf_44_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_44_wr_clk));
 CLKBUF_X3 clkbuf_leaf_45_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_45_wr_clk));
 CLKBUF_X3 clkbuf_leaf_46_wr_clk (.A(clknet_3_6__leaf_wr_clk),
    .Z(clknet_leaf_46_wr_clk));
 CLKBUF_X3 clkbuf_leaf_47_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_47_wr_clk));
 CLKBUF_X3 clkbuf_leaf_48_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_48_wr_clk));
 CLKBUF_X3 clkbuf_leaf_49_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_49_wr_clk));
 CLKBUF_X3 clkbuf_leaf_50_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_50_wr_clk));
 CLKBUF_X3 clkbuf_leaf_51_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_51_wr_clk));
 CLKBUF_X3 clkbuf_leaf_52_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_52_wr_clk));
 CLKBUF_X3 clkbuf_leaf_53_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_53_wr_clk));
 CLKBUF_X3 clkbuf_leaf_54_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_54_wr_clk));
 CLKBUF_X3 clkbuf_leaf_55_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_55_wr_clk));
 CLKBUF_X3 clkbuf_leaf_56_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_56_wr_clk));
 CLKBUF_X3 clkbuf_leaf_57_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_57_wr_clk));
 CLKBUF_X3 clkbuf_leaf_58_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_58_wr_clk));
 CLKBUF_X3 clkbuf_leaf_59_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_59_wr_clk));
 CLKBUF_X3 clkbuf_leaf_60_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_60_wr_clk));
 CLKBUF_X3 clkbuf_leaf_61_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_61_wr_clk));
 CLKBUF_X3 clkbuf_leaf_62_wr_clk (.A(clknet_3_3__leaf_wr_clk),
    .Z(clknet_leaf_62_wr_clk));
 CLKBUF_X3 clkbuf_leaf_63_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_63_wr_clk));
 CLKBUF_X3 clkbuf_leaf_64_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_64_wr_clk));
 CLKBUF_X3 clkbuf_leaf_65_wr_clk (.A(clknet_3_2__leaf_wr_clk),
    .Z(clknet_leaf_65_wr_clk));
 CLKBUF_X3 clkbuf_leaf_66_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_66_wr_clk));
 CLKBUF_X3 clkbuf_leaf_67_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_67_wr_clk));
 CLKBUF_X3 clkbuf_leaf_68_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_68_wr_clk));
 CLKBUF_X3 clkbuf_leaf_69_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_69_wr_clk));
 CLKBUF_X3 clkbuf_leaf_70_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_70_wr_clk));
 CLKBUF_X3 clkbuf_leaf_71_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_71_wr_clk));
 CLKBUF_X3 clkbuf_leaf_72_wr_clk (.A(clknet_3_0__leaf_wr_clk),
    .Z(clknet_leaf_72_wr_clk));
 CLKBUF_X3 clkbuf_leaf_73_wr_clk (.A(clknet_3_1__leaf_wr_clk),
    .Z(clknet_leaf_73_wr_clk));
 CLKBUF_X3 clkbuf_0_wr_clk (.A(wr_clk),
    .Z(clknet_0_wr_clk));
 CLKBUF_X3 clkbuf_3_0__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_0__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_1__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_1__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_2__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_2__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_3__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_3__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_4__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_4__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_5__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_5__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_6__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_6__leaf_wr_clk));
 CLKBUF_X3 clkbuf_3_7__f_wr_clk (.A(clknet_0_wr_clk),
    .Z(clknet_3_7__leaf_wr_clk));
 INV_X2 clkload0 (.A(clknet_3_0__leaf_wr_clk));
 INV_X2 clkload1 (.A(clknet_3_2__leaf_wr_clk));
 CLKBUF_X3 clkload2 (.A(clknet_3_3__leaf_wr_clk));
 CLKBUF_X3 clkload3 (.A(clknet_3_5__leaf_wr_clk));
 CLKBUF_X1 clkload4 (.A(clknet_leaf_64_wr_clk));
 CLKBUF_X1 clkload5 (.A(clknet_leaf_67_wr_clk));
 CLKBUF_X1 clkload6 (.A(clknet_leaf_68_wr_clk));
 CLKBUF_X1 clkload7 (.A(clknet_leaf_69_wr_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_70_wr_clk));
 CLKBUF_X1 clkload9 (.A(clknet_leaf_72_wr_clk));
 CLKBUF_X1 clkload10 (.A(clknet_leaf_1_wr_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_3_wr_clk));
 INV_X1 clkload12 (.A(clknet_leaf_4_wr_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_5_wr_clk));
 INV_X1 clkload14 (.A(clknet_leaf_7_wr_clk));
 INV_X2 clkload15 (.A(clknet_leaf_73_wr_clk));
 INV_X1 clkload16 (.A(clknet_leaf_53_wr_clk));
 INV_X1 clkload17 (.A(clknet_leaf_55_wr_clk));
 INV_X1 clkload18 (.A(clknet_leaf_56_wr_clk));
 INV_X1 clkload19 (.A(clknet_leaf_57_wr_clk));
 CLKBUF_X2 clkload20 (.A(clknet_leaf_58_wr_clk));
 CLKBUF_X2 clkload21 (.A(clknet_leaf_59_wr_clk));
 CLKBUF_X2 clkload22 (.A(clknet_leaf_65_wr_clk));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_47_wr_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_48_wr_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_49_wr_clk));
 INV_X2 clkload26 (.A(clknet_leaf_52_wr_clk));
 CLKBUF_X1 clkload27 (.A(clknet_leaf_61_wr_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_62_wr_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_8_wr_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_9_wr_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_10_wr_clk));
 INV_X1 clkload32 (.A(clknet_leaf_11_wr_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_12_wr_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_13_wr_clk));
 INV_X2 clkload35 (.A(clknet_leaf_24_wr_clk));
 INV_X1 clkload36 (.A(clknet_leaf_25_wr_clk));
 INV_X2 clkload37 (.A(clknet_leaf_26_wr_clk));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_15_wr_clk));
 INV_X1 clkload39 (.A(clknet_leaf_16_wr_clk));
 INV_X1 clkload40 (.A(clknet_leaf_17_wr_clk));
 INV_X1 clkload41 (.A(clknet_leaf_18_wr_clk));
 CLKBUF_X1 clkload42 (.A(clknet_leaf_19_wr_clk));
 CLKBUF_X1 clkload43 (.A(clknet_leaf_20_wr_clk));
 INV_X1 clkload44 (.A(clknet_leaf_21_wr_clk));
 CLKBUF_X1 clkload45 (.A(clknet_leaf_22_wr_clk));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_38_wr_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_39_wr_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_41_wr_clk));
 CLKBUF_X1 clkload49 (.A(clknet_leaf_42_wr_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_43_wr_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_44_wr_clk));
 INV_X1 clkload52 (.A(clknet_leaf_45_wr_clk));
 INV_X1 clkload53 (.A(clknet_leaf_46_wr_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_29_wr_clk));
 CLKBUF_X1 clkload55 (.A(clknet_leaf_30_wr_clk));
 INV_X1 clkload56 (.A(clknet_leaf_32_wr_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_33_wr_clk));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_34_wr_clk));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_36_wr_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_37_wr_clk));
 CLKBUF_X1 hold1 (.A(net54),
    .Z(net52));
 CLKBUF_X1 hold2 (.A(net56),
    .Z(net53));
 CLKBUF_X1 hold3 (.A(wr_rst_n),
    .Z(net54));
 CLKBUF_X1 hold4 (.A(net52),
    .Z(net55));
 CLKBUF_X1 hold5 (.A(net5),
    .Z(net56));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X1 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_133 ();
 FILLCELL_X32 FILLER_0_144 ();
 FILLCELL_X16 FILLER_0_182 ();
 FILLCELL_X2 FILLER_0_198 ();
 FILLCELL_X1 FILLER_0_200 ();
 FILLCELL_X8 FILLER_0_204 ();
 FILLCELL_X4 FILLER_0_212 ();
 FILLCELL_X1 FILLER_0_216 ();
 FILLCELL_X8 FILLER_0_220 ();
 FILLCELL_X4 FILLER_0_228 ();
 FILLCELL_X1 FILLER_0_232 ();
 FILLCELL_X4 FILLER_0_236 ();
 FILLCELL_X2 FILLER_0_240 ();
 FILLCELL_X8 FILLER_0_245 ();
 FILLCELL_X4 FILLER_0_253 ();
 FILLCELL_X2 FILLER_0_257 ();
 FILLCELL_X8 FILLER_0_262 ();
 FILLCELL_X1 FILLER_0_270 ();
 FILLCELL_X2 FILLER_0_278 ();
 FILLCELL_X8 FILLER_0_283 ();
 FILLCELL_X4 FILLER_0_291 ();
 FILLCELL_X1 FILLER_0_295 ();
 FILLCELL_X32 FILLER_0_299 ();
 FILLCELL_X2 FILLER_0_331 ();
 FILLCELL_X16 FILLER_0_355 ();
 FILLCELL_X8 FILLER_0_371 ();
 FILLCELL_X4 FILLER_0_379 ();
 FILLCELL_X2 FILLER_0_383 ();
 FILLCELL_X1 FILLER_0_385 ();
 FILLCELL_X16 FILLER_0_389 ();
 FILLCELL_X1 FILLER_0_431 ();
 FILLCELL_X32 FILLER_0_442 ();
 FILLCELL_X32 FILLER_0_474 ();
 FILLCELL_X8 FILLER_0_506 ();
 FILLCELL_X2 FILLER_0_514 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_133 ();
 FILLCELL_X8 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_169 ();
 FILLCELL_X2 FILLER_1_188 ();
 FILLCELL_X1 FILLER_1_190 ();
 FILLCELL_X4 FILLER_1_198 ();
 FILLCELL_X1 FILLER_1_202 ();
 FILLCELL_X2 FILLER_1_224 ();
 FILLCELL_X1 FILLER_1_226 ();
 FILLCELL_X4 FILLER_1_244 ();
 FILLCELL_X1 FILLER_1_248 ();
 FILLCELL_X2 FILLER_1_266 ();
 FILLCELL_X32 FILLER_1_275 ();
 FILLCELL_X32 FILLER_1_307 ();
 FILLCELL_X2 FILLER_1_339 ();
 FILLCELL_X2 FILLER_1_373 ();
 FILLCELL_X1 FILLER_1_375 ();
 FILLCELL_X2 FILLER_1_387 ();
 FILLCELL_X1 FILLER_1_399 ();
 FILLCELL_X2 FILLER_1_434 ();
 FILLCELL_X1 FILLER_1_436 ();
 FILLCELL_X32 FILLER_1_457 ();
 FILLCELL_X16 FILLER_1_489 ();
 FILLCELL_X8 FILLER_1_505 ();
 FILLCELL_X2 FILLER_1_513 ();
 FILLCELL_X1 FILLER_1_515 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X8 FILLER_2_129 ();
 FILLCELL_X8 FILLER_2_154 ();
 FILLCELL_X2 FILLER_2_186 ();
 FILLCELL_X1 FILLER_2_188 ();
 FILLCELL_X8 FILLER_2_237 ();
 FILLCELL_X2 FILLER_2_245 ();
 FILLCELL_X1 FILLER_2_247 ();
 FILLCELL_X32 FILLER_2_282 ();
 FILLCELL_X16 FILLER_2_314 ();
 FILLCELL_X4 FILLER_2_330 ();
 FILLCELL_X2 FILLER_2_350 ();
 FILLCELL_X2 FILLER_2_386 ();
 FILLCELL_X1 FILLER_2_388 ();
 FILLCELL_X1 FILLER_2_435 ();
 FILLCELL_X32 FILLER_2_456 ();
 FILLCELL_X16 FILLER_2_488 ();
 FILLCELL_X8 FILLER_2_504 ();
 FILLCELL_X4 FILLER_2_512 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_129 ();
 FILLCELL_X1 FILLER_3_133 ();
 FILLCELL_X2 FILLER_3_141 ();
 FILLCELL_X4 FILLER_3_150 ();
 FILLCELL_X4 FILLER_3_168 ();
 FILLCELL_X2 FILLER_3_179 ();
 FILLCELL_X1 FILLER_3_181 ();
 FILLCELL_X16 FILLER_3_196 ();
 FILLCELL_X4 FILLER_3_212 ();
 FILLCELL_X1 FILLER_3_216 ();
 FILLCELL_X2 FILLER_3_224 ();
 FILLCELL_X2 FILLER_3_240 ();
 FILLCELL_X2 FILLER_3_245 ();
 FILLCELL_X1 FILLER_3_247 ();
 FILLCELL_X1 FILLER_3_255 ();
 FILLCELL_X2 FILLER_3_263 ();
 FILLCELL_X1 FILLER_3_265 ();
 FILLCELL_X8 FILLER_3_280 ();
 FILLCELL_X4 FILLER_3_288 ();
 FILLCELL_X4 FILLER_3_326 ();
 FILLCELL_X2 FILLER_3_330 ();
 FILLCELL_X1 FILLER_3_349 ();
 FILLCELL_X8 FILLER_3_385 ();
 FILLCELL_X4 FILLER_3_393 ();
 FILLCELL_X2 FILLER_3_397 ();
 FILLCELL_X1 FILLER_3_429 ();
 FILLCELL_X16 FILLER_3_432 ();
 FILLCELL_X4 FILLER_3_448 ();
 FILLCELL_X32 FILLER_3_457 ();
 FILLCELL_X16 FILLER_3_489 ();
 FILLCELL_X8 FILLER_3_505 ();
 FILLCELL_X2 FILLER_3_513 ();
 FILLCELL_X1 FILLER_3_515 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X16 FILLER_4_97 ();
 FILLCELL_X1 FILLER_4_113 ();
 FILLCELL_X8 FILLER_4_134 ();
 FILLCELL_X2 FILLER_4_142 ();
 FILLCELL_X8 FILLER_4_161 ();
 FILLCELL_X16 FILLER_4_177 ();
 FILLCELL_X2 FILLER_4_197 ();
 FILLCELL_X8 FILLER_4_202 ();
 FILLCELL_X4 FILLER_4_210 ();
 FILLCELL_X2 FILLER_4_214 ();
 FILLCELL_X16 FILLER_4_256 ();
 FILLCELL_X2 FILLER_4_292 ();
 FILLCELL_X8 FILLER_4_301 ();
 FILLCELL_X4 FILLER_4_333 ();
 FILLCELL_X2 FILLER_4_337 ();
 FILLCELL_X4 FILLER_4_349 ();
 FILLCELL_X2 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_372 ();
 FILLCELL_X1 FILLER_4_404 ();
 FILLCELL_X2 FILLER_4_417 ();
 FILLCELL_X16 FILLER_4_429 ();
 FILLCELL_X1 FILLER_4_445 ();
 FILLCELL_X32 FILLER_4_468 ();
 FILLCELL_X16 FILLER_4_500 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X16 FILLER_5_97 ();
 FILLCELL_X2 FILLER_5_113 ();
 FILLCELL_X1 FILLER_5_115 ();
 FILLCELL_X16 FILLER_5_139 ();
 FILLCELL_X2 FILLER_5_155 ();
 FILLCELL_X8 FILLER_5_180 ();
 FILLCELL_X1 FILLER_5_208 ();
 FILLCELL_X2 FILLER_5_238 ();
 FILLCELL_X1 FILLER_5_240 ();
 FILLCELL_X8 FILLER_5_245 ();
 FILLCELL_X4 FILLER_5_253 ();
 FILLCELL_X1 FILLER_5_257 ();
 FILLCELL_X4 FILLER_5_272 ();
 FILLCELL_X2 FILLER_5_276 ();
 FILLCELL_X16 FILLER_5_285 ();
 FILLCELL_X4 FILLER_5_301 ();
 FILLCELL_X1 FILLER_5_305 ();
 FILLCELL_X2 FILLER_5_313 ();
 FILLCELL_X4 FILLER_5_329 ();
 FILLCELL_X1 FILLER_5_333 ();
 FILLCELL_X4 FILLER_5_349 ();
 FILLCELL_X1 FILLER_5_359 ();
 FILLCELL_X1 FILLER_5_366 ();
 FILLCELL_X2 FILLER_5_376 ();
 FILLCELL_X1 FILLER_5_378 ();
 FILLCELL_X8 FILLER_5_407 ();
 FILLCELL_X4 FILLER_5_415 ();
 FILLCELL_X4 FILLER_5_429 ();
 FILLCELL_X1 FILLER_5_433 ();
 FILLCELL_X32 FILLER_5_454 ();
 FILLCELL_X16 FILLER_5_486 ();
 FILLCELL_X8 FILLER_5_502 ();
 FILLCELL_X4 FILLER_5_510 ();
 FILLCELL_X2 FILLER_5_514 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X16 FILLER_6_97 ();
 FILLCELL_X2 FILLER_6_113 ();
 FILLCELL_X1 FILLER_6_115 ();
 FILLCELL_X4 FILLER_6_120 ();
 FILLCELL_X8 FILLER_6_131 ();
 FILLCELL_X1 FILLER_6_139 ();
 FILLCELL_X1 FILLER_6_151 ();
 FILLCELL_X1 FILLER_6_169 ();
 FILLCELL_X1 FILLER_6_174 ();
 FILLCELL_X2 FILLER_6_179 ();
 FILLCELL_X8 FILLER_6_198 ();
 FILLCELL_X4 FILLER_6_206 ();
 FILLCELL_X2 FILLER_6_210 ();
 FILLCELL_X4 FILLER_6_219 ();
 FILLCELL_X1 FILLER_6_223 ();
 FILLCELL_X32 FILLER_6_228 ();
 FILLCELL_X1 FILLER_6_274 ();
 FILLCELL_X16 FILLER_6_280 ();
 FILLCELL_X4 FILLER_6_296 ();
 FILLCELL_X2 FILLER_6_300 ();
 FILLCELL_X1 FILLER_6_311 ();
 FILLCELL_X2 FILLER_6_321 ();
 FILLCELL_X1 FILLER_6_342 ();
 FILLCELL_X2 FILLER_6_360 ();
 FILLCELL_X16 FILLER_6_390 ();
 FILLCELL_X4 FILLER_6_406 ();
 FILLCELL_X32 FILLER_6_469 ();
 FILLCELL_X8 FILLER_6_501 ();
 FILLCELL_X4 FILLER_6_509 ();
 FILLCELL_X2 FILLER_6_513 ();
 FILLCELL_X1 FILLER_6_515 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_17 ();
 FILLCELL_X4 FILLER_7_25 ();
 FILLCELL_X8 FILLER_7_46 ();
 FILLCELL_X2 FILLER_7_54 ();
 FILLCELL_X8 FILLER_7_83 ();
 FILLCELL_X2 FILLER_7_91 ();
 FILLCELL_X32 FILLER_7_110 ();
 FILLCELL_X1 FILLER_7_142 ();
 FILLCELL_X16 FILLER_7_160 ();
 FILLCELL_X8 FILLER_7_176 ();
 FILLCELL_X2 FILLER_7_184 ();
 FILLCELL_X16 FILLER_7_197 ();
 FILLCELL_X4 FILLER_7_213 ();
 FILLCELL_X2 FILLER_7_217 ();
 FILLCELL_X1 FILLER_7_219 ();
 FILLCELL_X16 FILLER_7_224 ();
 FILLCELL_X4 FILLER_7_240 ();
 FILLCELL_X1 FILLER_7_244 ();
 FILLCELL_X1 FILLER_7_262 ();
 FILLCELL_X16 FILLER_7_277 ();
 FILLCELL_X8 FILLER_7_293 ();
 FILLCELL_X2 FILLER_7_301 ();
 FILLCELL_X1 FILLER_7_330 ();
 FILLCELL_X1 FILLER_7_337 ();
 FILLCELL_X2 FILLER_7_351 ();
 FILLCELL_X1 FILLER_7_362 ();
 FILLCELL_X2 FILLER_7_373 ();
 FILLCELL_X1 FILLER_7_387 ();
 FILLCELL_X4 FILLER_7_400 ();
 FILLCELL_X4 FILLER_7_426 ();
 FILLCELL_X1 FILLER_7_430 ();
 FILLCELL_X32 FILLER_7_451 ();
 FILLCELL_X32 FILLER_7_483 ();
 FILLCELL_X1 FILLER_7_515 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_20 ();
 FILLCELL_X2 FILLER_8_28 ();
 FILLCELL_X1 FILLER_8_30 ();
 FILLCELL_X1 FILLER_8_55 ();
 FILLCELL_X1 FILLER_8_80 ();
 FILLCELL_X32 FILLER_8_105 ();
 FILLCELL_X2 FILLER_8_137 ();
 FILLCELL_X2 FILLER_8_146 ();
 FILLCELL_X1 FILLER_8_148 ();
 FILLCELL_X4 FILLER_8_166 ();
 FILLCELL_X1 FILLER_8_170 ();
 FILLCELL_X4 FILLER_8_199 ();
 FILLCELL_X8 FILLER_8_234 ();
 FILLCELL_X2 FILLER_8_242 ();
 FILLCELL_X4 FILLER_8_261 ();
 FILLCELL_X2 FILLER_8_265 ();
 FILLCELL_X1 FILLER_8_267 ();
 FILLCELL_X16 FILLER_8_285 ();
 FILLCELL_X4 FILLER_8_301 ();
 FILLCELL_X2 FILLER_8_305 ();
 FILLCELL_X1 FILLER_8_316 ();
 FILLCELL_X2 FILLER_8_326 ();
 FILLCELL_X2 FILLER_8_337 ();
 FILLCELL_X4 FILLER_8_352 ();
 FILLCELL_X1 FILLER_8_356 ();
 FILLCELL_X8 FILLER_8_366 ();
 FILLCELL_X4 FILLER_8_374 ();
 FILLCELL_X1 FILLER_8_378 ();
 FILLCELL_X8 FILLER_8_382 ();
 FILLCELL_X2 FILLER_8_390 ();
 FILLCELL_X16 FILLER_8_412 ();
 FILLCELL_X1 FILLER_8_428 ();
 FILLCELL_X1 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_470 ();
 FILLCELL_X8 FILLER_8_502 ();
 FILLCELL_X4 FILLER_8_510 ();
 FILLCELL_X2 FILLER_8_514 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_33 ();
 FILLCELL_X1 FILLER_9_41 ();
 FILLCELL_X2 FILLER_9_49 ();
 FILLCELL_X1 FILLER_9_84 ();
 FILLCELL_X8 FILLER_9_116 ();
 FILLCELL_X2 FILLER_9_124 ();
 FILLCELL_X1 FILLER_9_126 ();
 FILLCELL_X2 FILLER_9_144 ();
 FILLCELL_X1 FILLER_9_146 ();
 FILLCELL_X1 FILLER_9_154 ();
 FILLCELL_X1 FILLER_9_184 ();
 FILLCELL_X8 FILLER_9_202 ();
 FILLCELL_X4 FILLER_9_234 ();
 FILLCELL_X2 FILLER_9_238 ();
 FILLCELL_X1 FILLER_9_240 ();
 FILLCELL_X2 FILLER_9_262 ();
 FILLCELL_X8 FILLER_9_291 ();
 FILLCELL_X1 FILLER_9_299 ();
 FILLCELL_X4 FILLER_9_307 ();
 FILLCELL_X2 FILLER_9_311 ();
 FILLCELL_X1 FILLER_9_313 ();
 FILLCELL_X4 FILLER_9_321 ();
 FILLCELL_X2 FILLER_9_325 ();
 FILLCELL_X8 FILLER_9_331 ();
 FILLCELL_X4 FILLER_9_339 ();
 FILLCELL_X2 FILLER_9_343 ();
 FILLCELL_X1 FILLER_9_345 ();
 FILLCELL_X4 FILLER_9_359 ();
 FILLCELL_X1 FILLER_9_363 ();
 FILLCELL_X4 FILLER_9_378 ();
 FILLCELL_X2 FILLER_9_382 ();
 FILLCELL_X2 FILLER_9_411 ();
 FILLCELL_X1 FILLER_9_413 ();
 FILLCELL_X32 FILLER_9_434 ();
 FILLCELL_X32 FILLER_9_466 ();
 FILLCELL_X16 FILLER_9_498 ();
 FILLCELL_X2 FILLER_9_514 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_9 ();
 FILLCELL_X32 FILLER_10_14 ();
 FILLCELL_X32 FILLER_10_46 ();
 FILLCELL_X8 FILLER_10_78 ();
 FILLCELL_X4 FILLER_10_86 ();
 FILLCELL_X2 FILLER_10_90 ();
 FILLCELL_X1 FILLER_10_92 ();
 FILLCELL_X8 FILLER_10_100 ();
 FILLCELL_X2 FILLER_10_132 ();
 FILLCELL_X8 FILLER_10_141 ();
 FILLCELL_X2 FILLER_10_149 ();
 FILLCELL_X2 FILLER_10_153 ();
 FILLCELL_X16 FILLER_10_158 ();
 FILLCELL_X8 FILLER_10_174 ();
 FILLCELL_X4 FILLER_10_182 ();
 FILLCELL_X2 FILLER_10_186 ();
 FILLCELL_X8 FILLER_10_197 ();
 FILLCELL_X4 FILLER_10_205 ();
 FILLCELL_X2 FILLER_10_226 ();
 FILLCELL_X4 FILLER_10_230 ();
 FILLCELL_X2 FILLER_10_234 ();
 FILLCELL_X8 FILLER_10_250 ();
 FILLCELL_X4 FILLER_10_258 ();
 FILLCELL_X1 FILLER_10_262 ();
 FILLCELL_X4 FILLER_10_267 ();
 FILLCELL_X2 FILLER_10_271 ();
 FILLCELL_X8 FILLER_10_282 ();
 FILLCELL_X4 FILLER_10_290 ();
 FILLCELL_X2 FILLER_10_294 ();
 FILLCELL_X8 FILLER_10_347 ();
 FILLCELL_X2 FILLER_10_355 ();
 FILLCELL_X4 FILLER_10_364 ();
 FILLCELL_X8 FILLER_10_408 ();
 FILLCELL_X4 FILLER_10_416 ();
 FILLCELL_X2 FILLER_10_420 ();
 FILLCELL_X1 FILLER_10_422 ();
 FILLCELL_X2 FILLER_10_443 ();
 FILLCELL_X1 FILLER_10_445 ();
 FILLCELL_X16 FILLER_10_466 ();
 FILLCELL_X8 FILLER_10_482 ();
 FILLCELL_X8 FILLER_10_503 ();
 FILLCELL_X4 FILLER_10_511 ();
 FILLCELL_X1 FILLER_10_515 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X2 FILLER_11_13 ();
 FILLCELL_X32 FILLER_11_39 ();
 FILLCELL_X8 FILLER_11_71 ();
 FILLCELL_X4 FILLER_11_79 ();
 FILLCELL_X2 FILLER_11_83 ();
 FILLCELL_X1 FILLER_11_85 ();
 FILLCELL_X16 FILLER_11_113 ();
 FILLCELL_X8 FILLER_11_129 ();
 FILLCELL_X1 FILLER_11_161 ();
 FILLCELL_X2 FILLER_11_166 ();
 FILLCELL_X1 FILLER_11_168 ();
 FILLCELL_X4 FILLER_11_174 ();
 FILLCELL_X2 FILLER_11_178 ();
 FILLCELL_X1 FILLER_11_180 ();
 FILLCELL_X4 FILLER_11_185 ();
 FILLCELL_X2 FILLER_11_193 ();
 FILLCELL_X1 FILLER_11_195 ();
 FILLCELL_X4 FILLER_11_200 ();
 FILLCELL_X2 FILLER_11_204 ();
 FILLCELL_X1 FILLER_11_206 ();
 FILLCELL_X2 FILLER_11_214 ();
 FILLCELL_X1 FILLER_11_216 ();
 FILLCELL_X4 FILLER_11_222 ();
 FILLCELL_X2 FILLER_11_226 ();
 FILLCELL_X1 FILLER_11_228 ();
 FILLCELL_X8 FILLER_11_233 ();
 FILLCELL_X2 FILLER_11_241 ();
 FILLCELL_X4 FILLER_11_250 ();
 FILLCELL_X4 FILLER_11_263 ();
 FILLCELL_X2 FILLER_11_267 ();
 FILLCELL_X1 FILLER_11_280 ();
 FILLCELL_X16 FILLER_11_285 ();
 FILLCELL_X1 FILLER_11_325 ();
 FILLCELL_X16 FILLER_11_335 ();
 FILLCELL_X2 FILLER_11_351 ();
 FILLCELL_X1 FILLER_11_353 ();
 FILLCELL_X8 FILLER_11_366 ();
 FILLCELL_X2 FILLER_11_374 ();
 FILLCELL_X1 FILLER_11_396 ();
 FILLCELL_X16 FILLER_11_417 ();
 FILLCELL_X4 FILLER_11_433 ();
 FILLCELL_X1 FILLER_11_437 ();
 FILLCELL_X4 FILLER_11_458 ();
 FILLCELL_X1 FILLER_11_462 ();
 FILLCELL_X8 FILLER_11_478 ();
 FILLCELL_X4 FILLER_11_486 ();
 FILLCELL_X1 FILLER_11_490 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X1 FILLER_12_13 ();
 FILLCELL_X8 FILLER_12_38 ();
 FILLCELL_X2 FILLER_12_46 ();
 FILLCELL_X2 FILLER_12_55 ();
 FILLCELL_X2 FILLER_12_81 ();
 FILLCELL_X4 FILLER_12_100 ();
 FILLCELL_X8 FILLER_12_137 ();
 FILLCELL_X4 FILLER_12_145 ();
 FILLCELL_X2 FILLER_12_149 ();
 FILLCELL_X2 FILLER_12_180 ();
 FILLCELL_X1 FILLER_12_182 ();
 FILLCELL_X1 FILLER_12_201 ();
 FILLCELL_X1 FILLER_12_219 ();
 FILLCELL_X8 FILLER_12_231 ();
 FILLCELL_X1 FILLER_12_239 ();
 FILLCELL_X16 FILLER_12_292 ();
 FILLCELL_X4 FILLER_12_308 ();
 FILLCELL_X4 FILLER_12_316 ();
 FILLCELL_X2 FILLER_12_320 ();
 FILLCELL_X1 FILLER_12_322 ();
 FILLCELL_X1 FILLER_12_332 ();
 FILLCELL_X16 FILLER_12_374 ();
 FILLCELL_X2 FILLER_12_390 ();
 FILLCELL_X8 FILLER_12_412 ();
 FILLCELL_X4 FILLER_12_420 ();
 FILLCELL_X2 FILLER_12_424 ();
 FILLCELL_X4 FILLER_12_453 ();
 FILLCELL_X1 FILLER_12_457 ();
 FILLCELL_X4 FILLER_12_464 ();
 FILLCELL_X2 FILLER_12_468 ();
 FILLCELL_X32 FILLER_12_480 ();
 FILLCELL_X4 FILLER_12_512 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_19 ();
 FILLCELL_X1 FILLER_13_27 ();
 FILLCELL_X4 FILLER_13_56 ();
 FILLCELL_X1 FILLER_13_60 ();
 FILLCELL_X2 FILLER_13_92 ();
 FILLCELL_X4 FILLER_13_106 ();
 FILLCELL_X2 FILLER_13_110 ();
 FILLCELL_X4 FILLER_13_115 ();
 FILLCELL_X16 FILLER_13_143 ();
 FILLCELL_X2 FILLER_13_159 ();
 FILLCELL_X2 FILLER_13_173 ();
 FILLCELL_X2 FILLER_13_188 ();
 FILLCELL_X4 FILLER_13_193 ();
 FILLCELL_X1 FILLER_13_197 ();
 FILLCELL_X4 FILLER_13_201 ();
 FILLCELL_X2 FILLER_13_205 ();
 FILLCELL_X1 FILLER_13_207 ();
 FILLCELL_X2 FILLER_13_235 ();
 FILLCELL_X8 FILLER_13_244 ();
 FILLCELL_X4 FILLER_13_252 ();
 FILLCELL_X2 FILLER_13_263 ();
 FILLCELL_X4 FILLER_13_280 ();
 FILLCELL_X2 FILLER_13_284 ();
 FILLCELL_X1 FILLER_13_286 ();
 FILLCELL_X16 FILLER_13_304 ();
 FILLCELL_X2 FILLER_13_320 ();
 FILLCELL_X1 FILLER_13_355 ();
 FILLCELL_X16 FILLER_13_362 ();
 FILLCELL_X2 FILLER_13_378 ();
 FILLCELL_X8 FILLER_13_407 ();
 FILLCELL_X16 FILLER_13_435 ();
 FILLCELL_X2 FILLER_13_451 ();
 FILLCELL_X2 FILLER_13_467 ();
 FILLCELL_X1 FILLER_13_469 ();
 FILLCELL_X1 FILLER_13_483 ();
 FILLCELL_X16 FILLER_13_491 ();
 FILLCELL_X8 FILLER_13_507 ();
 FILLCELL_X1 FILLER_13_515 ();
 FILLCELL_X1 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_26 ();
 FILLCELL_X1 FILLER_14_52 ();
 FILLCELL_X4 FILLER_14_60 ();
 FILLCELL_X2 FILLER_14_64 ();
 FILLCELL_X2 FILLER_14_73 ();
 FILLCELL_X4 FILLER_14_85 ();
 FILLCELL_X2 FILLER_14_89 ();
 FILLCELL_X1 FILLER_14_97 ();
 FILLCELL_X1 FILLER_14_121 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X4 FILLER_14_161 ();
 FILLCELL_X2 FILLER_14_165 ();
 FILLCELL_X1 FILLER_14_167 ();
 FILLCELL_X1 FILLER_14_171 ();
 FILLCELL_X16 FILLER_14_189 ();
 FILLCELL_X8 FILLER_14_205 ();
 FILLCELL_X4 FILLER_14_227 ();
 FILLCELL_X1 FILLER_14_240 ();
 FILLCELL_X16 FILLER_14_258 ();
 FILLCELL_X4 FILLER_14_274 ();
 FILLCELL_X2 FILLER_14_278 ();
 FILLCELL_X1 FILLER_14_280 ();
 FILLCELL_X1 FILLER_14_290 ();
 FILLCELL_X4 FILLER_14_298 ();
 FILLCELL_X2 FILLER_14_302 ();
 FILLCELL_X1 FILLER_14_304 ();
 FILLCELL_X1 FILLER_14_312 ();
 FILLCELL_X8 FILLER_14_318 ();
 FILLCELL_X1 FILLER_14_343 ();
 FILLCELL_X2 FILLER_14_353 ();
 FILLCELL_X4 FILLER_14_362 ();
 FILLCELL_X2 FILLER_14_366 ();
 FILLCELL_X1 FILLER_14_368 ();
 FILLCELL_X32 FILLER_14_376 ();
 FILLCELL_X2 FILLER_14_408 ();
 FILLCELL_X1 FILLER_14_410 ();
 FILLCELL_X16 FILLER_14_431 ();
 FILLCELL_X4 FILLER_14_447 ();
 FILLCELL_X2 FILLER_14_451 ();
 FILLCELL_X1 FILLER_14_453 ();
 FILLCELL_X4 FILLER_14_475 ();
 FILLCELL_X2 FILLER_14_479 ();
 FILLCELL_X8 FILLER_14_502 ();
 FILLCELL_X4 FILLER_14_510 ();
 FILLCELL_X2 FILLER_14_514 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_25 ();
 FILLCELL_X32 FILLER_15_31 ();
 FILLCELL_X8 FILLER_15_63 ();
 FILLCELL_X2 FILLER_15_71 ();
 FILLCELL_X1 FILLER_15_73 ();
 FILLCELL_X32 FILLER_15_96 ();
 FILLCELL_X8 FILLER_15_128 ();
 FILLCELL_X4 FILLER_15_143 ();
 FILLCELL_X2 FILLER_15_147 ();
 FILLCELL_X1 FILLER_15_149 ();
 FILLCELL_X8 FILLER_15_184 ();
 FILLCELL_X2 FILLER_15_192 ();
 FILLCELL_X1 FILLER_15_194 ();
 FILLCELL_X8 FILLER_15_226 ();
 FILLCELL_X2 FILLER_15_234 ();
 FILLCELL_X8 FILLER_15_243 ();
 FILLCELL_X8 FILLER_15_275 ();
 FILLCELL_X4 FILLER_15_283 ();
 FILLCELL_X2 FILLER_15_287 ();
 FILLCELL_X1 FILLER_15_338 ();
 FILLCELL_X16 FILLER_15_348 ();
 FILLCELL_X8 FILLER_15_364 ();
 FILLCELL_X4 FILLER_15_372 ();
 FILLCELL_X2 FILLER_15_376 ();
 FILLCELL_X8 FILLER_15_385 ();
 FILLCELL_X2 FILLER_15_393 ();
 FILLCELL_X8 FILLER_15_422 ();
 FILLCELL_X4 FILLER_15_430 ();
 FILLCELL_X2 FILLER_15_434 ();
 FILLCELL_X1 FILLER_15_436 ();
 FILLCELL_X8 FILLER_15_457 ();
 FILLCELL_X1 FILLER_15_465 ();
 FILLCELL_X1 FILLER_15_476 ();
 FILLCELL_X1 FILLER_15_489 ();
 FILLCELL_X8 FILLER_15_496 ();
 FILLCELL_X8 FILLER_15_507 ();
 FILLCELL_X1 FILLER_15_515 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_5 ();
 FILLCELL_X1 FILLER_16_7 ();
 FILLCELL_X4 FILLER_16_32 ();
 FILLCELL_X1 FILLER_16_36 ();
 FILLCELL_X2 FILLER_16_61 ();
 FILLCELL_X2 FILLER_16_70 ();
 FILLCELL_X2 FILLER_16_87 ();
 FILLCELL_X1 FILLER_16_89 ();
 FILLCELL_X1 FILLER_16_107 ();
 FILLCELL_X2 FILLER_16_111 ();
 FILLCELL_X4 FILLER_16_130 ();
 FILLCELL_X2 FILLER_16_134 ();
 FILLCELL_X2 FILLER_16_153 ();
 FILLCELL_X4 FILLER_16_190 ();
 FILLCELL_X2 FILLER_16_194 ();
 FILLCELL_X4 FILLER_16_227 ();
 FILLCELL_X2 FILLER_16_231 ();
 FILLCELL_X1 FILLER_16_257 ();
 FILLCELL_X2 FILLER_16_275 ();
 FILLCELL_X8 FILLER_16_294 ();
 FILLCELL_X8 FILLER_16_319 ();
 FILLCELL_X1 FILLER_16_327 ();
 FILLCELL_X4 FILLER_16_355 ();
 FILLCELL_X16 FILLER_16_366 ();
 FILLCELL_X2 FILLER_16_382 ();
 FILLCELL_X1 FILLER_16_396 ();
 FILLCELL_X16 FILLER_16_408 ();
 FILLCELL_X2 FILLER_16_424 ();
 FILLCELL_X1 FILLER_16_426 ();
 FILLCELL_X4 FILLER_16_433 ();
 FILLCELL_X1 FILLER_16_437 ();
 FILLCELL_X8 FILLER_16_452 ();
 FILLCELL_X4 FILLER_16_460 ();
 FILLCELL_X2 FILLER_16_464 ();
 FILLCELL_X1 FILLER_16_466 ();
 FILLCELL_X2 FILLER_16_479 ();
 FILLCELL_X4 FILLER_16_487 ();
 FILLCELL_X2 FILLER_16_495 ();
 FILLCELL_X1 FILLER_16_511 ();
 FILLCELL_X1 FILLER_16_515 ();
 FILLCELL_X2 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_3 ();
 FILLCELL_X2 FILLER_17_7 ();
 FILLCELL_X4 FILLER_17_54 ();
 FILLCELL_X2 FILLER_17_75 ();
 FILLCELL_X1 FILLER_17_77 ();
 FILLCELL_X2 FILLER_17_107 ();
 FILLCELL_X8 FILLER_17_136 ();
 FILLCELL_X4 FILLER_17_144 ();
 FILLCELL_X2 FILLER_17_148 ();
 FILLCELL_X1 FILLER_17_155 ();
 FILLCELL_X2 FILLER_17_170 ();
 FILLCELL_X8 FILLER_17_189 ();
 FILLCELL_X4 FILLER_17_197 ();
 FILLCELL_X2 FILLER_17_201 ();
 FILLCELL_X8 FILLER_17_210 ();
 FILLCELL_X16 FILLER_17_235 ();
 FILLCELL_X2 FILLER_17_272 ();
 FILLCELL_X8 FILLER_17_293 ();
 FILLCELL_X2 FILLER_17_301 ();
 FILLCELL_X1 FILLER_17_303 ();
 FILLCELL_X2 FILLER_17_311 ();
 FILLCELL_X1 FILLER_17_313 ();
 FILLCELL_X1 FILLER_17_335 ();
 FILLCELL_X2 FILLER_17_379 ();
 FILLCELL_X16 FILLER_17_403 ();
 FILLCELL_X4 FILLER_17_419 ();
 FILLCELL_X2 FILLER_17_443 ();
 FILLCELL_X1 FILLER_17_445 ();
 FILLCELL_X2 FILLER_17_466 ();
 FILLCELL_X1 FILLER_17_477 ();
 FILLCELL_X8 FILLER_17_490 ();
 FILLCELL_X2 FILLER_17_498 ();
 FILLCELL_X1 FILLER_17_500 ();
 FILLCELL_X2 FILLER_17_514 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_5 ();
 FILLCELL_X16 FILLER_18_27 ();
 FILLCELL_X4 FILLER_18_43 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X8 FILLER_18_72 ();
 FILLCELL_X4 FILLER_18_87 ();
 FILLCELL_X1 FILLER_18_103 ();
 FILLCELL_X1 FILLER_18_108 ();
 FILLCELL_X1 FILLER_18_120 ();
 FILLCELL_X16 FILLER_18_124 ();
 FILLCELL_X8 FILLER_18_140 ();
 FILLCELL_X2 FILLER_18_148 ();
 FILLCELL_X1 FILLER_18_150 ();
 FILLCELL_X2 FILLER_18_158 ();
 FILLCELL_X1 FILLER_18_160 ();
 FILLCELL_X32 FILLER_18_168 ();
 FILLCELL_X4 FILLER_18_200 ();
 FILLCELL_X8 FILLER_18_221 ();
 FILLCELL_X1 FILLER_18_229 ();
 FILLCELL_X32 FILLER_18_237 ();
 FILLCELL_X8 FILLER_18_286 ();
 FILLCELL_X1 FILLER_18_294 ();
 FILLCELL_X8 FILLER_18_313 ();
 FILLCELL_X2 FILLER_18_321 ();
 FILLCELL_X16 FILLER_18_368 ();
 FILLCELL_X4 FILLER_18_387 ();
 FILLCELL_X2 FILLER_18_418 ();
 FILLCELL_X8 FILLER_18_455 ();
 FILLCELL_X4 FILLER_18_463 ();
 FILLCELL_X1 FILLER_18_467 ();
 FILLCELL_X4 FILLER_18_494 ();
 FILLCELL_X2 FILLER_18_498 ();
 FILLCELL_X2 FILLER_18_507 ();
 FILLCELL_X1 FILLER_18_509 ();
 FILLCELL_X2 FILLER_18_513 ();
 FILLCELL_X1 FILLER_18_515 ();
 FILLCELL_X32 FILLER_19_4 ();
 FILLCELL_X32 FILLER_19_36 ();
 FILLCELL_X16 FILLER_19_68 ();
 FILLCELL_X8 FILLER_19_84 ();
 FILLCELL_X2 FILLER_19_92 ();
 FILLCELL_X32 FILLER_19_98 ();
 FILLCELL_X16 FILLER_19_130 ();
 FILLCELL_X2 FILLER_19_146 ();
 FILLCELL_X4 FILLER_19_155 ();
 FILLCELL_X2 FILLER_19_176 ();
 FILLCELL_X8 FILLER_19_195 ();
 FILLCELL_X2 FILLER_19_227 ();
 FILLCELL_X1 FILLER_19_229 ();
 FILLCELL_X32 FILLER_19_259 ();
 FILLCELL_X4 FILLER_19_291 ();
 FILLCELL_X2 FILLER_19_295 ();
 FILLCELL_X1 FILLER_19_297 ();
 FILLCELL_X2 FILLER_19_303 ();
 FILLCELL_X4 FILLER_19_322 ();
 FILLCELL_X4 FILLER_19_336 ();
 FILLCELL_X32 FILLER_19_349 ();
 FILLCELL_X8 FILLER_19_381 ();
 FILLCELL_X16 FILLER_19_396 ();
 FILLCELL_X1 FILLER_19_412 ();
 FILLCELL_X4 FILLER_19_443 ();
 FILLCELL_X16 FILLER_19_457 ();
 FILLCELL_X2 FILLER_19_473 ();
 FILLCELL_X1 FILLER_19_475 ();
 FILLCELL_X16 FILLER_19_492 ();
 FILLCELL_X8 FILLER_19_508 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_27 ();
 FILLCELL_X1 FILLER_20_31 ();
 FILLCELL_X4 FILLER_20_60 ();
 FILLCELL_X2 FILLER_20_64 ();
 FILLCELL_X1 FILLER_20_66 ();
 FILLCELL_X2 FILLER_20_74 ();
 FILLCELL_X2 FILLER_20_108 ();
 FILLCELL_X1 FILLER_20_110 ();
 FILLCELL_X16 FILLER_20_118 ();
 FILLCELL_X8 FILLER_20_134 ();
 FILLCELL_X2 FILLER_20_142 ();
 FILLCELL_X4 FILLER_20_175 ();
 FILLCELL_X4 FILLER_20_186 ();
 FILLCELL_X2 FILLER_20_190 ();
 FILLCELL_X8 FILLER_20_199 ();
 FILLCELL_X2 FILLER_20_207 ();
 FILLCELL_X1 FILLER_20_209 ();
 FILLCELL_X4 FILLER_20_217 ();
 FILLCELL_X1 FILLER_20_221 ();
 FILLCELL_X8 FILLER_20_227 ();
 FILLCELL_X2 FILLER_20_235 ();
 FILLCELL_X1 FILLER_20_237 ();
 FILLCELL_X4 FILLER_20_266 ();
 FILLCELL_X2 FILLER_20_270 ();
 FILLCELL_X1 FILLER_20_272 ();
 FILLCELL_X2 FILLER_20_307 ();
 FILLCELL_X1 FILLER_20_309 ();
 FILLCELL_X4 FILLER_20_315 ();
 FILLCELL_X2 FILLER_20_319 ();
 FILLCELL_X1 FILLER_20_321 ();
 FILLCELL_X4 FILLER_20_346 ();
 FILLCELL_X1 FILLER_20_350 ();
 FILLCELL_X8 FILLER_20_382 ();
 FILLCELL_X4 FILLER_20_390 ();
 FILLCELL_X1 FILLER_20_394 ();
 FILLCELL_X2 FILLER_20_402 ();
 FILLCELL_X1 FILLER_20_404 ();
 FILLCELL_X16 FILLER_20_412 ();
 FILLCELL_X4 FILLER_20_428 ();
 FILLCELL_X2 FILLER_20_432 ();
 FILLCELL_X1 FILLER_20_434 ();
 FILLCELL_X32 FILLER_20_479 ();
 FILLCELL_X4 FILLER_20_511 ();
 FILLCELL_X1 FILLER_20_515 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_5 ();
 FILLCELL_X2 FILLER_21_52 ();
 FILLCELL_X1 FILLER_21_54 ();
 FILLCELL_X2 FILLER_21_111 ();
 FILLCELL_X1 FILLER_21_113 ();
 FILLCELL_X16 FILLER_21_131 ();
 FILLCELL_X1 FILLER_21_147 ();
 FILLCELL_X2 FILLER_21_203 ();
 FILLCELL_X1 FILLER_21_205 ();
 FILLCELL_X32 FILLER_21_227 ();
 FILLCELL_X8 FILLER_21_259 ();
 FILLCELL_X4 FILLER_21_267 ();
 FILLCELL_X2 FILLER_21_271 ();
 FILLCELL_X4 FILLER_21_306 ();
 FILLCELL_X2 FILLER_21_332 ();
 FILLCELL_X1 FILLER_21_334 ();
 FILLCELL_X4 FILLER_21_342 ();
 FILLCELL_X1 FILLER_21_346 ();
 FILLCELL_X1 FILLER_21_352 ();
 FILLCELL_X4 FILLER_21_370 ();
 FILLCELL_X2 FILLER_21_374 ();
 FILLCELL_X4 FILLER_21_383 ();
 FILLCELL_X1 FILLER_21_387 ();
 FILLCELL_X16 FILLER_21_395 ();
 FILLCELL_X2 FILLER_21_411 ();
 FILLCELL_X8 FILLER_21_430 ();
 FILLCELL_X4 FILLER_21_438 ();
 FILLCELL_X1 FILLER_21_442 ();
 FILLCELL_X1 FILLER_21_460 ();
 FILLCELL_X32 FILLER_21_471 ();
 FILLCELL_X8 FILLER_21_503 ();
 FILLCELL_X4 FILLER_21_511 ();
 FILLCELL_X1 FILLER_21_515 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_5 ();
 FILLCELL_X8 FILLER_22_13 ();
 FILLCELL_X1 FILLER_22_21 ();
 FILLCELL_X2 FILLER_22_39 ();
 FILLCELL_X1 FILLER_22_41 ();
 FILLCELL_X2 FILLER_22_47 ();
 FILLCELL_X4 FILLER_22_66 ();
 FILLCELL_X2 FILLER_22_70 ();
 FILLCELL_X1 FILLER_22_72 ();
 FILLCELL_X2 FILLER_22_92 ();
 FILLCELL_X8 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_114 ();
 FILLCELL_X8 FILLER_22_135 ();
 FILLCELL_X4 FILLER_22_143 ();
 FILLCELL_X2 FILLER_22_147 ();
 FILLCELL_X16 FILLER_22_154 ();
 FILLCELL_X4 FILLER_22_170 ();
 FILLCELL_X2 FILLER_22_174 ();
 FILLCELL_X4 FILLER_22_200 ();
 FILLCELL_X2 FILLER_22_211 ();
 FILLCELL_X4 FILLER_22_225 ();
 FILLCELL_X2 FILLER_22_229 ();
 FILLCELL_X1 FILLER_22_231 ();
 FILLCELL_X8 FILLER_22_247 ();
 FILLCELL_X2 FILLER_22_255 ();
 FILLCELL_X2 FILLER_22_262 ();
 FILLCELL_X16 FILLER_22_271 ();
 FILLCELL_X1 FILLER_22_298 ();
 FILLCELL_X4 FILLER_22_303 ();
 FILLCELL_X2 FILLER_22_307 ();
 FILLCELL_X1 FILLER_22_309 ();
 FILLCELL_X4 FILLER_22_319 ();
 FILLCELL_X2 FILLER_22_323 ();
 FILLCELL_X2 FILLER_22_353 ();
 FILLCELL_X1 FILLER_22_355 ();
 FILLCELL_X16 FILLER_22_361 ();
 FILLCELL_X8 FILLER_22_377 ();
 FILLCELL_X2 FILLER_22_385 ();
 FILLCELL_X4 FILLER_22_401 ();
 FILLCELL_X2 FILLER_22_405 ();
 FILLCELL_X32 FILLER_22_411 ();
 FILLCELL_X8 FILLER_22_443 ();
 FILLCELL_X1 FILLER_22_451 ();
 FILLCELL_X2 FILLER_22_459 ();
 FILLCELL_X32 FILLER_22_466 ();
 FILLCELL_X16 FILLER_22_498 ();
 FILLCELL_X2 FILLER_22_514 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X8 FILLER_23_17 ();
 FILLCELL_X4 FILLER_23_25 ();
 FILLCELL_X2 FILLER_23_29 ();
 FILLCELL_X4 FILLER_23_34 ();
 FILLCELL_X2 FILLER_23_38 ();
 FILLCELL_X16 FILLER_23_57 ();
 FILLCELL_X4 FILLER_23_73 ();
 FILLCELL_X8 FILLER_23_97 ();
 FILLCELL_X1 FILLER_23_105 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X1 FILLER_23_121 ();
 FILLCELL_X32 FILLER_23_125 ();
 FILLCELL_X16 FILLER_23_157 ();
 FILLCELL_X8 FILLER_23_173 ();
 FILLCELL_X2 FILLER_23_181 ();
 FILLCELL_X1 FILLER_23_183 ();
 FILLCELL_X4 FILLER_23_191 ();
 FILLCELL_X8 FILLER_23_200 ();
 FILLCELL_X8 FILLER_23_232 ();
 FILLCELL_X1 FILLER_23_240 ();
 FILLCELL_X2 FILLER_23_275 ();
 FILLCELL_X4 FILLER_23_289 ();
 FILLCELL_X4 FILLER_23_315 ();
 FILLCELL_X1 FILLER_23_319 ();
 FILLCELL_X8 FILLER_23_324 ();
 FILLCELL_X1 FILLER_23_332 ();
 FILLCELL_X32 FILLER_23_340 ();
 FILLCELL_X2 FILLER_23_389 ();
 FILLCELL_X16 FILLER_23_408 ();
 FILLCELL_X2 FILLER_23_424 ();
 FILLCELL_X2 FILLER_23_433 ();
 FILLCELL_X4 FILLER_23_452 ();
 FILLCELL_X32 FILLER_23_463 ();
 FILLCELL_X16 FILLER_23_495 ();
 FILLCELL_X4 FILLER_23_511 ();
 FILLCELL_X1 FILLER_23_515 ();
 FILLCELL_X4 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_5 ();
 FILLCELL_X1 FILLER_24_7 ();
 FILLCELL_X16 FILLER_24_25 ();
 FILLCELL_X1 FILLER_24_41 ();
 FILLCELL_X2 FILLER_24_49 ();
 FILLCELL_X1 FILLER_24_51 ();
 FILLCELL_X2 FILLER_24_59 ();
 FILLCELL_X2 FILLER_24_68 ();
 FILLCELL_X1 FILLER_24_70 ();
 FILLCELL_X4 FILLER_24_76 ();
 FILLCELL_X1 FILLER_24_80 ();
 FILLCELL_X4 FILLER_24_88 ();
 FILLCELL_X1 FILLER_24_92 ();
 FILLCELL_X4 FILLER_24_97 ();
 FILLCELL_X2 FILLER_24_111 ();
 FILLCELL_X1 FILLER_24_113 ();
 FILLCELL_X2 FILLER_24_118 ();
 FILLCELL_X16 FILLER_24_123 ();
 FILLCELL_X4 FILLER_24_141 ();
 FILLCELL_X1 FILLER_24_145 ();
 FILLCELL_X2 FILLER_24_151 ();
 FILLCELL_X1 FILLER_24_153 ();
 FILLCELL_X1 FILLER_24_175 ();
 FILLCELL_X16 FILLER_24_193 ();
 FILLCELL_X4 FILLER_24_209 ();
 FILLCELL_X8 FILLER_24_227 ();
 FILLCELL_X4 FILLER_24_235 ();
 FILLCELL_X1 FILLER_24_239 ();
 FILLCELL_X8 FILLER_24_247 ();
 FILLCELL_X2 FILLER_24_255 ();
 FILLCELL_X1 FILLER_24_257 ();
 FILLCELL_X8 FILLER_24_265 ();
 FILLCELL_X4 FILLER_24_273 ();
 FILLCELL_X1 FILLER_24_277 ();
 FILLCELL_X16 FILLER_24_295 ();
 FILLCELL_X2 FILLER_24_311 ();
 FILLCELL_X8 FILLER_24_320 ();
 FILLCELL_X1 FILLER_24_328 ();
 FILLCELL_X4 FILLER_24_346 ();
 FILLCELL_X1 FILLER_24_374 ();
 FILLCELL_X4 FILLER_24_382 ();
 FILLCELL_X2 FILLER_24_386 ();
 FILLCELL_X1 FILLER_24_388 ();
 FILLCELL_X8 FILLER_24_421 ();
 FILLCELL_X2 FILLER_24_453 ();
 FILLCELL_X32 FILLER_24_479 ();
 FILLCELL_X4 FILLER_24_511 ();
 FILLCELL_X1 FILLER_24_515 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_9 ();
 FILLCELL_X2 FILLER_25_20 ();
 FILLCELL_X1 FILLER_25_22 ();
 FILLCELL_X4 FILLER_25_30 ();
 FILLCELL_X2 FILLER_25_34 ();
 FILLCELL_X8 FILLER_25_73 ();
 FILLCELL_X4 FILLER_25_81 ();
 FILLCELL_X2 FILLER_25_85 ();
 FILLCELL_X4 FILLER_25_90 ();
 FILLCELL_X1 FILLER_25_94 ();
 FILLCELL_X4 FILLER_25_154 ();
 FILLCELL_X1 FILLER_25_158 ();
 FILLCELL_X32 FILLER_25_176 ();
 FILLCELL_X1 FILLER_25_208 ();
 FILLCELL_X1 FILLER_25_226 ();
 FILLCELL_X2 FILLER_25_234 ();
 FILLCELL_X1 FILLER_25_236 ();
 FILLCELL_X2 FILLER_25_254 ();
 FILLCELL_X8 FILLER_25_273 ();
 FILLCELL_X4 FILLER_25_281 ();
 FILLCELL_X1 FILLER_25_285 ();
 FILLCELL_X8 FILLER_25_313 ();
 FILLCELL_X4 FILLER_25_321 ();
 FILLCELL_X1 FILLER_25_325 ();
 FILLCELL_X2 FILLER_25_333 ();
 FILLCELL_X4 FILLER_25_342 ();
 FILLCELL_X2 FILLER_25_363 ();
 FILLCELL_X4 FILLER_25_393 ();
 FILLCELL_X1 FILLER_25_397 ();
 FILLCELL_X1 FILLER_25_415 ();
 FILLCELL_X2 FILLER_25_423 ();
 FILLCELL_X1 FILLER_25_436 ();
 FILLCELL_X2 FILLER_25_441 ();
 FILLCELL_X1 FILLER_25_443 ();
 FILLCELL_X32 FILLER_25_464 ();
 FILLCELL_X16 FILLER_25_496 ();
 FILLCELL_X4 FILLER_25_512 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_32 ();
 FILLCELL_X1 FILLER_26_34 ();
 FILLCELL_X8 FILLER_26_41 ();
 FILLCELL_X4 FILLER_26_49 ();
 FILLCELL_X4 FILLER_26_60 ();
 FILLCELL_X2 FILLER_26_64 ();
 FILLCELL_X1 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_70 ();
 FILLCELL_X1 FILLER_26_72 ();
 FILLCELL_X8 FILLER_26_80 ();
 FILLCELL_X2 FILLER_26_88 ();
 FILLCELL_X4 FILLER_26_99 ();
 FILLCELL_X16 FILLER_26_110 ();
 FILLCELL_X1 FILLER_26_171 ();
 FILLCELL_X2 FILLER_26_177 ();
 FILLCELL_X1 FILLER_26_179 ();
 FILLCELL_X4 FILLER_26_187 ();
 FILLCELL_X1 FILLER_26_191 ();
 FILLCELL_X2 FILLER_26_209 ();
 FILLCELL_X4 FILLER_26_218 ();
 FILLCELL_X2 FILLER_26_229 ();
 FILLCELL_X2 FILLER_26_238 ();
 FILLCELL_X2 FILLER_26_250 ();
 FILLCELL_X16 FILLER_26_259 ();
 FILLCELL_X4 FILLER_26_275 ();
 FILLCELL_X2 FILLER_26_279 ();
 FILLCELL_X2 FILLER_26_312 ();
 FILLCELL_X1 FILLER_26_314 ();
 FILLCELL_X4 FILLER_26_328 ();
 FILLCELL_X1 FILLER_26_332 ();
 FILLCELL_X1 FILLER_26_340 ();
 FILLCELL_X2 FILLER_26_352 ();
 FILLCELL_X16 FILLER_26_361 ();
 FILLCELL_X8 FILLER_26_377 ();
 FILLCELL_X4 FILLER_26_385 ();
 FILLCELL_X2 FILLER_26_389 ();
 FILLCELL_X1 FILLER_26_391 ();
 FILLCELL_X8 FILLER_26_399 ();
 FILLCELL_X4 FILLER_26_407 ();
 FILLCELL_X2 FILLER_26_411 ();
 FILLCELL_X1 FILLER_26_413 ();
 FILLCELL_X4 FILLER_26_421 ();
 FILLCELL_X2 FILLER_26_425 ();
 FILLCELL_X2 FILLER_26_437 ();
 FILLCELL_X2 FILLER_26_444 ();
 FILLCELL_X32 FILLER_26_474 ();
 FILLCELL_X8 FILLER_26_506 ();
 FILLCELL_X2 FILLER_26_514 ();
 FILLCELL_X8 FILLER_27_1 ();
 FILLCELL_X4 FILLER_27_9 ();
 FILLCELL_X2 FILLER_27_13 ();
 FILLCELL_X1 FILLER_27_15 ();
 FILLCELL_X1 FILLER_27_43 ();
 FILLCELL_X8 FILLER_27_55 ();
 FILLCELL_X2 FILLER_27_63 ();
 FILLCELL_X8 FILLER_27_101 ();
 FILLCELL_X1 FILLER_27_109 ();
 FILLCELL_X2 FILLER_27_119 ();
 FILLCELL_X8 FILLER_27_130 ();
 FILLCELL_X2 FILLER_27_138 ();
 FILLCELL_X1 FILLER_27_140 ();
 FILLCELL_X16 FILLER_27_155 ();
 FILLCELL_X2 FILLER_27_171 ();
 FILLCELL_X1 FILLER_27_173 ();
 FILLCELL_X1 FILLER_27_191 ();
 FILLCELL_X4 FILLER_27_199 ();
 FILLCELL_X2 FILLER_27_203 ();
 FILLCELL_X2 FILLER_27_212 ();
 FILLCELL_X1 FILLER_27_214 ();
 FILLCELL_X2 FILLER_27_249 ();
 FILLCELL_X16 FILLER_27_272 ();
 FILLCELL_X4 FILLER_27_288 ();
 FILLCELL_X1 FILLER_27_292 ();
 FILLCELL_X1 FILLER_27_300 ();
 FILLCELL_X2 FILLER_27_308 ();
 FILLCELL_X1 FILLER_27_317 ();
 FILLCELL_X4 FILLER_27_361 ();
 FILLCELL_X4 FILLER_27_367 ();
 FILLCELL_X2 FILLER_27_371 ();
 FILLCELL_X8 FILLER_27_380 ();
 FILLCELL_X4 FILLER_27_412 ();
 FILLCELL_X2 FILLER_27_416 ();
 FILLCELL_X1 FILLER_27_418 ();
 FILLCELL_X2 FILLER_27_453 ();
 FILLCELL_X1 FILLER_27_455 ();
 FILLCELL_X16 FILLER_27_490 ();
 FILLCELL_X4 FILLER_27_506 ();
 FILLCELL_X2 FILLER_27_510 ();
 FILLCELL_X1 FILLER_27_512 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_17 ();
 FILLCELL_X2 FILLER_28_21 ();
 FILLCELL_X1 FILLER_28_23 ();
 FILLCELL_X8 FILLER_28_31 ();
 FILLCELL_X4 FILLER_28_39 ();
 FILLCELL_X16 FILLER_28_67 ();
 FILLCELL_X4 FILLER_28_83 ();
 FILLCELL_X2 FILLER_28_87 ();
 FILLCELL_X1 FILLER_28_106 ();
 FILLCELL_X4 FILLER_28_124 ();
 FILLCELL_X2 FILLER_28_128 ();
 FILLCELL_X1 FILLER_28_130 ();
 FILLCELL_X8 FILLER_28_155 ();
 FILLCELL_X4 FILLER_28_163 ();
 FILLCELL_X2 FILLER_28_167 ();
 FILLCELL_X1 FILLER_28_169 ();
 FILLCELL_X2 FILLER_28_177 ();
 FILLCELL_X8 FILLER_28_186 ();
 FILLCELL_X2 FILLER_28_216 ();
 FILLCELL_X1 FILLER_28_218 ();
 FILLCELL_X8 FILLER_28_223 ();
 FILLCELL_X4 FILLER_28_231 ();
 FILLCELL_X16 FILLER_28_252 ();
 FILLCELL_X1 FILLER_28_268 ();
 FILLCELL_X2 FILLER_28_273 ();
 FILLCELL_X1 FILLER_28_275 ();
 FILLCELL_X8 FILLER_28_281 ();
 FILLCELL_X2 FILLER_28_289 ();
 FILLCELL_X1 FILLER_28_291 ();
 FILLCELL_X4 FILLER_28_297 ();
 FILLCELL_X2 FILLER_28_301 ();
 FILLCELL_X16 FILLER_28_310 ();
 FILLCELL_X2 FILLER_28_337 ();
 FILLCELL_X1 FILLER_28_339 ();
 FILLCELL_X1 FILLER_28_351 ();
 FILLCELL_X1 FILLER_28_359 ();
 FILLCELL_X1 FILLER_28_381 ();
 FILLCELL_X2 FILLER_28_399 ();
 FILLCELL_X1 FILLER_28_401 ();
 FILLCELL_X4 FILLER_28_419 ();
 FILLCELL_X1 FILLER_28_423 ();
 FILLCELL_X1 FILLER_28_431 ();
 FILLCELL_X2 FILLER_28_443 ();
 FILLCELL_X2 FILLER_28_471 ();
 FILLCELL_X1 FILLER_28_473 ();
 FILLCELL_X8 FILLER_28_481 ();
 FILLCELL_X2 FILLER_28_489 ();
 FILLCELL_X1 FILLER_28_515 ();
 FILLCELL_X1 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_19 ();
 FILLCELL_X1 FILLER_29_27 ();
 FILLCELL_X1 FILLER_29_42 ();
 FILLCELL_X16 FILLER_29_77 ();
 FILLCELL_X4 FILLER_29_93 ();
 FILLCELL_X2 FILLER_29_97 ();
 FILLCELL_X1 FILLER_29_99 ();
 FILLCELL_X8 FILLER_29_155 ();
 FILLCELL_X2 FILLER_29_163 ();
 FILLCELL_X1 FILLER_29_165 ();
 FILLCELL_X1 FILLER_29_190 ();
 FILLCELL_X4 FILLER_29_196 ();
 FILLCELL_X1 FILLER_29_200 ();
 FILLCELL_X4 FILLER_29_205 ();
 FILLCELL_X16 FILLER_29_215 ();
 FILLCELL_X4 FILLER_29_231 ();
 FILLCELL_X2 FILLER_29_235 ();
 FILLCELL_X2 FILLER_29_266 ();
 FILLCELL_X1 FILLER_29_268 ();
 FILLCELL_X2 FILLER_29_283 ();
 FILLCELL_X4 FILLER_29_316 ();
 FILLCELL_X2 FILLER_29_320 ();
 FILLCELL_X1 FILLER_29_322 ();
 FILLCELL_X4 FILLER_29_347 ();
 FILLCELL_X2 FILLER_29_351 ();
 FILLCELL_X4 FILLER_29_379 ();
 FILLCELL_X2 FILLER_29_383 ();
 FILLCELL_X1 FILLER_29_406 ();
 FILLCELL_X1 FILLER_29_436 ();
 FILLCELL_X1 FILLER_29_441 ();
 FILLCELL_X1 FILLER_29_454 ();
 FILLCELL_X2 FILLER_29_462 ();
 FILLCELL_X1 FILLER_29_464 ();
 FILLCELL_X16 FILLER_29_469 ();
 FILLCELL_X4 FILLER_29_485 ();
 FILLCELL_X2 FILLER_29_489 ();
 FILLCELL_X1 FILLER_29_515 ();
 FILLCELL_X2 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_3 ();
 FILLCELL_X8 FILLER_30_28 ();
 FILLCELL_X2 FILLER_30_36 ();
 FILLCELL_X4 FILLER_30_45 ();
 FILLCELL_X1 FILLER_30_49 ();
 FILLCELL_X1 FILLER_30_57 ();
 FILLCELL_X16 FILLER_30_72 ();
 FILLCELL_X8 FILLER_30_88 ();
 FILLCELL_X4 FILLER_30_127 ();
 FILLCELL_X2 FILLER_30_131 ();
 FILLCELL_X16 FILLER_30_147 ();
 FILLCELL_X4 FILLER_30_163 ();
 FILLCELL_X2 FILLER_30_167 ();
 FILLCELL_X1 FILLER_30_169 ();
 FILLCELL_X1 FILLER_30_204 ();
 FILLCELL_X16 FILLER_30_229 ();
 FILLCELL_X2 FILLER_30_245 ();
 FILLCELL_X1 FILLER_30_247 ();
 FILLCELL_X4 FILLER_30_251 ();
 FILLCELL_X2 FILLER_30_255 ();
 FILLCELL_X1 FILLER_30_264 ();
 FILLCELL_X4 FILLER_30_272 ();
 FILLCELL_X1 FILLER_30_276 ();
 FILLCELL_X4 FILLER_30_318 ();
 FILLCELL_X2 FILLER_30_322 ();
 FILLCELL_X1 FILLER_30_324 ();
 FILLCELL_X2 FILLER_30_332 ();
 FILLCELL_X8 FILLER_30_341 ();
 FILLCELL_X2 FILLER_30_349 ();
 FILLCELL_X8 FILLER_30_358 ();
 FILLCELL_X8 FILLER_30_380 ();
 FILLCELL_X4 FILLER_30_388 ();
 FILLCELL_X32 FILLER_30_399 ();
 FILLCELL_X16 FILLER_30_431 ();
 FILLCELL_X4 FILLER_30_447 ();
 FILLCELL_X2 FILLER_30_451 ();
 FILLCELL_X1 FILLER_30_453 ();
 FILLCELL_X2 FILLER_30_466 ();
 FILLCELL_X1 FILLER_30_468 ();
 FILLCELL_X2 FILLER_30_514 ();
 FILLCELL_X8 FILLER_31_1 ();
 FILLCELL_X16 FILLER_31_13 ();
 FILLCELL_X16 FILLER_31_53 ();
 FILLCELL_X2 FILLER_31_69 ();
 FILLCELL_X8 FILLER_31_93 ();
 FILLCELL_X4 FILLER_31_101 ();
 FILLCELL_X1 FILLER_31_105 ();
 FILLCELL_X8 FILLER_31_114 ();
 FILLCELL_X1 FILLER_31_122 ();
 FILLCELL_X8 FILLER_31_140 ();
 FILLCELL_X4 FILLER_31_148 ();
 FILLCELL_X1 FILLER_31_152 ();
 FILLCELL_X16 FILLER_31_161 ();
 FILLCELL_X4 FILLER_31_177 ();
 FILLCELL_X4 FILLER_31_222 ();
 FILLCELL_X2 FILLER_31_226 ();
 FILLCELL_X2 FILLER_31_242 ();
 FILLCELL_X1 FILLER_31_244 ();
 FILLCELL_X8 FILLER_31_252 ();
 FILLCELL_X4 FILLER_31_260 ();
 FILLCELL_X1 FILLER_31_264 ();
 FILLCELL_X16 FILLER_31_272 ();
 FILLCELL_X4 FILLER_31_288 ();
 FILLCELL_X4 FILLER_31_306 ();
 FILLCELL_X2 FILLER_31_310 ();
 FILLCELL_X2 FILLER_31_319 ();
 FILLCELL_X1 FILLER_31_321 ();
 FILLCELL_X4 FILLER_31_325 ();
 FILLCELL_X1 FILLER_31_329 ();
 FILLCELL_X8 FILLER_31_338 ();
 FILLCELL_X4 FILLER_31_346 ();
 FILLCELL_X2 FILLER_31_350 ();
 FILLCELL_X2 FILLER_31_369 ();
 FILLCELL_X2 FILLER_31_375 ();
 FILLCELL_X2 FILLER_31_384 ();
 FILLCELL_X1 FILLER_31_386 ();
 FILLCELL_X8 FILLER_31_404 ();
 FILLCELL_X4 FILLER_31_412 ();
 FILLCELL_X1 FILLER_31_416 ();
 FILLCELL_X4 FILLER_31_439 ();
 FILLCELL_X2 FILLER_31_443 ();
 FILLCELL_X1 FILLER_31_445 ();
 FILLCELL_X4 FILLER_31_464 ();
 FILLCELL_X1 FILLER_31_468 ();
 FILLCELL_X16 FILLER_31_497 ();
 FILLCELL_X2 FILLER_31_513 ();
 FILLCELL_X1 FILLER_31_515 ();
 FILLCELL_X8 FILLER_32_1 ();
 FILLCELL_X4 FILLER_32_9 ();
 FILLCELL_X2 FILLER_32_13 ();
 FILLCELL_X1 FILLER_32_15 ();
 FILLCELL_X8 FILLER_32_30 ();
 FILLCELL_X4 FILLER_32_38 ();
 FILLCELL_X4 FILLER_32_45 ();
 FILLCELL_X2 FILLER_32_49 ();
 FILLCELL_X1 FILLER_32_51 ();
 FILLCELL_X8 FILLER_32_60 ();
 FILLCELL_X2 FILLER_32_68 ();
 FILLCELL_X1 FILLER_32_70 ();
 FILLCELL_X4 FILLER_32_102 ();
 FILLCELL_X16 FILLER_32_115 ();
 FILLCELL_X8 FILLER_32_131 ();
 FILLCELL_X4 FILLER_32_139 ();
 FILLCELL_X1 FILLER_32_143 ();
 FILLCELL_X16 FILLER_32_168 ();
 FILLCELL_X4 FILLER_32_184 ();
 FILLCELL_X16 FILLER_32_195 ();
 FILLCELL_X1 FILLER_32_211 ();
 FILLCELL_X1 FILLER_32_236 ();
 FILLCELL_X2 FILLER_32_244 ();
 FILLCELL_X8 FILLER_32_253 ();
 FILLCELL_X1 FILLER_32_261 ();
 FILLCELL_X4 FILLER_32_269 ();
 FILLCELL_X2 FILLER_32_273 ();
 FILLCELL_X1 FILLER_32_275 ();
 FILLCELL_X2 FILLER_32_283 ();
 FILLCELL_X1 FILLER_32_285 ();
 FILLCELL_X16 FILLER_32_305 ();
 FILLCELL_X2 FILLER_32_321 ();
 FILLCELL_X1 FILLER_32_323 ();
 FILLCELL_X4 FILLER_32_331 ();
 FILLCELL_X2 FILLER_32_335 ();
 FILLCELL_X2 FILLER_32_344 ();
 FILLCELL_X1 FILLER_32_346 ();
 FILLCELL_X2 FILLER_32_361 ();
 FILLCELL_X1 FILLER_32_363 ();
 FILLCELL_X2 FILLER_32_398 ();
 FILLCELL_X1 FILLER_32_400 ();
 FILLCELL_X8 FILLER_32_406 ();
 FILLCELL_X2 FILLER_32_414 ();
 FILLCELL_X1 FILLER_32_416 ();
 FILLCELL_X4 FILLER_32_424 ();
 FILLCELL_X8 FILLER_32_442 ();
 FILLCELL_X32 FILLER_32_474 ();
 FILLCELL_X8 FILLER_32_506 ();
 FILLCELL_X2 FILLER_32_514 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X2 FILLER_33_5 ();
 FILLCELL_X2 FILLER_33_38 ();
 FILLCELL_X1 FILLER_33_40 ();
 FILLCELL_X4 FILLER_33_48 ();
 FILLCELL_X2 FILLER_33_52 ();
 FILLCELL_X4 FILLER_33_78 ();
 FILLCELL_X1 FILLER_33_96 ();
 FILLCELL_X1 FILLER_33_104 ();
 FILLCELL_X4 FILLER_33_133 ();
 FILLCELL_X2 FILLER_33_137 ();
 FILLCELL_X1 FILLER_33_139 ();
 FILLCELL_X1 FILLER_33_174 ();
 FILLCELL_X32 FILLER_33_182 ();
 FILLCELL_X16 FILLER_33_214 ();
 FILLCELL_X4 FILLER_33_230 ();
 FILLCELL_X1 FILLER_33_234 ();
 FILLCELL_X8 FILLER_33_249 ();
 FILLCELL_X1 FILLER_33_257 ();
 FILLCELL_X2 FILLER_33_265 ();
 FILLCELL_X4 FILLER_33_274 ();
 FILLCELL_X2 FILLER_33_278 ();
 FILLCELL_X1 FILLER_33_299 ();
 FILLCELL_X2 FILLER_33_321 ();
 FILLCELL_X16 FILLER_33_330 ();
 FILLCELL_X4 FILLER_33_346 ();
 FILLCELL_X2 FILLER_33_350 ();
 FILLCELL_X32 FILLER_33_376 ();
 FILLCELL_X8 FILLER_33_408 ();
 FILLCELL_X2 FILLER_33_416 ();
 FILLCELL_X2 FILLER_33_435 ();
 FILLCELL_X32 FILLER_33_454 ();
 FILLCELL_X16 FILLER_33_486 ();
 FILLCELL_X8 FILLER_33_502 ();
 FILLCELL_X4 FILLER_33_510 ();
 FILLCELL_X2 FILLER_33_514 ();
 FILLCELL_X16 FILLER_34_1 ();
 FILLCELL_X16 FILLER_34_45 ();
 FILLCELL_X4 FILLER_34_68 ();
 FILLCELL_X2 FILLER_34_72 ();
 FILLCELL_X4 FILLER_34_81 ();
 FILLCELL_X2 FILLER_34_85 ();
 FILLCELL_X4 FILLER_34_92 ();
 FILLCELL_X1 FILLER_34_96 ();
 FILLCELL_X8 FILLER_34_131 ();
 FILLCELL_X1 FILLER_34_139 ();
 FILLCELL_X4 FILLER_34_158 ();
 FILLCELL_X2 FILLER_34_219 ();
 FILLCELL_X4 FILLER_34_235 ();
 FILLCELL_X2 FILLER_34_239 ();
 FILLCELL_X2 FILLER_34_248 ();
 FILLCELL_X4 FILLER_34_257 ();
 FILLCELL_X8 FILLER_34_275 ();
 FILLCELL_X2 FILLER_34_283 ();
 FILLCELL_X4 FILLER_34_306 ();
 FILLCELL_X2 FILLER_34_310 ();
 FILLCELL_X1 FILLER_34_312 ();
 FILLCELL_X4 FILLER_34_320 ();
 FILLCELL_X8 FILLER_34_348 ();
 FILLCELL_X2 FILLER_34_356 ();
 FILLCELL_X8 FILLER_34_389 ();
 FILLCELL_X2 FILLER_34_397 ();
 FILLCELL_X1 FILLER_34_399 ();
 FILLCELL_X4 FILLER_34_424 ();
 FILLCELL_X2 FILLER_34_428 ();
 FILLCELL_X32 FILLER_34_437 ();
 FILLCELL_X32 FILLER_34_469 ();
 FILLCELL_X8 FILLER_34_501 ();
 FILLCELL_X4 FILLER_34_509 ();
 FILLCELL_X2 FILLER_34_513 ();
 FILLCELL_X1 FILLER_34_515 ();
 FILLCELL_X16 FILLER_35_1 ();
 FILLCELL_X8 FILLER_35_17 ();
 FILLCELL_X4 FILLER_35_25 ();
 FILLCELL_X1 FILLER_35_29 ();
 FILLCELL_X2 FILLER_35_47 ();
 FILLCELL_X1 FILLER_35_80 ();
 FILLCELL_X32 FILLER_35_119 ();
 FILLCELL_X16 FILLER_35_151 ();
 FILLCELL_X4 FILLER_35_167 ();
 FILLCELL_X2 FILLER_35_171 ();
 FILLCELL_X2 FILLER_35_184 ();
 FILLCELL_X1 FILLER_35_186 ();
 FILLCELL_X8 FILLER_35_238 ();
 FILLCELL_X4 FILLER_35_251 ();
 FILLCELL_X1 FILLER_35_255 ();
 FILLCELL_X8 FILLER_35_263 ();
 FILLCELL_X4 FILLER_35_271 ();
 FILLCELL_X4 FILLER_35_282 ();
 FILLCELL_X2 FILLER_35_286 ();
 FILLCELL_X1 FILLER_35_288 ();
 FILLCELL_X4 FILLER_35_341 ();
 FILLCELL_X1 FILLER_35_345 ();
 FILLCELL_X2 FILLER_35_353 ();
 FILLCELL_X4 FILLER_35_389 ();
 FILLCELL_X2 FILLER_35_393 ();
 FILLCELL_X1 FILLER_35_395 ();
 FILLCELL_X4 FILLER_35_420 ();
 FILLCELL_X2 FILLER_35_424 ();
 FILLCELL_X1 FILLER_35_426 ();
 FILLCELL_X8 FILLER_35_434 ();
 FILLCELL_X2 FILLER_35_442 ();
 FILLCELL_X2 FILLER_35_465 ();
 FILLCELL_X32 FILLER_35_484 ();
 FILLCELL_X8 FILLER_36_1 ();
 FILLCELL_X4 FILLER_36_9 ();
 FILLCELL_X2 FILLER_36_13 ();
 FILLCELL_X1 FILLER_36_15 ();
 FILLCELL_X1 FILLER_36_37 ();
 FILLCELL_X16 FILLER_36_42 ();
 FILLCELL_X8 FILLER_36_58 ();
 FILLCELL_X4 FILLER_36_66 ();
 FILLCELL_X2 FILLER_36_70 ();
 FILLCELL_X4 FILLER_36_79 ();
 FILLCELL_X1 FILLER_36_83 ();
 FILLCELL_X4 FILLER_36_101 ();
 FILLCELL_X2 FILLER_36_105 ();
 FILLCELL_X8 FILLER_36_114 ();
 FILLCELL_X4 FILLER_36_122 ();
 FILLCELL_X4 FILLER_36_133 ();
 FILLCELL_X2 FILLER_36_137 ();
 FILLCELL_X8 FILLER_36_156 ();
 FILLCELL_X4 FILLER_36_164 ();
 FILLCELL_X4 FILLER_36_185 ();
 FILLCELL_X2 FILLER_36_189 ();
 FILLCELL_X2 FILLER_36_205 ();
 FILLCELL_X32 FILLER_36_230 ();
 FILLCELL_X4 FILLER_36_262 ();
 FILLCELL_X2 FILLER_36_266 ();
 FILLCELL_X2 FILLER_36_285 ();
 FILLCELL_X16 FILLER_36_301 ();
 FILLCELL_X4 FILLER_36_317 ();
 FILLCELL_X2 FILLER_36_328 ();
 FILLCELL_X1 FILLER_36_330 ();
 FILLCELL_X2 FILLER_36_340 ();
 FILLCELL_X1 FILLER_36_342 ();
 FILLCELL_X4 FILLER_36_362 ();
 FILLCELL_X2 FILLER_36_366 ();
 FILLCELL_X1 FILLER_36_368 ();
 FILLCELL_X8 FILLER_36_390 ();
 FILLCELL_X4 FILLER_36_398 ();
 FILLCELL_X1 FILLER_36_402 ();
 FILLCELL_X4 FILLER_36_424 ();
 FILLCELL_X1 FILLER_36_428 ();
 FILLCELL_X2 FILLER_36_446 ();
 FILLCELL_X1 FILLER_36_448 ();
 FILLCELL_X2 FILLER_36_456 ();
 FILLCELL_X1 FILLER_36_458 ();
 FILLCELL_X16 FILLER_36_497 ();
 FILLCELL_X2 FILLER_36_513 ();
 FILLCELL_X1 FILLER_36_515 ();
 FILLCELL_X4 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_5 ();
 FILLCELL_X4 FILLER_37_31 ();
 FILLCELL_X2 FILLER_37_35 ();
 FILLCELL_X1 FILLER_37_37 ();
 FILLCELL_X8 FILLER_37_45 ();
 FILLCELL_X2 FILLER_37_53 ();
 FILLCELL_X2 FILLER_37_69 ();
 FILLCELL_X8 FILLER_37_88 ();
 FILLCELL_X4 FILLER_37_96 ();
 FILLCELL_X2 FILLER_37_100 ();
 FILLCELL_X2 FILLER_37_136 ();
 FILLCELL_X2 FILLER_37_145 ();
 FILLCELL_X1 FILLER_37_147 ();
 FILLCELL_X2 FILLER_37_165 ();
 FILLCELL_X1 FILLER_37_167 ();
 FILLCELL_X2 FILLER_37_175 ();
 FILLCELL_X16 FILLER_37_181 ();
 FILLCELL_X8 FILLER_37_197 ();
 FILLCELL_X4 FILLER_37_205 ();
 FILLCELL_X2 FILLER_37_209 ();
 FILLCELL_X1 FILLER_37_211 ();
 FILLCELL_X16 FILLER_37_229 ();
 FILLCELL_X4 FILLER_37_245 ();
 FILLCELL_X1 FILLER_37_249 ();
 FILLCELL_X4 FILLER_37_257 ();
 FILLCELL_X2 FILLER_37_261 ();
 FILLCELL_X1 FILLER_37_263 ();
 FILLCELL_X1 FILLER_37_302 ();
 FILLCELL_X2 FILLER_37_331 ();
 FILLCELL_X16 FILLER_37_344 ();
 FILLCELL_X1 FILLER_37_360 ();
 FILLCELL_X4 FILLER_37_365 ();
 FILLCELL_X2 FILLER_37_378 ();
 FILLCELL_X1 FILLER_37_390 ();
 FILLCELL_X32 FILLER_37_398 ();
 FILLCELL_X8 FILLER_37_430 ();
 FILLCELL_X2 FILLER_37_438 ();
 FILLCELL_X2 FILLER_37_445 ();
 FILLCELL_X1 FILLER_37_447 ();
 FILLCELL_X8 FILLER_37_455 ();
 FILLCELL_X2 FILLER_37_463 ();
 FILLCELL_X1 FILLER_37_465 ();
 FILLCELL_X8 FILLER_37_473 ();
 FILLCELL_X4 FILLER_37_481 ();
 FILLCELL_X2 FILLER_37_497 ();
 FILLCELL_X1 FILLER_37_499 ();
 FILLCELL_X8 FILLER_37_503 ();
 FILLCELL_X4 FILLER_37_511 ();
 FILLCELL_X1 FILLER_37_515 ();
 FILLCELL_X8 FILLER_38_1 ();
 FILLCELL_X2 FILLER_38_9 ();
 FILLCELL_X1 FILLER_38_11 ();
 FILLCELL_X2 FILLER_38_29 ();
 FILLCELL_X1 FILLER_38_31 ();
 FILLCELL_X2 FILLER_38_63 ();
 FILLCELL_X1 FILLER_38_65 ();
 FILLCELL_X8 FILLER_38_90 ();
 FILLCELL_X4 FILLER_38_98 ();
 FILLCELL_X8 FILLER_38_133 ();
 FILLCELL_X4 FILLER_38_141 ();
 FILLCELL_X2 FILLER_38_145 ();
 FILLCELL_X1 FILLER_38_147 ();
 FILLCELL_X2 FILLER_38_157 ();
 FILLCELL_X2 FILLER_38_185 ();
 FILLCELL_X1 FILLER_38_187 ();
 FILLCELL_X8 FILLER_38_191 ();
 FILLCELL_X8 FILLER_38_206 ();
 FILLCELL_X2 FILLER_38_225 ();
 FILLCELL_X4 FILLER_38_231 ();
 FILLCELL_X2 FILLER_38_235 ();
 FILLCELL_X1 FILLER_38_237 ();
 FILLCELL_X8 FILLER_38_259 ();
 FILLCELL_X2 FILLER_38_267 ();
 FILLCELL_X1 FILLER_38_269 ();
 FILLCELL_X4 FILLER_38_287 ();
 FILLCELL_X8 FILLER_38_293 ();
 FILLCELL_X2 FILLER_38_301 ();
 FILLCELL_X8 FILLER_38_310 ();
 FILLCELL_X1 FILLER_38_318 ();
 FILLCELL_X2 FILLER_38_326 ();
 FILLCELL_X1 FILLER_38_345 ();
 FILLCELL_X2 FILLER_38_353 ();
 FILLCELL_X1 FILLER_38_355 ();
 FILLCELL_X4 FILLER_38_363 ();
 FILLCELL_X2 FILLER_38_367 ();
 FILLCELL_X2 FILLER_38_373 ();
 FILLCELL_X1 FILLER_38_375 ();
 FILLCELL_X2 FILLER_38_393 ();
 FILLCELL_X1 FILLER_38_395 ();
 FILLCELL_X1 FILLER_38_415 ();
 FILLCELL_X4 FILLER_38_423 ();
 FILLCELL_X4 FILLER_38_458 ();
 FILLCELL_X1 FILLER_38_462 ();
 FILLCELL_X1 FILLER_38_515 ();
 FILLCELL_X4 FILLER_39_1 ();
 FILLCELL_X4 FILLER_39_29 ();
 FILLCELL_X4 FILLER_39_50 ();
 FILLCELL_X2 FILLER_39_54 ();
 FILLCELL_X1 FILLER_39_56 ();
 FILLCELL_X4 FILLER_39_88 ();
 FILLCELL_X2 FILLER_39_92 ();
 FILLCELL_X1 FILLER_39_94 ();
 FILLCELL_X1 FILLER_39_102 ();
 FILLCELL_X16 FILLER_39_127 ();
 FILLCELL_X4 FILLER_39_143 ();
 FILLCELL_X2 FILLER_39_154 ();
 FILLCELL_X1 FILLER_39_156 ();
 FILLCELL_X4 FILLER_39_188 ();
 FILLCELL_X2 FILLER_39_192 ();
 FILLCELL_X2 FILLER_39_211 ();
 FILLCELL_X1 FILLER_39_213 ();
 FILLCELL_X8 FILLER_39_230 ();
 FILLCELL_X1 FILLER_39_238 ();
 FILLCELL_X4 FILLER_39_263 ();
 FILLCELL_X4 FILLER_39_271 ();
 FILLCELL_X8 FILLER_39_318 ();
 FILLCELL_X4 FILLER_39_343 ();
 FILLCELL_X1 FILLER_39_347 ();
 FILLCELL_X2 FILLER_39_365 ();
 FILLCELL_X1 FILLER_39_367 ();
 FILLCELL_X2 FILLER_39_392 ();
 FILLCELL_X1 FILLER_39_394 ();
 FILLCELL_X4 FILLER_39_468 ();
 FILLCELL_X16 FILLER_39_479 ();
 FILLCELL_X8 FILLER_39_499 ();
 FILLCELL_X4 FILLER_39_507 ();
 FILLCELL_X2 FILLER_39_511 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X8 FILLER_40_17 ();
 FILLCELL_X4 FILLER_40_25 ();
 FILLCELL_X2 FILLER_40_29 ();
 FILLCELL_X32 FILLER_40_39 ();
 FILLCELL_X4 FILLER_40_71 ();
 FILLCELL_X2 FILLER_40_75 ();
 FILLCELL_X4 FILLER_40_94 ();
 FILLCELL_X16 FILLER_40_120 ();
 FILLCELL_X4 FILLER_40_136 ();
 FILLCELL_X2 FILLER_40_178 ();
 FILLCELL_X8 FILLER_40_190 ();
 FILLCELL_X1 FILLER_40_209 ();
 FILLCELL_X2 FILLER_40_215 ();
 FILLCELL_X1 FILLER_40_217 ();
 FILLCELL_X8 FILLER_40_233 ();
 FILLCELL_X1 FILLER_40_244 ();
 FILLCELL_X2 FILLER_40_265 ();
 FILLCELL_X4 FILLER_40_272 ();
 FILLCELL_X2 FILLER_40_276 ();
 FILLCELL_X1 FILLER_40_278 ();
 FILLCELL_X2 FILLER_40_282 ();
 FILLCELL_X1 FILLER_40_284 ();
 FILLCELL_X4 FILLER_40_302 ();
 FILLCELL_X2 FILLER_40_311 ();
 FILLCELL_X8 FILLER_40_330 ();
 FILLCELL_X4 FILLER_40_338 ();
 FILLCELL_X1 FILLER_40_371 ();
 FILLCELL_X16 FILLER_40_377 ();
 FILLCELL_X8 FILLER_40_400 ();
 FILLCELL_X1 FILLER_40_408 ();
 FILLCELL_X4 FILLER_40_417 ();
 FILLCELL_X1 FILLER_40_421 ();
 FILLCELL_X2 FILLER_40_441 ();
 FILLCELL_X1 FILLER_40_443 ();
 FILLCELL_X1 FILLER_40_451 ();
 FILLCELL_X32 FILLER_40_476 ();
 FILLCELL_X8 FILLER_40_508 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X1 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_51 ();
 FILLCELL_X32 FILLER_41_83 ();
 FILLCELL_X8 FILLER_41_115 ();
 FILLCELL_X2 FILLER_41_123 ();
 FILLCELL_X1 FILLER_41_149 ();
 FILLCELL_X2 FILLER_41_195 ();
 FILLCELL_X2 FILLER_41_214 ();
 FILLCELL_X1 FILLER_41_216 ();
 FILLCELL_X1 FILLER_41_234 ();
 FILLCELL_X2 FILLER_41_257 ();
 FILLCELL_X4 FILLER_41_292 ();
 FILLCELL_X4 FILLER_41_303 ();
 FILLCELL_X2 FILLER_41_314 ();
 FILLCELL_X1 FILLER_41_316 ();
 FILLCELL_X8 FILLER_41_324 ();
 FILLCELL_X2 FILLER_41_332 ();
 FILLCELL_X32 FILLER_41_341 ();
 FILLCELL_X16 FILLER_41_373 ();
 FILLCELL_X8 FILLER_41_420 ();
 FILLCELL_X4 FILLER_41_428 ();
 FILLCELL_X1 FILLER_41_432 ();
 FILLCELL_X32 FILLER_41_457 ();
 FILLCELL_X16 FILLER_41_489 ();
 FILLCELL_X8 FILLER_41_505 ();
 FILLCELL_X2 FILLER_41_513 ();
 FILLCELL_X1 FILLER_41_515 ();
 FILLCELL_X8 FILLER_42_1 ();
 FILLCELL_X4 FILLER_42_9 ();
 FILLCELL_X2 FILLER_42_13 ();
 FILLCELL_X8 FILLER_42_19 ();
 FILLCELL_X4 FILLER_42_27 ();
 FILLCELL_X2 FILLER_42_31 ();
 FILLCELL_X1 FILLER_42_33 ();
 FILLCELL_X4 FILLER_42_58 ();
 FILLCELL_X2 FILLER_42_62 ();
 FILLCELL_X1 FILLER_42_64 ();
 FILLCELL_X4 FILLER_42_82 ();
 FILLCELL_X2 FILLER_42_93 ();
 FILLCELL_X8 FILLER_42_112 ();
 FILLCELL_X4 FILLER_42_120 ();
 FILLCELL_X1 FILLER_42_168 ();
 FILLCELL_X32 FILLER_42_177 ();
 FILLCELL_X16 FILLER_42_209 ();
 FILLCELL_X8 FILLER_42_225 ();
 FILLCELL_X8 FILLER_42_247 ();
 FILLCELL_X8 FILLER_42_258 ();
 FILLCELL_X4 FILLER_42_266 ();
 FILLCELL_X2 FILLER_42_270 ();
 FILLCELL_X16 FILLER_42_279 ();
 FILLCELL_X1 FILLER_42_295 ();
 FILLCELL_X8 FILLER_42_313 ();
 FILLCELL_X16 FILLER_42_335 ();
 FILLCELL_X4 FILLER_42_358 ();
 FILLCELL_X4 FILLER_42_386 ();
 FILLCELL_X2 FILLER_42_390 ();
 FILLCELL_X4 FILLER_42_409 ();
 FILLCELL_X2 FILLER_42_413 ();
 FILLCELL_X16 FILLER_42_426 ();
 FILLCELL_X8 FILLER_42_442 ();
 FILLCELL_X4 FILLER_42_450 ();
 FILLCELL_X2 FILLER_42_454 ();
 FILLCELL_X16 FILLER_42_485 ();
 FILLCELL_X8 FILLER_42_501 ();
 FILLCELL_X4 FILLER_42_509 ();
 FILLCELL_X2 FILLER_42_513 ();
 FILLCELL_X1 FILLER_42_515 ();
 FILLCELL_X8 FILLER_43_1 ();
 FILLCELL_X4 FILLER_43_9 ();
 FILLCELL_X2 FILLER_43_13 ();
 FILLCELL_X1 FILLER_43_15 ();
 FILLCELL_X8 FILLER_43_33 ();
 FILLCELL_X4 FILLER_43_41 ();
 FILLCELL_X2 FILLER_43_45 ();
 FILLCELL_X1 FILLER_43_47 ();
 FILLCELL_X16 FILLER_43_58 ();
 FILLCELL_X4 FILLER_43_74 ();
 FILLCELL_X16 FILLER_43_119 ();
 FILLCELL_X1 FILLER_43_135 ();
 FILLCELL_X32 FILLER_43_141 ();
 FILLCELL_X16 FILLER_43_173 ();
 FILLCELL_X8 FILLER_43_189 ();
 FILLCELL_X2 FILLER_43_197 ();
 FILLCELL_X4 FILLER_43_223 ();
 FILLCELL_X2 FILLER_43_227 ();
 FILLCELL_X1 FILLER_43_229 ();
 FILLCELL_X2 FILLER_43_237 ();
 FILLCELL_X1 FILLER_43_239 ();
 FILLCELL_X8 FILLER_43_257 ();
 FILLCELL_X4 FILLER_43_265 ();
 FILLCELL_X1 FILLER_43_269 ();
 FILLCELL_X16 FILLER_43_277 ();
 FILLCELL_X4 FILLER_43_293 ();
 FILLCELL_X1 FILLER_43_297 ();
 FILLCELL_X4 FILLER_43_305 ();
 FILLCELL_X1 FILLER_43_309 ();
 FILLCELL_X1 FILLER_43_315 ();
 FILLCELL_X2 FILLER_43_333 ();
 FILLCELL_X16 FILLER_43_359 ();
 FILLCELL_X4 FILLER_43_375 ();
 FILLCELL_X2 FILLER_43_384 ();
 FILLCELL_X4 FILLER_43_390 ();
 FILLCELL_X4 FILLER_43_401 ();
 FILLCELL_X2 FILLER_43_405 ();
 FILLCELL_X1 FILLER_43_415 ();
 FILLCELL_X16 FILLER_43_433 ();
 FILLCELL_X2 FILLER_43_449 ();
 FILLCELL_X1 FILLER_43_468 ();
 FILLCELL_X16 FILLER_43_486 ();
 FILLCELL_X8 FILLER_43_502 ();
 FILLCELL_X4 FILLER_43_510 ();
 FILLCELL_X2 FILLER_43_514 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X1 FILLER_44_26 ();
 FILLCELL_X2 FILLER_44_48 ();
 FILLCELL_X1 FILLER_44_50 ();
 FILLCELL_X8 FILLER_44_58 ();
 FILLCELL_X2 FILLER_44_66 ();
 FILLCELL_X1 FILLER_44_68 ();
 FILLCELL_X2 FILLER_44_90 ();
 FILLCELL_X1 FILLER_44_92 ();
 FILLCELL_X8 FILLER_44_107 ();
 FILLCELL_X2 FILLER_44_120 ();
 FILLCELL_X2 FILLER_44_139 ();
 FILLCELL_X2 FILLER_44_148 ();
 FILLCELL_X1 FILLER_44_150 ();
 FILLCELL_X2 FILLER_44_168 ();
 FILLCELL_X2 FILLER_44_174 ();
 FILLCELL_X4 FILLER_44_193 ();
 FILLCELL_X4 FILLER_44_235 ();
 FILLCELL_X1 FILLER_44_239 ();
 FILLCELL_X4 FILLER_44_285 ();
 FILLCELL_X2 FILLER_44_289 ();
 FILLCELL_X1 FILLER_44_312 ();
 FILLCELL_X4 FILLER_44_317 ();
 FILLCELL_X4 FILLER_44_337 ();
 FILLCELL_X2 FILLER_44_341 ();
 FILLCELL_X1 FILLER_44_343 ();
 FILLCELL_X8 FILLER_44_359 ();
 FILLCELL_X4 FILLER_44_374 ();
 FILLCELL_X2 FILLER_44_378 ();
 FILLCELL_X1 FILLER_44_380 ();
 FILLCELL_X1 FILLER_44_394 ();
 FILLCELL_X4 FILLER_44_411 ();
 FILLCELL_X4 FILLER_44_422 ();
 FILLCELL_X2 FILLER_44_457 ();
 FILLCELL_X1 FILLER_44_459 ();
 FILLCELL_X8 FILLER_44_481 ();
 FILLCELL_X2 FILLER_44_489 ();
 FILLCELL_X16 FILLER_44_494 ();
 FILLCELL_X4 FILLER_44_510 ();
 FILLCELL_X2 FILLER_44_514 ();
 FILLCELL_X16 FILLER_45_1 ();
 FILLCELL_X8 FILLER_45_17 ();
 FILLCELL_X2 FILLER_45_25 ();
 FILLCELL_X1 FILLER_45_27 ();
 FILLCELL_X4 FILLER_45_35 ();
 FILLCELL_X1 FILLER_45_39 ();
 FILLCELL_X16 FILLER_45_44 ();
 FILLCELL_X8 FILLER_45_60 ();
 FILLCELL_X2 FILLER_45_68 ();
 FILLCELL_X1 FILLER_45_84 ();
 FILLCELL_X8 FILLER_45_90 ();
 FILLCELL_X2 FILLER_45_98 ();
 FILLCELL_X1 FILLER_45_100 ();
 FILLCELL_X4 FILLER_45_191 ();
 FILLCELL_X2 FILLER_45_195 ();
 FILLCELL_X1 FILLER_45_197 ();
 FILLCELL_X8 FILLER_45_222 ();
 FILLCELL_X4 FILLER_45_230 ();
 FILLCELL_X4 FILLER_45_251 ();
 FILLCELL_X2 FILLER_45_255 ();
 FILLCELL_X1 FILLER_45_257 ();
 FILLCELL_X4 FILLER_45_296 ();
 FILLCELL_X4 FILLER_45_307 ();
 FILLCELL_X4 FILLER_45_318 ();
 FILLCELL_X1 FILLER_45_322 ();
 FILLCELL_X16 FILLER_45_330 ();
 FILLCELL_X8 FILLER_45_346 ();
 FILLCELL_X2 FILLER_45_354 ();
 FILLCELL_X1 FILLER_45_363 ();
 FILLCELL_X4 FILLER_45_388 ();
 FILLCELL_X2 FILLER_45_392 ();
 FILLCELL_X8 FILLER_45_407 ();
 FILLCELL_X4 FILLER_45_415 ();
 FILLCELL_X2 FILLER_45_419 ();
 FILLCELL_X1 FILLER_45_421 ();
 FILLCELL_X4 FILLER_45_436 ();
 FILLCELL_X8 FILLER_45_457 ();
 FILLCELL_X1 FILLER_45_465 ();
 FILLCELL_X16 FILLER_45_473 ();
 FILLCELL_X2 FILLER_45_489 ();
 FILLCELL_X1 FILLER_45_491 ();
 FILLCELL_X2 FILLER_45_496 ();
 FILLCELL_X8 FILLER_45_501 ();
 FILLCELL_X4 FILLER_45_509 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X4 FILLER_46_33 ();
 FILLCELL_X2 FILLER_46_37 ();
 FILLCELL_X1 FILLER_46_39 ();
 FILLCELL_X1 FILLER_46_47 ();
 FILLCELL_X8 FILLER_46_89 ();
 FILLCELL_X4 FILLER_46_97 ();
 FILLCELL_X2 FILLER_46_101 ();
 FILLCELL_X1 FILLER_46_103 ();
 FILLCELL_X4 FILLER_46_109 ();
 FILLCELL_X1 FILLER_46_113 ();
 FILLCELL_X2 FILLER_46_117 ();
 FILLCELL_X2 FILLER_46_164 ();
 FILLCELL_X2 FILLER_46_171 ();
 FILLCELL_X32 FILLER_46_187 ();
 FILLCELL_X8 FILLER_46_219 ();
 FILLCELL_X4 FILLER_46_227 ();
 FILLCELL_X8 FILLER_46_245 ();
 FILLCELL_X2 FILLER_46_253 ();
 FILLCELL_X1 FILLER_46_255 ();
 FILLCELL_X8 FILLER_46_280 ();
 FILLCELL_X2 FILLER_46_288 ();
 FILLCELL_X1 FILLER_46_300 ();
 FILLCELL_X4 FILLER_46_306 ();
 FILLCELL_X1 FILLER_46_310 ();
 FILLCELL_X4 FILLER_46_318 ();
 FILLCELL_X2 FILLER_46_322 ();
 FILLCELL_X1 FILLER_46_324 ();
 FILLCELL_X32 FILLER_46_349 ();
 FILLCELL_X4 FILLER_46_381 ();
 FILLCELL_X2 FILLER_46_385 ();
 FILLCELL_X4 FILLER_46_394 ();
 FILLCELL_X1 FILLER_46_398 ();
 FILLCELL_X4 FILLER_46_416 ();
 FILLCELL_X8 FILLER_46_427 ();
 FILLCELL_X4 FILLER_46_435 ();
 FILLCELL_X1 FILLER_46_446 ();
 FILLCELL_X32 FILLER_46_451 ();
 FILLCELL_X4 FILLER_46_483 ();
 FILLCELL_X4 FILLER_46_512 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X8 FILLER_47_33 ();
 FILLCELL_X2 FILLER_47_41 ();
 FILLCELL_X1 FILLER_47_43 ();
 FILLCELL_X2 FILLER_47_51 ();
 FILLCELL_X1 FILLER_47_53 ();
 FILLCELL_X8 FILLER_47_61 ();
 FILLCELL_X1 FILLER_47_69 ();
 FILLCELL_X4 FILLER_47_87 ();
 FILLCELL_X2 FILLER_47_91 ();
 FILLCELL_X1 FILLER_47_103 ();
 FILLCELL_X8 FILLER_47_111 ();
 FILLCELL_X4 FILLER_47_119 ();
 FILLCELL_X32 FILLER_47_128 ();
 FILLCELL_X16 FILLER_47_160 ();
 FILLCELL_X2 FILLER_47_176 ();
 FILLCELL_X1 FILLER_47_178 ();
 FILLCELL_X8 FILLER_47_190 ();
 FILLCELL_X2 FILLER_47_198 ();
 FILLCELL_X16 FILLER_47_224 ();
 FILLCELL_X1 FILLER_47_240 ();
 FILLCELL_X4 FILLER_47_248 ();
 FILLCELL_X4 FILLER_47_261 ();
 FILLCELL_X2 FILLER_47_272 ();
 FILLCELL_X1 FILLER_47_274 ();
 FILLCELL_X4 FILLER_47_299 ();
 FILLCELL_X2 FILLER_47_303 ();
 FILLCELL_X8 FILLER_47_322 ();
 FILLCELL_X1 FILLER_47_330 ();
 FILLCELL_X8 FILLER_47_352 ();
 FILLCELL_X4 FILLER_47_360 ();
 FILLCELL_X1 FILLER_47_409 ();
 FILLCELL_X2 FILLER_47_413 ();
 FILLCELL_X8 FILLER_47_432 ();
 FILLCELL_X4 FILLER_47_440 ();
 FILLCELL_X4 FILLER_47_451 ();
 FILLCELL_X2 FILLER_47_455 ();
 FILLCELL_X1 FILLER_47_471 ();
 FILLCELL_X32 FILLER_47_479 ();
 FILLCELL_X4 FILLER_47_511 ();
 FILLCELL_X1 FILLER_47_515 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X8 FILLER_48_33 ();
 FILLCELL_X2 FILLER_48_41 ();
 FILLCELL_X2 FILLER_48_84 ();
 FILLCELL_X16 FILLER_48_113 ();
 FILLCELL_X8 FILLER_48_129 ();
 FILLCELL_X4 FILLER_48_137 ();
 FILLCELL_X1 FILLER_48_141 ();
 FILLCELL_X1 FILLER_48_166 ();
 FILLCELL_X2 FILLER_48_171 ();
 FILLCELL_X2 FILLER_48_178 ();
 FILLCELL_X2 FILLER_48_197 ();
 FILLCELL_X2 FILLER_48_207 ();
 FILLCELL_X1 FILLER_48_209 ();
 FILLCELL_X4 FILLER_48_217 ();
 FILLCELL_X8 FILLER_48_230 ();
 FILLCELL_X2 FILLER_48_238 ();
 FILLCELL_X16 FILLER_48_257 ();
 FILLCELL_X2 FILLER_48_273 ();
 FILLCELL_X16 FILLER_48_287 ();
 FILLCELL_X4 FILLER_48_303 ();
 FILLCELL_X1 FILLER_48_307 ();
 FILLCELL_X4 FILLER_48_356 ();
 FILLCELL_X2 FILLER_48_360 ();
 FILLCELL_X2 FILLER_48_384 ();
 FILLCELL_X8 FILLER_48_393 ();
 FILLCELL_X2 FILLER_48_401 ();
 FILLCELL_X1 FILLER_48_403 ();
 FILLCELL_X8 FILLER_48_411 ();
 FILLCELL_X4 FILLER_48_467 ();
 FILLCELL_X4 FILLER_48_488 ();
 FILLCELL_X8 FILLER_48_496 ();
 FILLCELL_X4 FILLER_48_504 ();
 FILLCELL_X1 FILLER_48_511 ();
 FILLCELL_X1 FILLER_48_515 ();
 FILLCELL_X8 FILLER_49_1 ();
 FILLCELL_X4 FILLER_49_29 ();
 FILLCELL_X32 FILLER_49_55 ();
 FILLCELL_X4 FILLER_49_87 ();
 FILLCELL_X2 FILLER_49_96 ();
 FILLCELL_X2 FILLER_49_109 ();
 FILLCELL_X1 FILLER_49_111 ();
 FILLCELL_X8 FILLER_49_123 ();
 FILLCELL_X2 FILLER_49_131 ();
 FILLCELL_X4 FILLER_49_140 ();
 FILLCELL_X2 FILLER_49_144 ();
 FILLCELL_X1 FILLER_49_146 ();
 FILLCELL_X8 FILLER_49_159 ();
 FILLCELL_X4 FILLER_49_167 ();
 FILLCELL_X1 FILLER_49_171 ();
 FILLCELL_X2 FILLER_49_188 ();
 FILLCELL_X1 FILLER_49_190 ();
 FILLCELL_X8 FILLER_49_194 ();
 FILLCELL_X4 FILLER_49_202 ();
 FILLCELL_X2 FILLER_49_206 ();
 FILLCELL_X1 FILLER_49_208 ();
 FILLCELL_X8 FILLER_49_226 ();
 FILLCELL_X4 FILLER_49_234 ();
 FILLCELL_X2 FILLER_49_238 ();
 FILLCELL_X2 FILLER_49_247 ();
 FILLCELL_X2 FILLER_49_254 ();
 FILLCELL_X4 FILLER_49_260 ();
 FILLCELL_X2 FILLER_49_264 ();
 FILLCELL_X1 FILLER_49_266 ();
 FILLCELL_X1 FILLER_49_274 ();
 FILLCELL_X16 FILLER_49_282 ();
 FILLCELL_X8 FILLER_49_298 ();
 FILLCELL_X1 FILLER_49_306 ();
 FILLCELL_X8 FILLER_49_317 ();
 FILLCELL_X16 FILLER_49_351 ();
 FILLCELL_X2 FILLER_49_367 ();
 FILLCELL_X16 FILLER_49_383 ();
 FILLCELL_X16 FILLER_49_406 ();
 FILLCELL_X8 FILLER_49_422 ();
 FILLCELL_X4 FILLER_49_430 ();
 FILLCELL_X2 FILLER_49_434 ();
 FILLCELL_X1 FILLER_49_436 ();
 FILLCELL_X1 FILLER_49_445 ();
 FILLCELL_X8 FILLER_49_477 ();
 FILLCELL_X4 FILLER_49_485 ();
 FILLCELL_X2 FILLER_49_489 ();
 FILLCELL_X4 FILLER_49_511 ();
 FILLCELL_X1 FILLER_49_515 ();
 FILLCELL_X8 FILLER_50_1 ();
 FILLCELL_X4 FILLER_50_9 ();
 FILLCELL_X2 FILLER_50_13 ();
 FILLCELL_X8 FILLER_50_56 ();
 FILLCELL_X1 FILLER_50_95 ();
 FILLCELL_X4 FILLER_50_133 ();
 FILLCELL_X4 FILLER_50_154 ();
 FILLCELL_X2 FILLER_50_158 ();
 FILLCELL_X4 FILLER_50_177 ();
 FILLCELL_X8 FILLER_50_201 ();
 FILLCELL_X1 FILLER_50_209 ();
 FILLCELL_X4 FILLER_50_229 ();
 FILLCELL_X2 FILLER_50_233 ();
 FILLCELL_X1 FILLER_50_235 ();
 FILLCELL_X4 FILLER_50_260 ();
 FILLCELL_X1 FILLER_50_264 ();
 FILLCELL_X8 FILLER_50_286 ();
 FILLCELL_X2 FILLER_50_294 ();
 FILLCELL_X1 FILLER_50_296 ();
 FILLCELL_X4 FILLER_50_304 ();
 FILLCELL_X2 FILLER_50_320 ();
 FILLCELL_X1 FILLER_50_327 ();
 FILLCELL_X16 FILLER_50_335 ();
 FILLCELL_X8 FILLER_50_351 ();
 FILLCELL_X4 FILLER_50_359 ();
 FILLCELL_X2 FILLER_50_363 ();
 FILLCELL_X1 FILLER_50_372 ();
 FILLCELL_X2 FILLER_50_378 ();
 FILLCELL_X2 FILLER_50_397 ();
 FILLCELL_X2 FILLER_50_416 ();
 FILLCELL_X4 FILLER_50_425 ();
 FILLCELL_X2 FILLER_50_429 ();
 FILLCELL_X8 FILLER_50_448 ();
 FILLCELL_X32 FILLER_50_463 ();
 FILLCELL_X16 FILLER_50_495 ();
 FILLCELL_X4 FILLER_50_511 ();
 FILLCELL_X1 FILLER_50_515 ();
 FILLCELL_X16 FILLER_51_1 ();
 FILLCELL_X2 FILLER_51_17 ();
 FILLCELL_X1 FILLER_51_19 ();
 FILLCELL_X4 FILLER_51_34 ();
 FILLCELL_X4 FILLER_51_45 ();
 FILLCELL_X2 FILLER_51_49 ();
 FILLCELL_X2 FILLER_51_71 ();
 FILLCELL_X32 FILLER_51_95 ();
 FILLCELL_X2 FILLER_51_127 ();
 FILLCELL_X4 FILLER_51_146 ();
 FILLCELL_X2 FILLER_51_150 ();
 FILLCELL_X1 FILLER_51_176 ();
 FILLCELL_X8 FILLER_51_185 ();
 FILLCELL_X8 FILLER_51_196 ();
 FILLCELL_X2 FILLER_51_204 ();
 FILLCELL_X8 FILLER_51_230 ();
 FILLCELL_X1 FILLER_51_238 ();
 FILLCELL_X8 FILLER_51_260 ();
 FILLCELL_X4 FILLER_51_268 ();
 FILLCELL_X16 FILLER_51_276 ();
 FILLCELL_X8 FILLER_51_338 ();
 FILLCELL_X1 FILLER_51_346 ();
 FILLCELL_X8 FILLER_51_381 ();
 FILLCELL_X4 FILLER_51_389 ();
 FILLCELL_X2 FILLER_51_393 ();
 FILLCELL_X1 FILLER_51_395 ();
 FILLCELL_X1 FILLER_51_421 ();
 FILLCELL_X2 FILLER_51_439 ();
 FILLCELL_X2 FILLER_51_448 ();
 FILLCELL_X32 FILLER_51_474 ();
 FILLCELL_X8 FILLER_51_506 ();
 FILLCELL_X2 FILLER_51_514 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X8 FILLER_52_33 ();
 FILLCELL_X2 FILLER_52_58 ();
 FILLCELL_X1 FILLER_52_60 ();
 FILLCELL_X1 FILLER_52_68 ();
 FILLCELL_X2 FILLER_52_76 ();
 FILLCELL_X2 FILLER_52_85 ();
 FILLCELL_X2 FILLER_52_104 ();
 FILLCELL_X1 FILLER_52_106 ();
 FILLCELL_X32 FILLER_52_124 ();
 FILLCELL_X4 FILLER_52_156 ();
 FILLCELL_X8 FILLER_52_165 ();
 FILLCELL_X2 FILLER_52_173 ();
 FILLCELL_X1 FILLER_52_175 ();
 FILLCELL_X8 FILLER_52_196 ();
 FILLCELL_X2 FILLER_52_204 ();
 FILLCELL_X8 FILLER_52_247 ();
 FILLCELL_X2 FILLER_52_255 ();
 FILLCELL_X32 FILLER_52_280 ();
 FILLCELL_X8 FILLER_52_312 ();
 FILLCELL_X4 FILLER_52_320 ();
 FILLCELL_X1 FILLER_52_324 ();
 FILLCELL_X8 FILLER_52_342 ();
 FILLCELL_X2 FILLER_52_350 ();
 FILLCELL_X2 FILLER_52_359 ();
 FILLCELL_X1 FILLER_52_361 ();
 FILLCELL_X16 FILLER_52_369 ();
 FILLCELL_X4 FILLER_52_385 ();
 FILLCELL_X16 FILLER_52_396 ();
 FILLCELL_X4 FILLER_52_412 ();
 FILLCELL_X2 FILLER_52_449 ();
 FILLCELL_X8 FILLER_52_465 ();
 FILLCELL_X16 FILLER_52_490 ();
 FILLCELL_X8 FILLER_52_506 ();
 FILLCELL_X2 FILLER_52_514 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X8 FILLER_53_33 ();
 FILLCELL_X4 FILLER_53_41 ();
 FILLCELL_X32 FILLER_53_52 ();
 FILLCELL_X1 FILLER_53_84 ();
 FILLCELL_X16 FILLER_53_116 ();
 FILLCELL_X8 FILLER_53_132 ();
 FILLCELL_X1 FILLER_53_140 ();
 FILLCELL_X32 FILLER_53_158 ();
 FILLCELL_X32 FILLER_53_190 ();
 FILLCELL_X8 FILLER_53_222 ();
 FILLCELL_X1 FILLER_53_230 ();
 FILLCELL_X8 FILLER_53_251 ();
 FILLCELL_X4 FILLER_53_259 ();
 FILLCELL_X2 FILLER_53_263 ();
 FILLCELL_X16 FILLER_53_268 ();
 FILLCELL_X8 FILLER_53_284 ();
 FILLCELL_X2 FILLER_53_292 ();
 FILLCELL_X8 FILLER_53_328 ();
 FILLCELL_X2 FILLER_53_336 ();
 FILLCELL_X4 FILLER_53_372 ();
 FILLCELL_X2 FILLER_53_383 ();
 FILLCELL_X1 FILLER_53_385 ();
 FILLCELL_X8 FILLER_53_403 ();
 FILLCELL_X2 FILLER_53_411 ();
 FILLCELL_X8 FILLER_53_444 ();
 FILLCELL_X2 FILLER_53_452 ();
 FILLCELL_X32 FILLER_53_478 ();
 FILLCELL_X4 FILLER_53_510 ();
 FILLCELL_X2 FILLER_53_514 ();
 FILLCELL_X8 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_9 ();
 FILLCELL_X2 FILLER_54_13 ();
 FILLCELL_X1 FILLER_54_15 ();
 FILLCELL_X2 FILLER_54_37 ();
 FILLCELL_X1 FILLER_54_39 ();
 FILLCELL_X8 FILLER_54_74 ();
 FILLCELL_X4 FILLER_54_89 ();
 FILLCELL_X2 FILLER_54_93 ();
 FILLCELL_X1 FILLER_54_95 ();
 FILLCELL_X1 FILLER_54_110 ();
 FILLCELL_X16 FILLER_54_116 ();
 FILLCELL_X2 FILLER_54_132 ();
 FILLCELL_X1 FILLER_54_134 ();
 FILLCELL_X2 FILLER_54_142 ();
 FILLCELL_X1 FILLER_54_144 ();
 FILLCELL_X8 FILLER_54_162 ();
 FILLCELL_X4 FILLER_54_170 ();
 FILLCELL_X2 FILLER_54_174 ();
 FILLCELL_X1 FILLER_54_176 ();
 FILLCELL_X8 FILLER_54_201 ();
 FILLCELL_X1 FILLER_54_209 ();
 FILLCELL_X16 FILLER_54_217 ();
 FILLCELL_X1 FILLER_54_233 ();
 FILLCELL_X16 FILLER_54_241 ();
 FILLCELL_X1 FILLER_54_295 ();
 FILLCELL_X4 FILLER_54_301 ();
 FILLCELL_X2 FILLER_54_312 ();
 FILLCELL_X2 FILLER_54_331 ();
 FILLCELL_X2 FILLER_54_340 ();
 FILLCELL_X2 FILLER_54_349 ();
 FILLCELL_X1 FILLER_54_351 ();
 FILLCELL_X2 FILLER_54_366 ();
 FILLCELL_X1 FILLER_54_368 ();
 FILLCELL_X2 FILLER_54_386 ();
 FILLCELL_X4 FILLER_54_446 ();
 FILLCELL_X4 FILLER_54_458 ();
 FILLCELL_X1 FILLER_54_462 ();
 FILLCELL_X32 FILLER_54_470 ();
 FILLCELL_X8 FILLER_54_502 ();
 FILLCELL_X4 FILLER_54_510 ();
 FILLCELL_X2 FILLER_54_514 ();
 FILLCELL_X8 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_9 ();
 FILLCELL_X1 FILLER_55_13 ();
 FILLCELL_X1 FILLER_55_31 ();
 FILLCELL_X2 FILLER_55_68 ();
 FILLCELL_X2 FILLER_55_77 ();
 FILLCELL_X16 FILLER_55_96 ();
 FILLCELL_X4 FILLER_55_112 ();
 FILLCELL_X2 FILLER_55_116 ();
 FILLCELL_X1 FILLER_55_118 ();
 FILLCELL_X4 FILLER_55_136 ();
 FILLCELL_X2 FILLER_55_140 ();
 FILLCELL_X2 FILLER_55_180 ();
 FILLCELL_X2 FILLER_55_223 ();
 FILLCELL_X4 FILLER_55_228 ();
 FILLCELL_X2 FILLER_55_232 ();
 FILLCELL_X1 FILLER_55_234 ();
 FILLCELL_X8 FILLER_55_252 ();
 FILLCELL_X2 FILLER_55_308 ();
 FILLCELL_X4 FILLER_55_324 ();
 FILLCELL_X2 FILLER_55_328 ();
 FILLCELL_X1 FILLER_55_330 ();
 FILLCELL_X16 FILLER_55_360 ();
 FILLCELL_X4 FILLER_55_376 ();
 FILLCELL_X16 FILLER_55_401 ();
 FILLCELL_X4 FILLER_55_417 ();
 FILLCELL_X8 FILLER_55_435 ();
 FILLCELL_X2 FILLER_55_443 ();
 FILLCELL_X8 FILLER_55_455 ();
 FILLCELL_X1 FILLER_55_463 ();
 FILLCELL_X16 FILLER_55_481 ();
 FILLCELL_X8 FILLER_55_497 ();
 FILLCELL_X2 FILLER_55_505 ();
 FILLCELL_X1 FILLER_55_507 ();
 FILLCELL_X4 FILLER_55_511 ();
 FILLCELL_X1 FILLER_55_515 ();
 FILLCELL_X16 FILLER_56_1 ();
 FILLCELL_X4 FILLER_56_17 ();
 FILLCELL_X1 FILLER_56_21 ();
 FILLCELL_X1 FILLER_56_36 ();
 FILLCELL_X4 FILLER_56_44 ();
 FILLCELL_X1 FILLER_56_48 ();
 FILLCELL_X4 FILLER_56_62 ();
 FILLCELL_X1 FILLER_56_66 ();
 FILLCELL_X4 FILLER_56_74 ();
 FILLCELL_X16 FILLER_56_92 ();
 FILLCELL_X2 FILLER_56_108 ();
 FILLCELL_X1 FILLER_56_110 ();
 FILLCELL_X2 FILLER_56_186 ();
 FILLCELL_X4 FILLER_56_202 ();
 FILLCELL_X2 FILLER_56_232 ();
 FILLCELL_X8 FILLER_56_248 ();
 FILLCELL_X4 FILLER_56_256 ();
 FILLCELL_X1 FILLER_56_260 ();
 FILLCELL_X16 FILLER_56_278 ();
 FILLCELL_X2 FILLER_56_294 ();
 FILLCELL_X2 FILLER_56_299 ();
 FILLCELL_X1 FILLER_56_313 ();
 FILLCELL_X2 FILLER_56_331 ();
 FILLCELL_X2 FILLER_56_347 ();
 FILLCELL_X2 FILLER_56_366 ();
 FILLCELL_X1 FILLER_56_368 ();
 FILLCELL_X2 FILLER_56_374 ();
 FILLCELL_X1 FILLER_56_376 ();
 FILLCELL_X32 FILLER_56_384 ();
 FILLCELL_X1 FILLER_56_416 ();
 FILLCELL_X2 FILLER_56_422 ();
 FILLCELL_X8 FILLER_56_431 ();
 FILLCELL_X1 FILLER_56_439 ();
 FILLCELL_X16 FILLER_56_471 ();
 FILLCELL_X1 FILLER_56_487 ();
 FILLCELL_X8 FILLER_56_508 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X16 FILLER_57_65 ();
 FILLCELL_X8 FILLER_57_81 ();
 FILLCELL_X1 FILLER_57_89 ();
 FILLCELL_X2 FILLER_57_102 ();
 FILLCELL_X8 FILLER_57_111 ();
 FILLCELL_X8 FILLER_57_143 ();
 FILLCELL_X2 FILLER_57_151 ();
 FILLCELL_X8 FILLER_57_172 ();
 FILLCELL_X2 FILLER_57_187 ();
 FILLCELL_X1 FILLER_57_189 ();
 FILLCELL_X1 FILLER_57_197 ();
 FILLCELL_X2 FILLER_57_203 ();
 FILLCELL_X1 FILLER_57_212 ();
 FILLCELL_X1 FILLER_57_230 ();
 FILLCELL_X4 FILLER_57_238 ();
 FILLCELL_X4 FILLER_57_259 ();
 FILLCELL_X1 FILLER_57_263 ();
 FILLCELL_X4 FILLER_57_269 ();
 FILLCELL_X2 FILLER_57_273 ();
 FILLCELL_X8 FILLER_57_282 ();
 FILLCELL_X2 FILLER_57_290 ();
 FILLCELL_X1 FILLER_57_292 ();
 FILLCELL_X2 FILLER_57_300 ();
 FILLCELL_X16 FILLER_57_305 ();
 FILLCELL_X8 FILLER_57_321 ();
 FILLCELL_X4 FILLER_57_329 ();
 FILLCELL_X8 FILLER_57_340 ();
 FILLCELL_X4 FILLER_57_348 ();
 FILLCELL_X1 FILLER_57_352 ();
 FILLCELL_X8 FILLER_57_383 ();
 FILLCELL_X1 FILLER_57_391 ();
 FILLCELL_X8 FILLER_57_399 ();
 FILLCELL_X2 FILLER_57_407 ();
 FILLCELL_X8 FILLER_57_416 ();
 FILLCELL_X2 FILLER_57_424 ();
 FILLCELL_X1 FILLER_57_426 ();
 FILLCELL_X4 FILLER_57_430 ();
 FILLCELL_X8 FILLER_57_441 ();
 FILLCELL_X1 FILLER_57_449 ();
 FILLCELL_X4 FILLER_57_457 ();
 FILLCELL_X2 FILLER_57_461 ();
 FILLCELL_X2 FILLER_57_491 ();
 FILLCELL_X1 FILLER_57_493 ();
 FILLCELL_X16 FILLER_57_497 ();
 FILLCELL_X2 FILLER_57_513 ();
 FILLCELL_X1 FILLER_57_515 ();
 FILLCELL_X16 FILLER_58_1 ();
 FILLCELL_X8 FILLER_58_17 ();
 FILLCELL_X2 FILLER_58_25 ();
 FILLCELL_X1 FILLER_58_27 ();
 FILLCELL_X32 FILLER_58_32 ();
 FILLCELL_X2 FILLER_58_64 ();
 FILLCELL_X8 FILLER_58_83 ();
 FILLCELL_X2 FILLER_58_91 ();
 FILLCELL_X16 FILLER_58_110 ();
 FILLCELL_X16 FILLER_58_133 ();
 FILLCELL_X1 FILLER_58_149 ();
 FILLCELL_X16 FILLER_58_170 ();
 FILLCELL_X4 FILLER_58_186 ();
 FILLCELL_X1 FILLER_58_190 ();
 FILLCELL_X8 FILLER_58_194 ();
 FILLCELL_X2 FILLER_58_202 ();
 FILLCELL_X4 FILLER_58_221 ();
 FILLCELL_X2 FILLER_58_225 ();
 FILLCELL_X1 FILLER_58_227 ();
 FILLCELL_X2 FILLER_58_252 ();
 FILLCELL_X2 FILLER_58_271 ();
 FILLCELL_X1 FILLER_58_273 ();
 FILLCELL_X8 FILLER_58_277 ();
 FILLCELL_X2 FILLER_58_285 ();
 FILLCELL_X8 FILLER_58_304 ();
 FILLCELL_X32 FILLER_58_319 ();
 FILLCELL_X8 FILLER_58_351 ();
 FILLCELL_X1 FILLER_58_359 ();
 FILLCELL_X16 FILLER_58_365 ();
 FILLCELL_X1 FILLER_58_388 ();
 FILLCELL_X8 FILLER_58_423 ();
 FILLCELL_X1 FILLER_58_431 ();
 FILLCELL_X32 FILLER_58_466 ();
 FILLCELL_X16 FILLER_58_498 ();
 FILLCELL_X2 FILLER_58_514 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X8 FILLER_59_17 ();
 FILLCELL_X4 FILLER_59_66 ();
 FILLCELL_X1 FILLER_59_70 ();
 FILLCELL_X2 FILLER_59_85 ();
 FILLCELL_X1 FILLER_59_87 ();
 FILLCELL_X4 FILLER_59_93 ();
 FILLCELL_X1 FILLER_59_97 ();
 FILLCELL_X16 FILLER_59_118 ();
 FILLCELL_X1 FILLER_59_134 ();
 FILLCELL_X2 FILLER_59_142 ();
 FILLCELL_X16 FILLER_59_158 ();
 FILLCELL_X16 FILLER_59_205 ();
 FILLCELL_X8 FILLER_59_221 ();
 FILLCELL_X4 FILLER_59_229 ();
 FILLCELL_X2 FILLER_59_233 ();
 FILLCELL_X1 FILLER_59_235 ();
 FILLCELL_X4 FILLER_59_253 ();
 FILLCELL_X1 FILLER_59_257 ();
 FILLCELL_X16 FILLER_59_265 ();
 FILLCELL_X4 FILLER_59_281 ();
 FILLCELL_X2 FILLER_59_285 ();
 FILLCELL_X1 FILLER_59_287 ();
 FILLCELL_X8 FILLER_59_327 ();
 FILLCELL_X2 FILLER_59_335 ();
 FILLCELL_X8 FILLER_59_361 ();
 FILLCELL_X4 FILLER_59_369 ();
 FILLCELL_X2 FILLER_59_373 ();
 FILLCELL_X1 FILLER_59_375 ();
 FILLCELL_X2 FILLER_59_393 ();
 FILLCELL_X1 FILLER_59_395 ();
 FILLCELL_X4 FILLER_59_401 ();
 FILLCELL_X2 FILLER_59_405 ();
 FILLCELL_X32 FILLER_59_431 ();
 FILLCELL_X32 FILLER_59_463 ();
 FILLCELL_X16 FILLER_59_495 ();
 FILLCELL_X4 FILLER_59_511 ();
 FILLCELL_X1 FILLER_59_515 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X2 FILLER_60_54 ();
 FILLCELL_X2 FILLER_60_73 ();
 FILLCELL_X1 FILLER_60_75 ();
 FILLCELL_X2 FILLER_60_93 ();
 FILLCELL_X1 FILLER_60_95 ();
 FILLCELL_X4 FILLER_60_99 ();
 FILLCELL_X2 FILLER_60_103 ();
 FILLCELL_X1 FILLER_60_105 ();
 FILLCELL_X1 FILLER_60_123 ();
 FILLCELL_X16 FILLER_60_163 ();
 FILLCELL_X8 FILLER_60_179 ();
 FILLCELL_X1 FILLER_60_187 ();
 FILLCELL_X16 FILLER_60_217 ();
 FILLCELL_X2 FILLER_60_233 ();
 FILLCELL_X1 FILLER_60_242 ();
 FILLCELL_X2 FILLER_60_250 ();
 FILLCELL_X1 FILLER_60_252 ();
 FILLCELL_X16 FILLER_60_258 ();
 FILLCELL_X1 FILLER_60_274 ();
 FILLCELL_X8 FILLER_60_283 ();
 FILLCELL_X1 FILLER_60_291 ();
 FILLCELL_X32 FILLER_60_308 ();
 FILLCELL_X2 FILLER_60_340 ();
 FILLCELL_X4 FILLER_60_349 ();
 FILLCELL_X1 FILLER_60_353 ();
 FILLCELL_X4 FILLER_60_376 ();
 FILLCELL_X1 FILLER_60_380 ();
 FILLCELL_X2 FILLER_60_388 ();
 FILLCELL_X4 FILLER_60_411 ();
 FILLCELL_X32 FILLER_60_422 ();
 FILLCELL_X4 FILLER_60_454 ();
 FILLCELL_X2 FILLER_60_458 ();
 FILLCELL_X32 FILLER_60_465 ();
 FILLCELL_X16 FILLER_60_497 ();
 FILLCELL_X2 FILLER_60_513 ();
 FILLCELL_X1 FILLER_60_515 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X16 FILLER_61_33 ();
 FILLCELL_X4 FILLER_61_49 ();
 FILLCELL_X2 FILLER_61_53 ();
 FILLCELL_X1 FILLER_61_86 ();
 FILLCELL_X2 FILLER_61_92 ();
 FILLCELL_X1 FILLER_61_94 ();
 FILLCELL_X2 FILLER_61_99 ();
 FILLCELL_X1 FILLER_61_101 ();
 FILLCELL_X32 FILLER_61_113 ();
 FILLCELL_X8 FILLER_61_145 ();
 FILLCELL_X4 FILLER_61_153 ();
 FILLCELL_X2 FILLER_61_157 ();
 FILLCELL_X1 FILLER_61_159 ();
 FILLCELL_X16 FILLER_61_164 ();
 FILLCELL_X8 FILLER_61_187 ();
 FILLCELL_X4 FILLER_61_195 ();
 FILLCELL_X2 FILLER_61_199 ();
 FILLCELL_X1 FILLER_61_201 ();
 FILLCELL_X16 FILLER_61_223 ();
 FILLCELL_X1 FILLER_61_239 ();
 FILLCELL_X2 FILLER_61_268 ();
 FILLCELL_X16 FILLER_61_274 ();
 FILLCELL_X8 FILLER_61_290 ();
 FILLCELL_X1 FILLER_61_302 ();
 FILLCELL_X2 FILLER_61_308 ();
 FILLCELL_X1 FILLER_61_310 ();
 FILLCELL_X8 FILLER_61_314 ();
 FILLCELL_X16 FILLER_61_329 ();
 FILLCELL_X8 FILLER_61_345 ();
 FILLCELL_X4 FILLER_61_353 ();
 FILLCELL_X1 FILLER_61_357 ();
 FILLCELL_X2 FILLER_61_362 ();
 FILLCELL_X1 FILLER_61_364 ();
 FILLCELL_X4 FILLER_61_372 ();
 FILLCELL_X1 FILLER_61_376 ();
 FILLCELL_X4 FILLER_61_426 ();
 FILLCELL_X2 FILLER_61_430 ();
 FILLCELL_X32 FILLER_61_480 ();
 FILLCELL_X4 FILLER_61_512 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X8 FILLER_62_33 ();
 FILLCELL_X2 FILLER_62_41 ();
 FILLCELL_X1 FILLER_62_43 ();
 FILLCELL_X1 FILLER_62_78 ();
 FILLCELL_X4 FILLER_62_86 ();
 FILLCELL_X2 FILLER_62_90 ();
 FILLCELL_X1 FILLER_62_92 ();
 FILLCELL_X2 FILLER_62_118 ();
 FILLCELL_X1 FILLER_62_120 ();
 FILLCELL_X4 FILLER_62_145 ();
 FILLCELL_X2 FILLER_62_149 ();
 FILLCELL_X1 FILLER_62_151 ();
 FILLCELL_X1 FILLER_62_159 ();
 FILLCELL_X4 FILLER_62_169 ();
 FILLCELL_X2 FILLER_62_173 ();
 FILLCELL_X1 FILLER_62_175 ();
 FILLCELL_X1 FILLER_62_193 ();
 FILLCELL_X4 FILLER_62_198 ();
 FILLCELL_X8 FILLER_62_217 ();
 FILLCELL_X4 FILLER_62_225 ();
 FILLCELL_X2 FILLER_62_229 ();
 FILLCELL_X1 FILLER_62_231 ();
 FILLCELL_X8 FILLER_62_271 ();
 FILLCELL_X4 FILLER_62_279 ();
 FILLCELL_X1 FILLER_62_314 ();
 FILLCELL_X4 FILLER_62_332 ();
 FILLCELL_X2 FILLER_62_353 ();
 FILLCELL_X1 FILLER_62_355 ();
 FILLCELL_X1 FILLER_62_365 ();
 FILLCELL_X4 FILLER_62_383 ();
 FILLCELL_X2 FILLER_62_398 ();
 FILLCELL_X4 FILLER_62_405 ();
 FILLCELL_X1 FILLER_62_409 ();
 FILLCELL_X1 FILLER_62_413 ();
 FILLCELL_X8 FILLER_62_442 ();
 FILLCELL_X4 FILLER_62_450 ();
 FILLCELL_X32 FILLER_62_464 ();
 FILLCELL_X16 FILLER_62_496 ();
 FILLCELL_X4 FILLER_62_512 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X8 FILLER_63_33 ();
 FILLCELL_X1 FILLER_63_41 ();
 FILLCELL_X8 FILLER_63_49 ();
 FILLCELL_X2 FILLER_63_57 ();
 FILLCELL_X2 FILLER_63_73 ();
 FILLCELL_X4 FILLER_63_99 ();
 FILLCELL_X2 FILLER_63_103 ();
 FILLCELL_X8 FILLER_63_112 ();
 FILLCELL_X4 FILLER_63_120 ();
 FILLCELL_X1 FILLER_63_124 ();
 FILLCELL_X1 FILLER_63_149 ();
 FILLCELL_X8 FILLER_63_167 ();
 FILLCELL_X4 FILLER_63_175 ();
 FILLCELL_X2 FILLER_63_179 ();
 FILLCELL_X2 FILLER_63_205 ();
 FILLCELL_X8 FILLER_63_214 ();
 FILLCELL_X2 FILLER_63_222 ();
 FILLCELL_X2 FILLER_63_238 ();
 FILLCELL_X2 FILLER_63_247 ();
 FILLCELL_X1 FILLER_63_249 ();
 FILLCELL_X2 FILLER_63_257 ();
 FILLCELL_X1 FILLER_63_259 ();
 FILLCELL_X2 FILLER_63_263 ();
 FILLCELL_X8 FILLER_63_272 ();
 FILLCELL_X4 FILLER_63_280 ();
 FILLCELL_X2 FILLER_63_284 ();
 FILLCELL_X2 FILLER_63_310 ();
 FILLCELL_X8 FILLER_63_319 ();
 FILLCELL_X4 FILLER_63_327 ();
 FILLCELL_X2 FILLER_63_331 ();
 FILLCELL_X16 FILLER_63_360 ();
 FILLCELL_X2 FILLER_63_376 ();
 FILLCELL_X2 FILLER_63_399 ();
 FILLCELL_X1 FILLER_63_404 ();
 FILLCELL_X16 FILLER_63_424 ();
 FILLCELL_X1 FILLER_63_440 ();
 FILLCELL_X8 FILLER_63_448 ();
 FILLCELL_X1 FILLER_63_456 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X2 FILLER_63_513 ();
 FILLCELL_X1 FILLER_63_515 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X1 FILLER_64_65 ();
 FILLCELL_X16 FILLER_64_70 ();
 FILLCELL_X4 FILLER_64_86 ();
 FILLCELL_X1 FILLER_64_90 ();
 FILLCELL_X2 FILLER_64_108 ();
 FILLCELL_X1 FILLER_64_110 ();
 FILLCELL_X16 FILLER_64_114 ();
 FILLCELL_X8 FILLER_64_130 ();
 FILLCELL_X1 FILLER_64_138 ();
 FILLCELL_X2 FILLER_64_146 ();
 FILLCELL_X16 FILLER_64_173 ();
 FILLCELL_X4 FILLER_64_189 ();
 FILLCELL_X1 FILLER_64_193 ();
 FILLCELL_X1 FILLER_64_198 ();
 FILLCELL_X16 FILLER_64_216 ();
 FILLCELL_X8 FILLER_64_232 ();
 FILLCELL_X2 FILLER_64_240 ();
 FILLCELL_X4 FILLER_64_259 ();
 FILLCELL_X1 FILLER_64_263 ();
 FILLCELL_X16 FILLER_64_281 ();
 FILLCELL_X4 FILLER_64_297 ();
 FILLCELL_X2 FILLER_64_301 ();
 FILLCELL_X8 FILLER_64_331 ();
 FILLCELL_X1 FILLER_64_339 ();
 FILLCELL_X8 FILLER_64_354 ();
 FILLCELL_X2 FILLER_64_362 ();
 FILLCELL_X1 FILLER_64_364 ();
 FILLCELL_X8 FILLER_64_379 ();
 FILLCELL_X4 FILLER_64_387 ();
 FILLCELL_X2 FILLER_64_391 ();
 FILLCELL_X4 FILLER_64_407 ();
 FILLCELL_X4 FILLER_64_414 ();
 FILLCELL_X4 FILLER_64_435 ();
 FILLCELL_X2 FILLER_64_439 ();
 FILLCELL_X32 FILLER_64_448 ();
 FILLCELL_X32 FILLER_64_480 ();
 FILLCELL_X4 FILLER_64_512 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X16 FILLER_65_65 ();
 FILLCELL_X4 FILLER_65_81 ();
 FILLCELL_X8 FILLER_65_92 ();
 FILLCELL_X4 FILLER_65_100 ();
 FILLCELL_X2 FILLER_65_104 ();
 FILLCELL_X16 FILLER_65_113 ();
 FILLCELL_X8 FILLER_65_129 ();
 FILLCELL_X4 FILLER_65_137 ();
 FILLCELL_X2 FILLER_65_141 ();
 FILLCELL_X4 FILLER_65_164 ();
 FILLCELL_X1 FILLER_65_168 ();
 FILLCELL_X8 FILLER_65_176 ();
 FILLCELL_X4 FILLER_65_184 ();
 FILLCELL_X1 FILLER_65_188 ();
 FILLCELL_X32 FILLER_65_218 ();
 FILLCELL_X2 FILLER_65_250 ();
 FILLCELL_X1 FILLER_65_252 ();
 FILLCELL_X8 FILLER_65_257 ();
 FILLCELL_X2 FILLER_65_265 ();
 FILLCELL_X16 FILLER_65_274 ();
 FILLCELL_X4 FILLER_65_290 ();
 FILLCELL_X8 FILLER_65_299 ();
 FILLCELL_X2 FILLER_65_307 ();
 FILLCELL_X4 FILLER_65_312 ();
 FILLCELL_X16 FILLER_65_323 ();
 FILLCELL_X8 FILLER_65_339 ();
 FILLCELL_X4 FILLER_65_347 ();
 FILLCELL_X2 FILLER_65_351 ();
 FILLCELL_X2 FILLER_65_360 ();
 FILLCELL_X4 FILLER_65_383 ();
 FILLCELL_X2 FILLER_65_387 ();
 FILLCELL_X4 FILLER_65_406 ();
 FILLCELL_X2 FILLER_65_410 ();
 FILLCELL_X16 FILLER_65_417 ();
 FILLCELL_X4 FILLER_65_433 ();
 FILLCELL_X2 FILLER_65_437 ();
 FILLCELL_X1 FILLER_65_439 ();
 FILLCELL_X32 FILLER_65_461 ();
 FILLCELL_X16 FILLER_65_493 ();
 FILLCELL_X4 FILLER_65_509 ();
 FILLCELL_X2 FILLER_65_513 ();
 FILLCELL_X1 FILLER_65_515 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X16 FILLER_66_65 ();
 FILLCELL_X4 FILLER_66_105 ();
 FILLCELL_X1 FILLER_66_125 ();
 FILLCELL_X8 FILLER_66_129 ();
 FILLCELL_X4 FILLER_66_137 ();
 FILLCELL_X1 FILLER_66_141 ();
 FILLCELL_X8 FILLER_66_174 ();
 FILLCELL_X4 FILLER_66_209 ();
 FILLCELL_X2 FILLER_66_230 ();
 FILLCELL_X2 FILLER_66_246 ();
 FILLCELL_X2 FILLER_66_255 ();
 FILLCELL_X16 FILLER_66_265 ();
 FILLCELL_X1 FILLER_66_281 ();
 FILLCELL_X1 FILLER_66_311 ();
 FILLCELL_X8 FILLER_66_329 ();
 FILLCELL_X4 FILLER_66_337 ();
 FILLCELL_X1 FILLER_66_341 ();
 FILLCELL_X2 FILLER_66_368 ();
 FILLCELL_X16 FILLER_66_373 ();
 FILLCELL_X8 FILLER_66_396 ();
 FILLCELL_X4 FILLER_66_404 ();
 FILLCELL_X1 FILLER_66_408 ();
 FILLCELL_X4 FILLER_66_428 ();
 FILLCELL_X2 FILLER_66_432 ();
 FILLCELL_X1 FILLER_66_434 ();
 FILLCELL_X32 FILLER_66_442 ();
 FILLCELL_X32 FILLER_66_474 ();
 FILLCELL_X8 FILLER_66_506 ();
 FILLCELL_X2 FILLER_66_514 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X16 FILLER_67_65 ();
 FILLCELL_X4 FILLER_67_81 ();
 FILLCELL_X2 FILLER_67_85 ();
 FILLCELL_X1 FILLER_67_87 ();
 FILLCELL_X2 FILLER_67_132 ();
 FILLCELL_X1 FILLER_67_151 ();
 FILLCELL_X8 FILLER_67_159 ();
 FILLCELL_X4 FILLER_67_167 ();
 FILLCELL_X2 FILLER_67_171 ();
 FILLCELL_X1 FILLER_67_173 ();
 FILLCELL_X2 FILLER_67_178 ();
 FILLCELL_X2 FILLER_67_197 ();
 FILLCELL_X2 FILLER_67_206 ();
 FILLCELL_X4 FILLER_67_213 ();
 FILLCELL_X1 FILLER_67_221 ();
 FILLCELL_X4 FILLER_67_225 ();
 FILLCELL_X2 FILLER_67_229 ();
 FILLCELL_X2 FILLER_67_248 ();
 FILLCELL_X2 FILLER_67_267 ();
 FILLCELL_X1 FILLER_67_269 ();
 FILLCELL_X4 FILLER_67_277 ();
 FILLCELL_X2 FILLER_67_281 ();
 FILLCELL_X1 FILLER_67_315 ();
 FILLCELL_X4 FILLER_67_336 ();
 FILLCELL_X2 FILLER_67_340 ();
 FILLCELL_X4 FILLER_67_380 ();
 FILLCELL_X2 FILLER_67_384 ();
 FILLCELL_X1 FILLER_67_410 ();
 FILLCELL_X4 FILLER_67_415 ();
 FILLCELL_X2 FILLER_67_419 ();
 FILLCELL_X1 FILLER_67_421 ();
 FILLCELL_X32 FILLER_67_456 ();
 FILLCELL_X16 FILLER_67_488 ();
 FILLCELL_X8 FILLER_67_504 ();
 FILLCELL_X4 FILLER_67_512 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X16 FILLER_68_65 ();
 FILLCELL_X4 FILLER_68_81 ();
 FILLCELL_X1 FILLER_68_85 ();
 FILLCELL_X2 FILLER_68_110 ();
 FILLCELL_X1 FILLER_68_112 ();
 FILLCELL_X4 FILLER_68_133 ();
 FILLCELL_X1 FILLER_68_137 ();
 FILLCELL_X4 FILLER_68_145 ();
 FILLCELL_X2 FILLER_68_193 ();
 FILLCELL_X1 FILLER_68_235 ();
 FILLCELL_X2 FILLER_68_253 ();
 FILLCELL_X1 FILLER_68_255 ();
 FILLCELL_X4 FILLER_68_263 ();
 FILLCELL_X1 FILLER_68_267 ();
 FILLCELL_X4 FILLER_68_288 ();
 FILLCELL_X1 FILLER_68_292 ();
 FILLCELL_X4 FILLER_68_300 ();
 FILLCELL_X4 FILLER_68_330 ();
 FILLCELL_X2 FILLER_68_334 ();
 FILLCELL_X1 FILLER_68_360 ();
 FILLCELL_X8 FILLER_68_381 ();
 FILLCELL_X2 FILLER_68_389 ();
 FILLCELL_X1 FILLER_68_391 ();
 FILLCELL_X1 FILLER_68_409 ();
 FILLCELL_X4 FILLER_68_434 ();
 FILLCELL_X2 FILLER_68_438 ();
 FILLCELL_X1 FILLER_68_440 ();
 FILLCELL_X32 FILLER_68_445 ();
 FILLCELL_X32 FILLER_68_477 ();
 FILLCELL_X4 FILLER_68_509 ();
 FILLCELL_X2 FILLER_68_513 ();
 FILLCELL_X1 FILLER_68_515 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X16 FILLER_69_33 ();
 FILLCELL_X4 FILLER_69_49 ();
 FILLCELL_X1 FILLER_69_53 ();
 FILLCELL_X32 FILLER_69_58 ();
 FILLCELL_X32 FILLER_69_90 ();
 FILLCELL_X2 FILLER_69_122 ();
 FILLCELL_X4 FILLER_69_130 ();
 FILLCELL_X1 FILLER_69_134 ();
 FILLCELL_X32 FILLER_69_138 ();
 FILLCELL_X4 FILLER_69_170 ();
 FILLCELL_X2 FILLER_69_174 ();
 FILLCELL_X4 FILLER_69_179 ();
 FILLCELL_X4 FILLER_69_186 ();
 FILLCELL_X1 FILLER_69_190 ();
 FILLCELL_X2 FILLER_69_194 ();
 FILLCELL_X32 FILLER_69_199 ();
 FILLCELL_X4 FILLER_69_231 ();
 FILLCELL_X8 FILLER_69_238 ();
 FILLCELL_X2 FILLER_69_246 ();
 FILLCELL_X2 FILLER_69_251 ();
 FILLCELL_X1 FILLER_69_253 ();
 FILLCELL_X16 FILLER_69_257 ();
 FILLCELL_X8 FILLER_69_273 ();
 FILLCELL_X1 FILLER_69_281 ();
 FILLCELL_X4 FILLER_69_285 ();
 FILLCELL_X4 FILLER_69_292 ();
 FILLCELL_X1 FILLER_69_296 ();
 FILLCELL_X16 FILLER_69_300 ();
 FILLCELL_X2 FILLER_69_316 ();
 FILLCELL_X32 FILLER_69_324 ();
 FILLCELL_X16 FILLER_69_356 ();
 FILLCELL_X2 FILLER_69_372 ();
 FILLCELL_X1 FILLER_69_374 ();
 FILLCELL_X4 FILLER_69_381 ();
 FILLCELL_X16 FILLER_69_389 ();
 FILLCELL_X4 FILLER_69_405 ();
 FILLCELL_X1 FILLER_69_412 ();
 FILLCELL_X32 FILLER_69_416 ();
 FILLCELL_X32 FILLER_69_448 ();
 FILLCELL_X32 FILLER_69_480 ();
 FILLCELL_X4 FILLER_69_512 ();
endmodule
