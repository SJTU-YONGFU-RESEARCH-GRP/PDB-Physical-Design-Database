module hamming_code (single_bit_error,
    corrected_code,
    data_in,
    data_out,
    encoded_out,
    received_in);
 output single_bit_error;
 output [6:0] corrected_code;
 input [3:0] data_in;
 output [3:0] data_out;
 output [6:0] encoded_out;
 input [6:0] received_in;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire p1;
 wire p2;
 wire p3;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;

 BUF_X2 _081_ (.A(received_in[5]),
    .Z(_010_));
 CLKBUF_X3 _082_ (.A(received_in[3]),
    .Z(_011_));
 XNOR2_X1 _083_ (.A(_010_),
    .B(_011_),
    .ZN(_012_));
 XNOR2_X1 _084_ (.A(net6),
    .B(net7),
    .ZN(_013_));
 NOR2_X1 _085_ (.A1(_012_),
    .A2(_013_),
    .ZN(_014_));
 AND2_X1 _086_ (.A1(_012_),
    .A2(_013_),
    .ZN(_015_));
 BUF_X4 _087_ (.A(received_in[2]),
    .Z(_016_));
 XOR2_X2 _088_ (.A(_016_),
    .B(net5),
    .Z(_017_));
 BUF_X4 _089_ (.A(_017_),
    .Z(_018_));
 MUX2_X1 _090_ (.A(_014_),
    .B(_015_),
    .S(_018_),
    .Z(_019_));
 CLKBUF_X2 _091_ (.A(received_in[1]),
    .Z(_020_));
 XNOR2_X2 _092_ (.A(_016_),
    .B(_020_),
    .ZN(_021_));
 BUF_X4 _093_ (.A(_021_),
    .Z(_022_));
 BUF_X4 _094_ (.A(net7),
    .Z(_023_));
 XNOR2_X2 _095_ (.A(_023_),
    .B(_010_),
    .ZN(_024_));
 XNOR2_X1 _096_ (.A(_022_),
    .B(_024_),
    .ZN(_025_));
 NAND2_X1 _097_ (.A1(_019_),
    .A2(_025_),
    .ZN(_026_));
 XNOR2_X1 _098_ (.A(net5),
    .B(_026_),
    .ZN(net8));
 XNOR2_X1 _099_ (.A(_016_),
    .B(_024_),
    .ZN(_027_));
 XNOR2_X2 _100_ (.A(_016_),
    .B(net5),
    .ZN(_028_));
 MUX2_X1 _101_ (.A(_014_),
    .B(_015_),
    .S(_028_),
    .Z(_029_));
 MUX2_X1 _102_ (.A(_020_),
    .B(_027_),
    .S(_029_),
    .Z(net9));
 XNOR2_X1 _103_ (.A(_020_),
    .B(_024_),
    .ZN(_030_));
 MUX2_X1 _104_ (.A(_016_),
    .B(_030_),
    .S(_019_),
    .Z(net10));
 NOR2_X1 _105_ (.A1(_011_),
    .A2(_028_),
    .ZN(_031_));
 CLKBUF_X3 _106_ (.A(_011_),
    .Z(_032_));
 XOR2_X2 _107_ (.A(_016_),
    .B(_020_),
    .Z(_033_));
 OAI21_X1 _108_ (.A(_032_),
    .B1(_018_),
    .B2(_033_),
    .ZN(_034_));
 INV_X2 _109_ (.A(_010_),
    .ZN(_035_));
 AOI21_X1 _110_ (.A(_031_),
    .B1(_034_),
    .B2(_035_),
    .ZN(_036_));
 NOR2_X1 _111_ (.A1(_023_),
    .A2(_036_),
    .ZN(_037_));
 INV_X1 _112_ (.A(_023_),
    .ZN(_038_));
 INV_X2 _113_ (.A(_011_),
    .ZN(_039_));
 AOI21_X1 _114_ (.A(_039_),
    .B1(_018_),
    .B2(_022_),
    .ZN(_040_));
 CLKBUF_X3 _115_ (.A(_010_),
    .Z(_041_));
 NOR2_X1 _116_ (.A1(_041_),
    .A2(_028_),
    .ZN(_042_));
 NOR3_X1 _117_ (.A1(_038_),
    .A2(_040_),
    .A3(_042_),
    .ZN(_043_));
 CLKBUF_X3 _118_ (.A(net6),
    .Z(_044_));
 INV_X1 _119_ (.A(_044_),
    .ZN(_045_));
 OAI21_X1 _120_ (.A(_045_),
    .B1(_032_),
    .B2(_033_),
    .ZN(_046_));
 NOR2_X2 _121_ (.A1(_028_),
    .A2(_021_),
    .ZN(_047_));
 NOR2_X1 _122_ (.A1(_039_),
    .A2(_047_),
    .ZN(_048_));
 NOR3_X1 _123_ (.A1(_023_),
    .A2(_042_),
    .A3(_048_),
    .ZN(_049_));
 OAI21_X1 _124_ (.A(_011_),
    .B1(_018_),
    .B2(_021_),
    .ZN(_050_));
 AOI21_X1 _125_ (.A(_031_),
    .B1(_050_),
    .B2(_035_),
    .ZN(_051_));
 OAI22_X1 _126_ (.A1(_032_),
    .A2(_022_),
    .B1(_051_),
    .B2(_038_),
    .ZN(_052_));
 OAI33_X1 _127_ (.A1(_037_),
    .A2(_043_),
    .A3(_046_),
    .B1(_049_),
    .B2(_052_),
    .B3(_045_),
    .ZN(net11));
 AOI21_X1 _128_ (.A(_044_),
    .B1(_039_),
    .B2(_033_),
    .ZN(_053_));
 NOR3_X1 _129_ (.A1(_039_),
    .A2(_018_),
    .A3(_022_),
    .ZN(_054_));
 OAI21_X1 _130_ (.A(_041_),
    .B1(_053_),
    .B2(_054_),
    .ZN(_055_));
 AOI21_X1 _131_ (.A(_044_),
    .B1(_011_),
    .B2(_022_),
    .ZN(_056_));
 NOR2_X2 _132_ (.A1(_017_),
    .A2(_033_),
    .ZN(_057_));
 AOI21_X1 _133_ (.A(_056_),
    .B1(_057_),
    .B2(_039_),
    .ZN(_058_));
 OAI221_X1 _134_ (.A(_055_),
    .B1(_058_),
    .B2(_041_),
    .C1(_044_),
    .C2(_018_),
    .ZN(_059_));
 NOR3_X1 _135_ (.A1(_032_),
    .A2(_028_),
    .A3(_033_),
    .ZN(_060_));
 OAI21_X1 _136_ (.A(_041_),
    .B1(_056_),
    .B2(_060_),
    .ZN(_061_));
 OAI21_X1 _137_ (.A(_061_),
    .B1(_028_),
    .B2(_044_),
    .ZN(_062_));
 AOI21_X1 _138_ (.A(_053_),
    .B1(_047_),
    .B2(_032_),
    .ZN(_063_));
 OAI21_X1 _139_ (.A(_023_),
    .B1(_041_),
    .B2(_063_),
    .ZN(_064_));
 OAI22_X1 _140_ (.A1(_023_),
    .A2(_059_),
    .B1(_062_),
    .B2(_064_),
    .ZN(net12));
 AOI21_X1 _141_ (.A(_041_),
    .B1(_011_),
    .B2(_028_),
    .ZN(_065_));
 AOI21_X1 _142_ (.A(_065_),
    .B1(_057_),
    .B2(_039_),
    .ZN(_066_));
 OAI22_X1 _143_ (.A1(_041_),
    .A2(_033_),
    .B1(_066_),
    .B2(_044_),
    .ZN(_067_));
 OAI21_X1 _144_ (.A(_035_),
    .B1(_032_),
    .B2(_028_),
    .ZN(_068_));
 NAND3_X1 _145_ (.A1(_032_),
    .A2(_018_),
    .A3(_022_),
    .ZN(_069_));
 AOI21_X1 _146_ (.A(_045_),
    .B1(_068_),
    .B2(_069_),
    .ZN(_070_));
 NOR3_X1 _147_ (.A1(_032_),
    .A2(_018_),
    .A3(_022_),
    .ZN(_071_));
 OAI21_X1 _148_ (.A(_044_),
    .B1(_065_),
    .B2(_071_),
    .ZN(_072_));
 INV_X1 _149_ (.A(_072_),
    .ZN(_073_));
 NAND2_X1 _150_ (.A1(_032_),
    .A2(_047_),
    .ZN(_074_));
 AOI21_X1 _151_ (.A(_044_),
    .B1(_074_),
    .B2(_068_),
    .ZN(_075_));
 OAI21_X1 _152_ (.A(_023_),
    .B1(_041_),
    .B2(_022_),
    .ZN(_076_));
 OAI33_X1 _153_ (.A1(_023_),
    .A2(_067_),
    .A3(_070_),
    .B1(_073_),
    .B2(_075_),
    .B3(_076_),
    .ZN(net13));
 OAI21_X1 _154_ (.A(_023_),
    .B1(_017_),
    .B2(_021_),
    .ZN(_077_));
 NAND3_X1 _155_ (.A1(_041_),
    .A2(_032_),
    .A3(_077_),
    .ZN(_078_));
 NOR2_X1 _156_ (.A1(_010_),
    .A2(_011_),
    .ZN(_079_));
 OR2_X1 _157_ (.A1(_028_),
    .A2(_079_),
    .ZN(_080_));
 AOI22_X1 _158_ (.A1(_057_),
    .A2(_079_),
    .B1(_080_),
    .B2(_038_),
    .ZN(_000_));
 AOI21_X1 _159_ (.A(_044_),
    .B1(_078_),
    .B2(_000_),
    .ZN(_001_));
 XNOR2_X1 _160_ (.A(_035_),
    .B(_022_),
    .ZN(_002_));
 NAND4_X1 _161_ (.A1(_035_),
    .A2(_011_),
    .A3(_018_),
    .A4(_022_),
    .ZN(_003_));
 NOR2_X1 _162_ (.A1(_038_),
    .A2(_047_),
    .ZN(_004_));
 NAND2_X1 _163_ (.A1(_041_),
    .A2(_039_),
    .ZN(_005_));
 AOI21_X1 _164_ (.A(_018_),
    .B1(_011_),
    .B2(_035_),
    .ZN(_006_));
 OAI221_X2 _165_ (.A(_003_),
    .B1(_004_),
    .B2(_005_),
    .C1(_006_),
    .C2(_023_),
    .ZN(_007_));
 AOI221_X2 _166_ (.A(_001_),
    .B1(_002_),
    .B2(_038_),
    .C1(_044_),
    .C2(_007_),
    .ZN(net14));
 XNOR2_X2 _167_ (.A(net4),
    .B(net2),
    .ZN(_008_));
 XNOR2_X1 _168_ (.A(net1),
    .B(_008_),
    .ZN(p1));
 XNOR2_X1 _169_ (.A(net1),
    .B(net3),
    .ZN(_009_));
 XNOR2_X1 _170_ (.A(net4),
    .B(_009_),
    .ZN(p2));
 XNOR2_X1 _171_ (.A(net3),
    .B(_008_),
    .ZN(p3));
 NAND2_X1 _172_ (.A1(_025_),
    .A2(_029_),
    .ZN(net26));
 BUF_X1 _173_ (.A(net10),
    .Z(net15));
 BUF_X1 _174_ (.A(net12),
    .Z(net16));
 BUF_X1 _175_ (.A(net13),
    .Z(net17));
 BUF_X1 _176_ (.A(net14),
    .Z(net18));
 BUF_X1 _177_ (.A(p1),
    .Z(net19));
 BUF_X1 _178_ (.A(p2),
    .Z(net20));
 BUF_X1 _179_ (.A(net1),
    .Z(net21));
 BUF_X1 _180_ (.A(p3),
    .Z(net22));
 BUF_X1 _181_ (.A(net2),
    .Z(net23));
 BUF_X1 _182_ (.A(net3),
    .Z(net24));
 BUF_X1 _183_ (.A(net4),
    .Z(net25));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[2]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[3]),
    .Z(net4));
 BUF_X2 input5 (.A(received_in[0]),
    .Z(net5));
 BUF_X1 input6 (.A(received_in[4]),
    .Z(net6));
 BUF_X1 input7 (.A(received_in[6]),
    .Z(net7));
 BUF_X1 output8 (.A(net8),
    .Z(corrected_code[0]));
 BUF_X1 output9 (.A(net9),
    .Z(corrected_code[1]));
 BUF_X1 output10 (.A(net10),
    .Z(corrected_code[2]));
 BUF_X1 output11 (.A(net11),
    .Z(corrected_code[3]));
 BUF_X1 output12 (.A(net12),
    .Z(corrected_code[4]));
 BUF_X1 output13 (.A(net13),
    .Z(corrected_code[5]));
 BUF_X1 output14 (.A(net14),
    .Z(corrected_code[6]));
 BUF_X1 output15 (.A(net15),
    .Z(data_out[0]));
 BUF_X1 output16 (.A(net16),
    .Z(data_out[1]));
 BUF_X1 output17 (.A(net17),
    .Z(data_out[2]));
 BUF_X1 output18 (.A(net18),
    .Z(data_out[3]));
 BUF_X1 output19 (.A(net19),
    .Z(encoded_out[0]));
 BUF_X1 output20 (.A(net20),
    .Z(encoded_out[1]));
 BUF_X1 output21 (.A(net21),
    .Z(encoded_out[2]));
 BUF_X1 output22 (.A(net22),
    .Z(encoded_out[3]));
 BUF_X1 output23 (.A(net23),
    .Z(encoded_out[4]));
 BUF_X1 output24 (.A(net24),
    .Z(encoded_out[5]));
 BUF_X1 output25 (.A(net25),
    .Z(encoded_out[6]));
 BUF_X1 output26 (.A(net26),
    .Z(single_bit_error));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X2 FILLER_0_33 ();
 FILLCELL_X1 FILLER_0_35 ();
 FILLCELL_X2 FILLER_0_63 ();
 FILLCELL_X4 FILLER_0_77 ();
 FILLCELL_X1 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X8 FILLER_0_89 ();
 FILLCELL_X1 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_110 ();
 FILLCELL_X32 FILLER_0_123 ();
 FILLCELL_X16 FILLER_0_155 ();
 FILLCELL_X8 FILLER_0_171 ();
 FILLCELL_X4 FILLER_0_179 ();
 FILLCELL_X1 FILLER_0_183 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X1 FILLER_1_33 ();
 FILLCELL_X2 FILLER_1_46 ();
 FILLCELL_X1 FILLER_1_48 ();
 FILLCELL_X16 FILLER_1_71 ();
 FILLCELL_X4 FILLER_1_87 ();
 FILLCELL_X2 FILLER_1_91 ();
 FILLCELL_X1 FILLER_1_93 ();
 FILLCELL_X2 FILLER_1_101 ();
 FILLCELL_X1 FILLER_1_103 ();
 FILLCELL_X32 FILLER_1_114 ();
 FILLCELL_X32 FILLER_1_146 ();
 FILLCELL_X4 FILLER_1_178 ();
 FILLCELL_X2 FILLER_1_182 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_41 ();
 FILLCELL_X1 FILLER_2_51 ();
 FILLCELL_X2 FILLER_2_58 ();
 FILLCELL_X16 FILLER_2_63 ();
 FILLCELL_X2 FILLER_2_79 ();
 FILLCELL_X1 FILLER_2_81 ();
 FILLCELL_X4 FILLER_2_85 ();
 FILLCELL_X32 FILLER_2_98 ();
 FILLCELL_X32 FILLER_2_130 ();
 FILLCELL_X16 FILLER_2_162 ();
 FILLCELL_X4 FILLER_2_178 ();
 FILLCELL_X2 FILLER_2_182 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X16 FILLER_3_65 ();
 FILLCELL_X2 FILLER_3_81 ();
 FILLCELL_X32 FILLER_3_96 ();
 FILLCELL_X32 FILLER_3_128 ();
 FILLCELL_X16 FILLER_3_160 ();
 FILLCELL_X8 FILLER_3_176 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X16 FILLER_4_161 ();
 FILLCELL_X4 FILLER_4_177 ();
 FILLCELL_X2 FILLER_4_181 ();
 FILLCELL_X1 FILLER_4_183 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X2 FILLER_5_81 ();
 FILLCELL_X1 FILLER_5_83 ();
 FILLCELL_X8 FILLER_5_90 ();
 FILLCELL_X4 FILLER_5_98 ();
 FILLCELL_X1 FILLER_5_102 ();
 FILLCELL_X32 FILLER_5_112 ();
 FILLCELL_X32 FILLER_5_144 ();
 FILLCELL_X8 FILLER_5_176 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X2 FILLER_6_73 ();
 FILLCELL_X1 FILLER_6_75 ();
 FILLCELL_X8 FILLER_6_83 ();
 FILLCELL_X2 FILLER_6_91 ();
 FILLCELL_X32 FILLER_6_122 ();
 FILLCELL_X16 FILLER_6_154 ();
 FILLCELL_X8 FILLER_6_170 ();
 FILLCELL_X4 FILLER_6_178 ();
 FILLCELL_X2 FILLER_6_182 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_73 ();
 FILLCELL_X2 FILLER_7_77 ();
 FILLCELL_X32 FILLER_7_86 ();
 FILLCELL_X32 FILLER_7_118 ();
 FILLCELL_X32 FILLER_7_150 ();
 FILLCELL_X2 FILLER_7_182 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X2 FILLER_8_65 ();
 FILLCELL_X16 FILLER_8_74 ();
 FILLCELL_X4 FILLER_8_90 ();
 FILLCELL_X2 FILLER_8_94 ();
 FILLCELL_X1 FILLER_8_96 ();
 FILLCELL_X32 FILLER_8_111 ();
 FILLCELL_X32 FILLER_8_143 ();
 FILLCELL_X8 FILLER_8_175 ();
 FILLCELL_X1 FILLER_8_183 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X4 FILLER_9_25 ();
 FILLCELL_X2 FILLER_9_29 ();
 FILLCELL_X16 FILLER_9_34 ();
 FILLCELL_X4 FILLER_9_50 ();
 FILLCELL_X8 FILLER_9_71 ();
 FILLCELL_X1 FILLER_9_79 ();
 FILLCELL_X4 FILLER_9_90 ();
 FILLCELL_X2 FILLER_9_94 ();
 FILLCELL_X8 FILLER_9_108 ();
 FILLCELL_X2 FILLER_9_116 ();
 FILLCELL_X4 FILLER_9_122 ();
 FILLCELL_X2 FILLER_9_126 ();
 FILLCELL_X1 FILLER_9_128 ();
 FILLCELL_X32 FILLER_9_133 ();
 FILLCELL_X16 FILLER_9_165 ();
 FILLCELL_X2 FILLER_9_181 ();
 FILLCELL_X1 FILLER_9_183 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_3 ();
 FILLCELL_X32 FILLER_10_7 ();
 FILLCELL_X16 FILLER_10_39 ();
 FILLCELL_X8 FILLER_10_55 ();
 FILLCELL_X2 FILLER_10_63 ();
 FILLCELL_X1 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_73 ();
 FILLCELL_X2 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_91 ();
 FILLCELL_X4 FILLER_10_97 ();
 FILLCELL_X1 FILLER_10_101 ();
 FILLCELL_X4 FILLER_10_106 ();
 FILLCELL_X2 FILLER_10_110 ();
 FILLCELL_X1 FILLER_10_112 ();
 FILLCELL_X1 FILLER_10_117 ();
 FILLCELL_X1 FILLER_10_122 ();
 FILLCELL_X1 FILLER_10_127 ();
 FILLCELL_X1 FILLER_10_132 ();
 FILLCELL_X32 FILLER_10_137 ();
 FILLCELL_X8 FILLER_10_169 ();
 FILLCELL_X4 FILLER_10_177 ();
 FILLCELL_X2 FILLER_10_181 ();
 FILLCELL_X1 FILLER_10_183 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X16 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_81 ();
 FILLCELL_X4 FILLER_11_89 ();
 FILLCELL_X2 FILLER_11_93 ();
 FILLCELL_X8 FILLER_11_104 ();
 FILLCELL_X4 FILLER_11_112 ();
 FILLCELL_X1 FILLER_11_116 ();
 FILLCELL_X8 FILLER_11_121 ();
 FILLCELL_X1 FILLER_11_129 ();
 FILLCELL_X2 FILLER_11_144 ();
 FILLCELL_X1 FILLER_11_146 ();
 FILLCELL_X16 FILLER_11_152 ();
 FILLCELL_X8 FILLER_11_168 ();
 FILLCELL_X2 FILLER_11_182 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X16 FILLER_12_65 ();
 FILLCELL_X1 FILLER_12_81 ();
 FILLCELL_X16 FILLER_12_85 ();
 FILLCELL_X8 FILLER_12_101 ();
 FILLCELL_X2 FILLER_12_109 ();
 FILLCELL_X32 FILLER_12_115 ();
 FILLCELL_X16 FILLER_12_147 ();
 FILLCELL_X8 FILLER_12_163 ();
 FILLCELL_X4 FILLER_12_171 ();
 FILLCELL_X2 FILLER_12_175 ();
 FILLCELL_X1 FILLER_12_177 ();
 FILLCELL_X2 FILLER_12_181 ();
 FILLCELL_X1 FILLER_12_183 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_38 ();
 FILLCELL_X4 FILLER_13_70 ();
 FILLCELL_X2 FILLER_13_74 ();
 FILLCELL_X1 FILLER_13_76 ();
 FILLCELL_X2 FILLER_13_88 ();
 FILLCELL_X8 FILLER_13_94 ();
 FILLCELL_X4 FILLER_13_113 ();
 FILLCELL_X2 FILLER_13_117 ();
 FILLCELL_X2 FILLER_13_123 ();
 FILLCELL_X1 FILLER_13_133 ();
 FILLCELL_X32 FILLER_13_138 ();
 FILLCELL_X8 FILLER_13_170 ();
 FILLCELL_X4 FILLER_13_178 ();
 FILLCELL_X2 FILLER_13_182 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X8 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_76 ();
 FILLCELL_X4 FILLER_14_92 ();
 FILLCELL_X2 FILLER_14_96 ();
 FILLCELL_X1 FILLER_14_101 ();
 FILLCELL_X1 FILLER_14_107 ();
 FILLCELL_X4 FILLER_14_111 ();
 FILLCELL_X2 FILLER_14_115 ();
 FILLCELL_X1 FILLER_14_117 ();
 FILLCELL_X2 FILLER_14_122 ();
 FILLCELL_X1 FILLER_14_124 ();
 FILLCELL_X4 FILLER_14_130 ();
 FILLCELL_X1 FILLER_14_134 ();
 FILLCELL_X32 FILLER_14_137 ();
 FILLCELL_X8 FILLER_14_169 ();
 FILLCELL_X4 FILLER_14_177 ();
 FILLCELL_X2 FILLER_14_181 ();
 FILLCELL_X1 FILLER_14_183 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X4 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_69 ();
 FILLCELL_X4 FILLER_15_77 ();
 FILLCELL_X4 FILLER_15_85 ();
 FILLCELL_X1 FILLER_15_97 ();
 FILLCELL_X1 FILLER_15_102 ();
 FILLCELL_X1 FILLER_15_110 ();
 FILLCELL_X8 FILLER_15_115 ();
 FILLCELL_X2 FILLER_15_123 ();
 FILLCELL_X1 FILLER_15_125 ();
 FILLCELL_X2 FILLER_15_132 ();
 FILLCELL_X1 FILLER_15_137 ();
 FILLCELL_X32 FILLER_15_142 ();
 FILLCELL_X4 FILLER_15_174 ();
 FILLCELL_X2 FILLER_15_181 ();
 FILLCELL_X1 FILLER_15_183 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X4 FILLER_16_65 ();
 FILLCELL_X2 FILLER_16_80 ();
 FILLCELL_X1 FILLER_16_93 ();
 FILLCELL_X2 FILLER_16_97 ();
 FILLCELL_X2 FILLER_16_103 ();
 FILLCELL_X1 FILLER_16_105 ();
 FILLCELL_X16 FILLER_16_113 ();
 FILLCELL_X1 FILLER_16_129 ();
 FILLCELL_X1 FILLER_16_134 ();
 FILLCELL_X2 FILLER_16_139 ();
 FILLCELL_X16 FILLER_16_148 ();
 FILLCELL_X8 FILLER_16_164 ();
 FILLCELL_X2 FILLER_16_172 ();
 FILLCELL_X1 FILLER_16_174 ();
 FILLCELL_X2 FILLER_16_178 ();
 FILLCELL_X1 FILLER_16_180 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X4 FILLER_17_97 ();
 FILLCELL_X2 FILLER_17_101 ();
 FILLCELL_X32 FILLER_17_108 ();
 FILLCELL_X32 FILLER_17_140 ();
 FILLCELL_X8 FILLER_17_172 ();
 FILLCELL_X4 FILLER_17_180 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_70 ();
 FILLCELL_X32 FILLER_18_102 ();
 FILLCELL_X32 FILLER_18_134 ();
 FILLCELL_X16 FILLER_18_166 ();
 FILLCELL_X2 FILLER_18_182 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_177 ();
 FILLCELL_X2 FILLER_19_181 ();
 FILLCELL_X1 FILLER_19_183 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_177 ();
 FILLCELL_X2 FILLER_20_181 ();
 FILLCELL_X1 FILLER_20_183 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_177 ();
 FILLCELL_X2 FILLER_21_181 ();
 FILLCELL_X1 FILLER_21_183 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X16 FILLER_22_33 ();
 FILLCELL_X8 FILLER_22_49 ();
 FILLCELL_X4 FILLER_22_57 ();
 FILLCELL_X2 FILLER_22_61 ();
 FILLCELL_X32 FILLER_22_69 ();
 FILLCELL_X32 FILLER_22_101 ();
 FILLCELL_X32 FILLER_22_133 ();
 FILLCELL_X16 FILLER_22_165 ();
 FILLCELL_X2 FILLER_22_181 ();
 FILLCELL_X1 FILLER_22_183 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_68 ();
 FILLCELL_X8 FILLER_23_100 ();
 FILLCELL_X32 FILLER_23_111 ();
 FILLCELL_X32 FILLER_23_143 ();
 FILLCELL_X8 FILLER_23_175 ();
 FILLCELL_X1 FILLER_23_183 ();
endmodule
