module parameterized_gray_counter (clk,
    enable,
    rst_n,
    binary_out,
    gray_out);
 input clk;
 input enable;
 input rst_n;
 output [3:0] binary_out;
 output [3:0] gray_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _17_ (.A(enable),
    .Z(_05_));
 MUX2_X1 _18_ (.A(net2),
    .B(_00_),
    .S(_05_),
    .Z(_06_));
 AND2_X1 _19_ (.A1(net1),
    .A2(_06_),
    .ZN(_01_));
 MUX2_X1 _20_ (.A(net3),
    .B(net6),
    .S(_05_),
    .Z(_07_));
 AND2_X1 _21_ (.A1(net1),
    .A2(_07_),
    .ZN(_02_));
 NAND2_X1 _22_ (.A1(_15_),
    .A2(_05_),
    .ZN(_08_));
 XNOR2_X1 _23_ (.A(net4),
    .B(_08_),
    .ZN(_09_));
 AND2_X1 _24_ (.A1(net1),
    .A2(_09_),
    .ZN(_03_));
 NAND3_X1 _25_ (.A1(net2),
    .A2(_16_),
    .A3(_05_),
    .ZN(_10_));
 XNOR2_X1 _26_ (.A(net5),
    .B(_10_),
    .ZN(_11_));
 AND2_X1 _27_ (.A1(net1),
    .A2(_11_),
    .ZN(_04_));
 XOR2_X1 _28_ (.A(net4),
    .B(net5),
    .Z(net8));
 HA_X1 _29_ (.A(net2),
    .B(net3),
    .CO(_15_),
    .S(net6));
 HA_X1 _30_ (.A(net3),
    .B(net4),
    .CO(_16_),
    .S(net7));
 BUF_X1 _31_ (.A(net5),
    .Z(net9));
 DFF_X2 \binary_count[0]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_00_));
 DFF_X2 \binary_count[1]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net3),
    .QN(_14_));
 DFF_X2 \binary_count[2]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_13_));
 DFF_X1 \binary_count[3]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_12_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_53 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(binary_out[0]));
 BUF_X1 output3 (.A(net3),
    .Z(binary_out[1]));
 BUF_X1 output4 (.A(net4),
    .Z(binary_out[2]));
 BUF_X1 output5 (.A(net5),
    .Z(binary_out[3]));
 BUF_X1 output6 (.A(net6),
    .Z(gray_out[0]));
 BUF_X1 output7 (.A(net7),
    .Z(gray_out[1]));
 BUF_X1 output8 (.A(net8),
    .Z(gray_out[2]));
 BUF_X1 output9 (.A(net9),
    .Z(gray_out[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X1 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X1 FILLER_0_103 ();
 FILLCELL_X32 FILLER_0_107 ();
 FILLCELL_X32 FILLER_0_139 ();
 FILLCELL_X32 FILLER_0_171 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_100 ();
 FILLCELL_X32 FILLER_1_132 ();
 FILLCELL_X32 FILLER_1_164 ();
 FILLCELL_X4 FILLER_1_196 ();
 FILLCELL_X2 FILLER_1_200 ();
 FILLCELL_X1 FILLER_1_202 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X8 FILLER_2_193 ();
 FILLCELL_X2 FILLER_2_201 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X8 FILLER_3_193 ();
 FILLCELL_X2 FILLER_3_201 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X8 FILLER_4_193 ();
 FILLCELL_X2 FILLER_4_201 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X8 FILLER_5_193 ();
 FILLCELL_X2 FILLER_5_201 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X8 FILLER_6_193 ();
 FILLCELL_X2 FILLER_6_201 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X8 FILLER_7_193 ();
 FILLCELL_X2 FILLER_7_201 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X8 FILLER_8_193 ();
 FILLCELL_X2 FILLER_8_201 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X8 FILLER_9_193 ();
 FILLCELL_X2 FILLER_9_201 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X8 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_112 ();
 FILLCELL_X32 FILLER_10_144 ();
 FILLCELL_X16 FILLER_10_176 ();
 FILLCELL_X8 FILLER_10_192 ();
 FILLCELL_X2 FILLER_10_200 ();
 FILLCELL_X1 FILLER_10_202 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X16 FILLER_11_65 ();
 FILLCELL_X8 FILLER_11_81 ();
 FILLCELL_X4 FILLER_11_89 ();
 FILLCELL_X2 FILLER_11_93 ();
 FILLCELL_X1 FILLER_11_95 ();
 FILLCELL_X32 FILLER_11_113 ();
 FILLCELL_X32 FILLER_11_145 ();
 FILLCELL_X16 FILLER_11_177 ();
 FILLCELL_X8 FILLER_11_193 ();
 FILLCELL_X2 FILLER_11_201 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X16 FILLER_12_65 ();
 FILLCELL_X4 FILLER_12_81 ();
 FILLCELL_X32 FILLER_12_111 ();
 FILLCELL_X32 FILLER_12_143 ();
 FILLCELL_X16 FILLER_12_175 ();
 FILLCELL_X8 FILLER_12_191 ();
 FILLCELL_X4 FILLER_12_199 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X16 FILLER_13_65 ();
 FILLCELL_X8 FILLER_13_81 ();
 FILLCELL_X2 FILLER_13_89 ();
 FILLCELL_X32 FILLER_13_121 ();
 FILLCELL_X32 FILLER_13_153 ();
 FILLCELL_X16 FILLER_13_185 ();
 FILLCELL_X2 FILLER_13_201 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X16 FILLER_14_65 ();
 FILLCELL_X8 FILLER_14_81 ();
 FILLCELL_X4 FILLER_14_89 ();
 FILLCELL_X2 FILLER_14_93 ();
 FILLCELL_X1 FILLER_14_113 ();
 FILLCELL_X32 FILLER_14_120 ();
 FILLCELL_X32 FILLER_14_152 ();
 FILLCELL_X16 FILLER_14_184 ();
 FILLCELL_X2 FILLER_14_200 ();
 FILLCELL_X1 FILLER_14_202 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X16 FILLER_15_65 ();
 FILLCELL_X8 FILLER_15_81 ();
 FILLCELL_X2 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_91 ();
 FILLCELL_X32 FILLER_15_119 ();
 FILLCELL_X32 FILLER_15_151 ();
 FILLCELL_X16 FILLER_15_183 ();
 FILLCELL_X4 FILLER_15_199 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X8 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_201 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X8 FILLER_17_193 ();
 FILLCELL_X2 FILLER_17_201 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X2 FILLER_18_97 ();
 FILLCELL_X1 FILLER_18_99 ();
 FILLCELL_X32 FILLER_18_105 ();
 FILLCELL_X32 FILLER_18_137 ();
 FILLCELL_X32 FILLER_18_169 ();
 FILLCELL_X2 FILLER_18_201 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X8 FILLER_19_193 ();
 FILLCELL_X2 FILLER_19_201 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X8 FILLER_20_193 ();
 FILLCELL_X2 FILLER_20_201 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X8 FILLER_21_193 ();
 FILLCELL_X2 FILLER_21_201 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X8 FILLER_22_193 ();
 FILLCELL_X2 FILLER_22_201 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X4 FILLER_23_97 ();
 FILLCELL_X1 FILLER_23_101 ();
 FILLCELL_X1 FILLER_23_106 ();
 FILLCELL_X32 FILLER_23_118 ();
 FILLCELL_X32 FILLER_23_150 ();
 FILLCELL_X16 FILLER_23_182 ();
 FILLCELL_X4 FILLER_23_198 ();
 FILLCELL_X1 FILLER_23_202 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X16 FILLER_24_65 ();
 FILLCELL_X8 FILLER_24_81 ();
 FILLCELL_X4 FILLER_24_89 ();
 FILLCELL_X32 FILLER_24_110 ();
 FILLCELL_X32 FILLER_24_142 ();
 FILLCELL_X16 FILLER_24_174 ();
 FILLCELL_X8 FILLER_24_190 ();
 FILLCELL_X4 FILLER_24_198 ();
 FILLCELL_X1 FILLER_24_202 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X16 FILLER_25_65 ();
 FILLCELL_X8 FILLER_25_81 ();
 FILLCELL_X4 FILLER_25_89 ();
 FILLCELL_X1 FILLER_25_93 ();
 FILLCELL_X2 FILLER_25_97 ();
 FILLCELL_X2 FILLER_25_102 ();
 FILLCELL_X1 FILLER_25_104 ();
 FILLCELL_X32 FILLER_25_114 ();
 FILLCELL_X32 FILLER_25_146 ();
 FILLCELL_X16 FILLER_25_178 ();
 FILLCELL_X8 FILLER_25_194 ();
 FILLCELL_X1 FILLER_25_202 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X4 FILLER_26_97 ();
 FILLCELL_X2 FILLER_26_104 ();
 FILLCELL_X1 FILLER_26_109 ();
 FILLCELL_X32 FILLER_26_116 ();
 FILLCELL_X32 FILLER_26_148 ();
 FILLCELL_X16 FILLER_26_180 ();
 FILLCELL_X4 FILLER_26_196 ();
 FILLCELL_X2 FILLER_26_200 ();
 FILLCELL_X1 FILLER_26_202 ();
endmodule
