module leading_zero_counter (valid_input,
    data_in,
    zero_count);
 output valid_input;
 input [31:0] data_in;
 output [5:0] zero_count;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;

 NOR4_X2 _067_ (.A1(net31),
    .A2(net30),
    .A3(net3),
    .A4(net2),
    .ZN(_011_));
 NOR4_X2 _068_ (.A1(net5),
    .A2(net4),
    .A3(net7),
    .A4(net6),
    .ZN(_012_));
 NAND2_X1 _069_ (.A1(_011_),
    .A2(_012_),
    .ZN(_013_));
 NOR4_X2 _070_ (.A1(net25),
    .A2(net22),
    .A3(net29),
    .A4(net28),
    .ZN(_014_));
 NOR2_X1 _071_ (.A1(net12),
    .A2(net1),
    .ZN(_015_));
 NOR2_X1 _072_ (.A1(net27),
    .A2(net26),
    .ZN(_016_));
 NAND3_X1 _073_ (.A1(_014_),
    .A2(_015_),
    .A3(_016_),
    .ZN(_017_));
 OR2_X1 _074_ (.A1(_013_),
    .A2(_017_),
    .ZN(net37));
 INV_X1 _075_ (.A(net37),
    .ZN(_018_));
 NOR4_X1 _076_ (.A1(net9),
    .A2(net8),
    .A3(net11),
    .A4(net10),
    .ZN(_019_));
 BUF_X1 _077_ (.A(data_in[20]),
    .Z(_020_));
 NOR2_X1 _078_ (.A1(net13),
    .A2(_020_),
    .ZN(_021_));
 NOR2_X1 _079_ (.A1(net15),
    .A2(net14),
    .ZN(_022_));
 AND3_X1 _080_ (.A1(_019_),
    .A2(_021_),
    .A3(_022_),
    .ZN(_023_));
 NOR4_X2 _081_ (.A1(net17),
    .A2(net16),
    .A3(net19),
    .A4(net18),
    .ZN(_024_));
 NOR4_X1 _082_ (.A1(net21),
    .A2(net20),
    .A3(net24),
    .A4(net23),
    .ZN(_025_));
 AND4_X1 _083_ (.A1(_018_),
    .A2(_023_),
    .A3(_024_),
    .A4(_025_),
    .ZN(net38));
 NAND4_X1 _084_ (.A1(_018_),
    .A2(_023_),
    .A3(_024_),
    .A4(_025_),
    .ZN(net32));
 INV_X1 _085_ (.A(net22),
    .ZN(_026_));
 AOI21_X1 _086_ (.A(net12),
    .B1(net25),
    .B2(_026_),
    .ZN(_027_));
 NOR3_X1 _087_ (.A1(net1),
    .A2(net22),
    .A3(net26),
    .ZN(_028_));
 INV_X1 _088_ (.A(net29),
    .ZN(_029_));
 AOI21_X1 _089_ (.A(net28),
    .B1(net30),
    .B2(_029_),
    .ZN(_030_));
 OAI21_X1 _090_ (.A(_028_),
    .B1(_030_),
    .B2(net27),
    .ZN(_031_));
 OR3_X1 _091_ (.A1(net27),
    .A2(net29),
    .A3(net31),
    .ZN(_032_));
 INV_X1 _092_ (.A(net3),
    .ZN(_033_));
 INV_X1 _093_ (.A(net5),
    .ZN(_034_));
 OAI21_X1 _094_ (.A(_033_),
    .B1(_034_),
    .B2(net4),
    .ZN(_035_));
 INV_X1 _095_ (.A(net2),
    .ZN(_036_));
 AOI21_X1 _096_ (.A(_032_),
    .B1(_035_),
    .B2(_036_),
    .ZN(_037_));
 OAI22_X1 _097_ (.A1(net1),
    .A2(_027_),
    .B1(_031_),
    .B2(_037_),
    .ZN(_038_));
 NOR3_X1 _098_ (.A1(net2),
    .A2(net4),
    .A3(net6),
    .ZN(_039_));
 INV_X1 _099_ (.A(net9),
    .ZN(_040_));
 AOI21_X1 _100_ (.A(net8),
    .B1(net10),
    .B2(_040_),
    .ZN(_041_));
 OAI21_X1 _101_ (.A(_039_),
    .B1(_041_),
    .B2(net7),
    .ZN(_042_));
 NOR2_X1 _102_ (.A1(_031_),
    .A2(_042_),
    .ZN(_043_));
 OR3_X1 _103_ (.A1(net7),
    .A2(net9),
    .A3(net11),
    .ZN(_044_));
 NOR2_X1 _104_ (.A1(_020_),
    .A2(net14),
    .ZN(_045_));
 INV_X1 _105_ (.A(_020_),
    .ZN(_046_));
 AOI221_X2 _106_ (.A(_044_),
    .B1(_045_),
    .B2(net15),
    .C1(net13),
    .C2(_046_),
    .ZN(_047_));
 OR3_X1 _107_ (.A1(_020_),
    .A2(net14),
    .A3(net16),
    .ZN(_048_));
 INV_X1 _108_ (.A(net18),
    .ZN(_049_));
 INV_X1 _109_ (.A(net21),
    .ZN(_050_));
 NAND2_X1 _110_ (.A1(_050_),
    .A2(net23),
    .ZN(_051_));
 NOR2_X1 _111_ (.A1(net18),
    .A2(net20),
    .ZN(_052_));
 AOI221_X2 _112_ (.A(net17),
    .B1(net19),
    .B2(_049_),
    .C1(_051_),
    .C2(_052_),
    .ZN(_053_));
 OAI21_X1 _113_ (.A(_047_),
    .B1(_048_),
    .B2(_053_),
    .ZN(_054_));
 AOI21_X1 _114_ (.A(_038_),
    .B1(_043_),
    .B2(_054_),
    .ZN(net33));
 INV_X1 _115_ (.A(net8),
    .ZN(_055_));
 NOR2_X1 _116_ (.A1(net5),
    .A2(net4),
    .ZN(_056_));
 NAND3_X1 _117_ (.A1(_040_),
    .A2(_055_),
    .A3(_056_),
    .ZN(_057_));
 NOR3_X1 _118_ (.A1(net13),
    .A2(_020_),
    .A3(_022_),
    .ZN(_058_));
 NOR3_X1 _119_ (.A1(net11),
    .A2(net10),
    .A3(_058_),
    .ZN(_059_));
 NOR2_X1 _120_ (.A1(net17),
    .A2(net16),
    .ZN(_060_));
 NOR2_X1 _121_ (.A1(net19),
    .A2(net18),
    .ZN(_061_));
 OAI21_X1 _122_ (.A(_061_),
    .B1(net20),
    .B2(net21),
    .ZN(_062_));
 NAND3_X1 _123_ (.A1(_021_),
    .A2(_060_),
    .A3(_062_),
    .ZN(_063_));
 AOI21_X1 _124_ (.A(_057_),
    .B1(_059_),
    .B2(_063_),
    .ZN(_064_));
 OAI21_X1 _125_ (.A(_056_),
    .B1(net6),
    .B2(net7),
    .ZN(_065_));
 NAND4_X1 _126_ (.A1(_033_),
    .A2(_036_),
    .A3(_014_),
    .A4(_065_),
    .ZN(_066_));
 NOR2_X1 _127_ (.A1(net29),
    .A2(net28),
    .ZN(_000_));
 OAI21_X1 _128_ (.A(_000_),
    .B1(net30),
    .B2(net31),
    .ZN(_001_));
 AND2_X1 _129_ (.A1(_016_),
    .A2(_001_),
    .ZN(_002_));
 OR2_X1 _130_ (.A1(net25),
    .A2(net22),
    .ZN(_003_));
 OAI221_X1 _131_ (.A(_015_),
    .B1(_064_),
    .B2(_066_),
    .C1(_002_),
    .C2(_003_),
    .ZN(net34));
 INV_X1 _132_ (.A(net28),
    .ZN(_004_));
 NAND3_X1 _133_ (.A1(_029_),
    .A2(_004_),
    .A3(_016_),
    .ZN(_005_));
 OR4_X1 _134_ (.A1(net13),
    .A2(_020_),
    .A3(net15),
    .A4(net14),
    .ZN(_006_));
 OAI21_X1 _135_ (.A(_019_),
    .B1(_006_),
    .B2(_024_),
    .ZN(_007_));
 NAND2_X1 _136_ (.A1(_012_),
    .A2(_007_),
    .ZN(_008_));
 AOI21_X1 _137_ (.A(_005_),
    .B1(_008_),
    .B2(_011_),
    .ZN(_009_));
 OR4_X1 _138_ (.A1(net12),
    .A2(net1),
    .A3(_003_),
    .A4(_009_),
    .ZN(net35));
 INV_X1 _139_ (.A(_017_),
    .ZN(_010_));
 OAI21_X1 _140_ (.A(_010_),
    .B1(_023_),
    .B2(_013_),
    .ZN(net36));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_55 ();
 BUF_X1 input1 (.A(data_in[0]),
    .Z(net1));
 BUF_X1 input2 (.A(data_in[10]),
    .Z(net2));
 BUF_X1 input3 (.A(data_in[11]),
    .Z(net3));
 BUF_X1 input4 (.A(data_in[12]),
    .Z(net4));
 BUF_X1 input5 (.A(data_in[13]),
    .Z(net5));
 BUF_X1 input6 (.A(data_in[14]),
    .Z(net6));
 BUF_X1 input7 (.A(data_in[15]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[16]),
    .Z(net8));
 BUF_X1 input9 (.A(data_in[17]),
    .Z(net9));
 BUF_X1 input10 (.A(data_in[18]),
    .Z(net10));
 BUF_X1 input11 (.A(data_in[19]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[1]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[21]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[22]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[23]),
    .Z(net15));
 BUF_X1 input16 (.A(data_in[24]),
    .Z(net16));
 BUF_X1 input17 (.A(data_in[25]),
    .Z(net17));
 BUF_X1 input18 (.A(data_in[26]),
    .Z(net18));
 BUF_X1 input19 (.A(data_in[27]),
    .Z(net19));
 BUF_X1 input20 (.A(data_in[28]),
    .Z(net20));
 BUF_X1 input21 (.A(data_in[29]),
    .Z(net21));
 BUF_X1 input22 (.A(data_in[2]),
    .Z(net22));
 BUF_X1 input23 (.A(data_in[30]),
    .Z(net23));
 BUF_X1 input24 (.A(data_in[31]),
    .Z(net24));
 BUF_X1 input25 (.A(data_in[3]),
    .Z(net25));
 BUF_X1 input26 (.A(data_in[4]),
    .Z(net26));
 BUF_X1 input27 (.A(data_in[5]),
    .Z(net27));
 CLKBUF_X2 input28 (.A(data_in[6]),
    .Z(net28));
 BUF_X1 input29 (.A(data_in[7]),
    .Z(net29));
 BUF_X1 input30 (.A(data_in[8]),
    .Z(net30));
 BUF_X1 input31 (.A(data_in[9]),
    .Z(net31));
 BUF_X1 output32 (.A(net32),
    .Z(valid_input));
 BUF_X1 output33 (.A(net33),
    .Z(zero_count[0]));
 BUF_X1 output34 (.A(net34),
    .Z(zero_count[1]));
 BUF_X1 output35 (.A(net35),
    .Z(zero_count[2]));
 BUF_X1 output36 (.A(net36),
    .Z(zero_count[3]));
 BUF_X1 output37 (.A(net37),
    .Z(zero_count[4]));
 BUF_X1 output38 (.A(net38),
    .Z(zero_count[5]));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_94 ();
 FILLCELL_X2 FILLER_0_101 ();
 FILLCELL_X32 FILLER_0_121 ();
 FILLCELL_X32 FILLER_0_153 ();
 FILLCELL_X16 FILLER_0_185 ();
 FILLCELL_X8 FILLER_0_201 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_81 ();
 FILLCELL_X2 FILLER_1_85 ();
 FILLCELL_X1 FILLER_1_87 ();
 FILLCELL_X1 FILLER_1_111 ();
 FILLCELL_X32 FILLER_1_117 ();
 FILLCELL_X32 FILLER_1_149 ();
 FILLCELL_X16 FILLER_1_181 ();
 FILLCELL_X8 FILLER_1_197 ();
 FILLCELL_X4 FILLER_1_205 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X16 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_81 ();
 FILLCELL_X32 FILLER_2_94 ();
 FILLCELL_X32 FILLER_2_126 ();
 FILLCELL_X32 FILLER_2_158 ();
 FILLCELL_X16 FILLER_2_190 ();
 FILLCELL_X2 FILLER_2_206 ();
 FILLCELL_X1 FILLER_2_208 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_105 ();
 FILLCELL_X1 FILLER_3_109 ();
 FILLCELL_X32 FILLER_3_121 ();
 FILLCELL_X32 FILLER_3_153 ();
 FILLCELL_X16 FILLER_3_185 ();
 FILLCELL_X8 FILLER_3_201 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X16 FILLER_4_193 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X16 FILLER_5_193 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X16 FILLER_6_193 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X16 FILLER_7_193 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_65 ();
 FILLCELL_X4 FILLER_8_81 ();
 FILLCELL_X1 FILLER_8_85 ();
 FILLCELL_X32 FILLER_8_89 ();
 FILLCELL_X32 FILLER_8_121 ();
 FILLCELL_X32 FILLER_8_153 ();
 FILLCELL_X16 FILLER_8_185 ();
 FILLCELL_X8 FILLER_8_201 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X1 FILLER_9_85 ();
 FILLCELL_X32 FILLER_9_90 ();
 FILLCELL_X32 FILLER_9_122 ();
 FILLCELL_X32 FILLER_9_154 ();
 FILLCELL_X16 FILLER_9_186 ();
 FILLCELL_X4 FILLER_9_202 ();
 FILLCELL_X2 FILLER_9_206 ();
 FILLCELL_X1 FILLER_9_208 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X16 FILLER_10_97 ();
 FILLCELL_X8 FILLER_10_113 ();
 FILLCELL_X32 FILLER_10_123 ();
 FILLCELL_X32 FILLER_10_155 ();
 FILLCELL_X16 FILLER_10_187 ();
 FILLCELL_X4 FILLER_10_203 ();
 FILLCELL_X2 FILLER_10_207 ();
 FILLCELL_X16 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_17 ();
 FILLCELL_X4 FILLER_11_25 ();
 FILLCELL_X2 FILLER_11_29 ();
 FILLCELL_X1 FILLER_11_31 ();
 FILLCELL_X2 FILLER_11_35 ();
 FILLCELL_X32 FILLER_11_40 ();
 FILLCELL_X2 FILLER_11_72 ();
 FILLCELL_X1 FILLER_11_74 ();
 FILLCELL_X2 FILLER_11_78 ();
 FILLCELL_X2 FILLER_11_82 ();
 FILLCELL_X1 FILLER_11_84 ();
 FILLCELL_X32 FILLER_11_90 ();
 FILLCELL_X32 FILLER_11_122 ();
 FILLCELL_X16 FILLER_11_154 ();
 FILLCELL_X32 FILLER_11_173 ();
 FILLCELL_X4 FILLER_11_205 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_17 ();
 FILLCELL_X2 FILLER_12_21 ();
 FILLCELL_X4 FILLER_12_26 ();
 FILLCELL_X1 FILLER_12_30 ();
 FILLCELL_X32 FILLER_12_34 ();
 FILLCELL_X4 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_73 ();
 FILLCELL_X2 FILLER_12_91 ();
 FILLCELL_X1 FILLER_12_93 ();
 FILLCELL_X32 FILLER_12_98 ();
 FILLCELL_X32 FILLER_12_130 ();
 FILLCELL_X16 FILLER_12_162 ();
 FILLCELL_X16 FILLER_12_181 ();
 FILLCELL_X8 FILLER_12_197 ();
 FILLCELL_X4 FILLER_12_205 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X4 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_69 ();
 FILLCELL_X8 FILLER_13_74 ();
 FILLCELL_X2 FILLER_13_82 ();
 FILLCELL_X2 FILLER_13_87 ();
 FILLCELL_X2 FILLER_13_94 ();
 FILLCELL_X16 FILLER_13_100 ();
 FILLCELL_X1 FILLER_13_116 ();
 FILLCELL_X32 FILLER_13_127 ();
 FILLCELL_X32 FILLER_13_159 ();
 FILLCELL_X16 FILLER_13_191 ();
 FILLCELL_X2 FILLER_13_207 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X16 FILLER_14_193 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_5 ();
 FILLCELL_X8 FILLER_15_9 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_21 ();
 FILLCELL_X1 FILLER_15_25 ();
 FILLCELL_X32 FILLER_15_29 ();
 FILLCELL_X8 FILLER_15_61 ();
 FILLCELL_X2 FILLER_15_69 ();
 FILLCELL_X1 FILLER_15_71 ();
 FILLCELL_X8 FILLER_15_76 ();
 FILLCELL_X4 FILLER_15_84 ();
 FILLCELL_X8 FILLER_15_92 ();
 FILLCELL_X1 FILLER_15_100 ();
 FILLCELL_X8 FILLER_15_104 ();
 FILLCELL_X4 FILLER_15_112 ();
 FILLCELL_X2 FILLER_15_116 ();
 FILLCELL_X4 FILLER_15_121 ();
 FILLCELL_X1 FILLER_15_125 ();
 FILLCELL_X32 FILLER_15_136 ();
 FILLCELL_X4 FILLER_15_168 ();
 FILLCELL_X2 FILLER_15_172 ();
 FILLCELL_X4 FILLER_15_177 ();
 FILLCELL_X2 FILLER_15_181 ();
 FILLCELL_X1 FILLER_15_183 ();
 FILLCELL_X4 FILLER_15_187 ();
 FILLCELL_X1 FILLER_15_191 ();
 FILLCELL_X8 FILLER_15_195 ();
 FILLCELL_X4 FILLER_15_203 ();
 FILLCELL_X2 FILLER_15_207 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_40 ();
 FILLCELL_X8 FILLER_16_56 ();
 FILLCELL_X4 FILLER_16_64 ();
 FILLCELL_X2 FILLER_16_68 ();
 FILLCELL_X1 FILLER_16_70 ();
 FILLCELL_X32 FILLER_16_93 ();
 FILLCELL_X4 FILLER_16_125 ();
 FILLCELL_X32 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_174 ();
 FILLCELL_X1 FILLER_16_178 ();
 FILLCELL_X1 FILLER_16_182 ();
 FILLCELL_X16 FILLER_16_186 ();
 FILLCELL_X4 FILLER_16_202 ();
 FILLCELL_X2 FILLER_16_206 ();
 FILLCELL_X1 FILLER_16_208 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X16 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_81 ();
 FILLCELL_X4 FILLER_17_89 ();
 FILLCELL_X2 FILLER_17_93 ();
 FILLCELL_X1 FILLER_17_95 ();
 FILLCELL_X2 FILLER_17_100 ();
 FILLCELL_X8 FILLER_17_109 ();
 FILLCELL_X1 FILLER_17_117 ();
 FILLCELL_X2 FILLER_17_129 ();
 FILLCELL_X1 FILLER_17_134 ();
 FILLCELL_X32 FILLER_17_143 ();
 FILLCELL_X8 FILLER_17_175 ();
 FILLCELL_X4 FILLER_17_183 ();
 FILLCELL_X1 FILLER_17_187 ();
 FILLCELL_X16 FILLER_17_191 ();
 FILLCELL_X2 FILLER_17_207 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X16 FILLER_18_97 ();
 FILLCELL_X4 FILLER_18_113 ();
 FILLCELL_X2 FILLER_18_117 ();
 FILLCELL_X1 FILLER_18_119 ();
 FILLCELL_X4 FILLER_18_124 ();
 FILLCELL_X2 FILLER_18_128 ();
 FILLCELL_X32 FILLER_18_139 ();
 FILLCELL_X32 FILLER_18_171 ();
 FILLCELL_X4 FILLER_18_203 ();
 FILLCELL_X2 FILLER_18_207 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X16 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_81 ();
 FILLCELL_X4 FILLER_19_89 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X2 FILLER_19_113 ();
 FILLCELL_X1 FILLER_19_115 ();
 FILLCELL_X4 FILLER_19_125 ();
 FILLCELL_X2 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_139 ();
 FILLCELL_X32 FILLER_19_171 ();
 FILLCELL_X4 FILLER_19_203 ();
 FILLCELL_X2 FILLER_19_207 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X16 FILLER_20_65 ();
 FILLCELL_X8 FILLER_20_81 ();
 FILLCELL_X2 FILLER_20_89 ();
 FILLCELL_X1 FILLER_20_91 ();
 FILLCELL_X4 FILLER_20_108 ();
 FILLCELL_X2 FILLER_20_112 ();
 FILLCELL_X1 FILLER_20_114 ();
 FILLCELL_X16 FILLER_20_117 ();
 FILLCELL_X2 FILLER_20_133 ();
 FILLCELL_X32 FILLER_20_139 ();
 FILLCELL_X32 FILLER_20_171 ();
 FILLCELL_X4 FILLER_20_203 ();
 FILLCELL_X2 FILLER_20_207 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X2 FILLER_21_97 ();
 FILLCELL_X1 FILLER_21_99 ();
 FILLCELL_X8 FILLER_21_102 ();
 FILLCELL_X2 FILLER_21_110 ();
 FILLCELL_X2 FILLER_21_116 ();
 FILLCELL_X2 FILLER_21_122 ();
 FILLCELL_X1 FILLER_21_124 ();
 FILLCELL_X32 FILLER_21_137 ();
 FILLCELL_X32 FILLER_21_169 ();
 FILLCELL_X8 FILLER_21_201 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X16 FILLER_22_97 ();
 FILLCELL_X2 FILLER_22_113 ();
 FILLCELL_X1 FILLER_22_117 ();
 FILLCELL_X32 FILLER_22_127 ();
 FILLCELL_X32 FILLER_22_159 ();
 FILLCELL_X16 FILLER_22_191 ();
 FILLCELL_X2 FILLER_22_207 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X16 FILLER_23_193 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X16 FILLER_24_193 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X16 FILLER_25_193 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X16 FILLER_26_65 ();
 FILLCELL_X8 FILLER_26_81 ();
 FILLCELL_X4 FILLER_26_89 ();
 FILLCELL_X1 FILLER_26_93 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X4 FILLER_26_129 ();
 FILLCELL_X2 FILLER_26_133 ();
 FILLCELL_X1 FILLER_26_135 ();
 FILLCELL_X32 FILLER_26_140 ();
 FILLCELL_X32 FILLER_26_172 ();
 FILLCELL_X4 FILLER_26_204 ();
 FILLCELL_X1 FILLER_26_208 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X4 FILLER_27_81 ();
 FILLCELL_X2 FILLER_27_85 ();
 FILLCELL_X1 FILLER_27_87 ();
 FILLCELL_X1 FILLER_27_91 ();
 FILLCELL_X2 FILLER_27_95 ();
 FILLCELL_X2 FILLER_27_100 ();
 FILLCELL_X4 FILLER_27_105 ();
 FILLCELL_X1 FILLER_27_115 ();
 FILLCELL_X4 FILLER_27_119 ();
 FILLCELL_X2 FILLER_27_123 ();
 FILLCELL_X1 FILLER_27_125 ();
 FILLCELL_X2 FILLER_27_129 ();
 FILLCELL_X1 FILLER_27_131 ();
 FILLCELL_X1 FILLER_27_138 ();
 FILLCELL_X32 FILLER_27_142 ();
 FILLCELL_X32 FILLER_27_174 ();
 FILLCELL_X2 FILLER_27_206 ();
 FILLCELL_X1 FILLER_27_208 ();
endmodule
