module mesh_router (clk,
    east_in_ready,
    east_in_valid,
    east_out_ready,
    east_out_valid,
    local_in_ready,
    local_in_valid,
    local_out_ready,
    local_out_valid,
    north_in_ready,
    north_in_valid,
    north_out_ready,
    north_out_valid,
    rst_n,
    south_in_ready,
    south_in_valid,
    south_out_ready,
    south_out_valid,
    west_in_ready,
    west_in_valid,
    west_out_ready,
    west_out_valid,
    east_in_data,
    east_out_data,
    local_in_data,
    local_out_data,
    north_in_data,
    north_out_data,
    south_in_data,
    south_out_data,
    west_in_data,
    west_out_data);
 input clk;
 output east_in_ready;
 input east_in_valid;
 input east_out_ready;
 output east_out_valid;
 output local_in_ready;
 input local_in_valid;
 input local_out_ready;
 output local_out_valid;
 output north_in_ready;
 input north_in_valid;
 input north_out_ready;
 output north_out_valid;
 input rst_n;
 output south_in_ready;
 input south_in_valid;
 input south_out_ready;
 output south_out_valid;
 output west_in_ready;
 input west_in_valid;
 input west_out_ready;
 output west_out_valid;
 input [31:0] east_in_data;
 output [31:0] east_out_data;
 input [31:0] local_in_data;
 output [31:0] local_out_data;
 input [31:0] north_in_data;
 output [31:0] north_out_data;
 input [31:0] south_in_data;
 output [31:0] south_out_data;
 input [31:0] west_in_data;
 output [31:0] west_out_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire net343;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire \dest_id[0][0] ;
 wire \dest_id[0][1] ;
 wire \dest_id[0][2] ;
 wire \dest_id[0][3] ;
 wire \dest_id[0][4] ;
 wire \dest_id[0][5] ;
 wire \dest_id[0][6] ;
 wire \dest_id[0][7] ;
 wire \dest_id[1][0] ;
 wire \dest_id[1][1] ;
 wire \dest_id[1][2] ;
 wire \dest_id[1][3] ;
 wire \dest_id[1][4] ;
 wire \dest_id[1][5] ;
 wire \dest_id[1][6] ;
 wire \dest_id[1][7] ;
 wire \dest_id[2][0] ;
 wire \dest_id[2][1] ;
 wire \dest_id[2][2] ;
 wire \dest_id[2][3] ;
 wire \dest_id[2][4] ;
 wire \dest_id[2][5] ;
 wire \dest_id[2][6] ;
 wire \dest_id[2][7] ;
 wire \dest_id[3][0] ;
 wire \dest_id[3][1] ;
 wire \dest_id[3][2] ;
 wire \dest_id[3][3] ;
 wire \dest_id[3][4] ;
 wire \dest_id[3][5] ;
 wire \dest_id[3][6] ;
 wire \dest_id[3][7] ;
 wire \dest_id[4][0] ;
 wire \dest_id[4][1] ;
 wire \dest_id[4][2] ;
 wire \dest_id[4][3] ;
 wire \dest_id[4][4] ;
 wire \dest_id[4][5] ;
 wire \dest_id[4][6] ;
 wire \dest_id[4][7] ;
 wire \input_buffer[0][0] ;
 wire \input_buffer[0][10] ;
 wire \input_buffer[0][11] ;
 wire \input_buffer[0][12] ;
 wire \input_buffer[0][13] ;
 wire \input_buffer[0][14] ;
 wire \input_buffer[0][15] ;
 wire \input_buffer[0][16] ;
 wire \input_buffer[0][17] ;
 wire \input_buffer[0][18] ;
 wire \input_buffer[0][19] ;
 wire \input_buffer[0][1] ;
 wire \input_buffer[0][20] ;
 wire \input_buffer[0][21] ;
 wire \input_buffer[0][22] ;
 wire \input_buffer[0][23] ;
 wire \input_buffer[0][2] ;
 wire \input_buffer[0][3] ;
 wire \input_buffer[0][4] ;
 wire \input_buffer[0][5] ;
 wire \input_buffer[0][6] ;
 wire \input_buffer[0][7] ;
 wire \input_buffer[0][8] ;
 wire \input_buffer[0][9] ;
 wire \input_buffer[1][0] ;
 wire \input_buffer[1][10] ;
 wire \input_buffer[1][11] ;
 wire \input_buffer[1][12] ;
 wire \input_buffer[1][13] ;
 wire \input_buffer[1][14] ;
 wire \input_buffer[1][15] ;
 wire \input_buffer[1][16] ;
 wire \input_buffer[1][17] ;
 wire \input_buffer[1][18] ;
 wire \input_buffer[1][19] ;
 wire \input_buffer[1][1] ;
 wire \input_buffer[1][20] ;
 wire \input_buffer[1][21] ;
 wire \input_buffer[1][22] ;
 wire \input_buffer[1][23] ;
 wire \input_buffer[1][2] ;
 wire \input_buffer[1][3] ;
 wire \input_buffer[1][4] ;
 wire \input_buffer[1][5] ;
 wire \input_buffer[1][6] ;
 wire \input_buffer[1][7] ;
 wire \input_buffer[1][8] ;
 wire \input_buffer[1][9] ;
 wire \input_buffer[2][0] ;
 wire \input_buffer[2][10] ;
 wire \input_buffer[2][11] ;
 wire \input_buffer[2][12] ;
 wire \input_buffer[2][13] ;
 wire \input_buffer[2][14] ;
 wire \input_buffer[2][15] ;
 wire \input_buffer[2][16] ;
 wire \input_buffer[2][17] ;
 wire \input_buffer[2][18] ;
 wire \input_buffer[2][19] ;
 wire \input_buffer[2][1] ;
 wire \input_buffer[2][20] ;
 wire \input_buffer[2][21] ;
 wire \input_buffer[2][22] ;
 wire \input_buffer[2][23] ;
 wire \input_buffer[2][2] ;
 wire \input_buffer[2][3] ;
 wire \input_buffer[2][4] ;
 wire \input_buffer[2][5] ;
 wire \input_buffer[2][6] ;
 wire \input_buffer[2][7] ;
 wire \input_buffer[2][8] ;
 wire \input_buffer[2][9] ;
 wire \input_buffer[3][0] ;
 wire \input_buffer[3][10] ;
 wire \input_buffer[3][11] ;
 wire \input_buffer[3][12] ;
 wire \input_buffer[3][13] ;
 wire \input_buffer[3][14] ;
 wire \input_buffer[3][15] ;
 wire \input_buffer[3][16] ;
 wire \input_buffer[3][17] ;
 wire \input_buffer[3][18] ;
 wire \input_buffer[3][19] ;
 wire \input_buffer[3][1] ;
 wire \input_buffer[3][20] ;
 wire \input_buffer[3][21] ;
 wire \input_buffer[3][22] ;
 wire \input_buffer[3][23] ;
 wire \input_buffer[3][2] ;
 wire \input_buffer[3][3] ;
 wire \input_buffer[3][4] ;
 wire \input_buffer[3][5] ;
 wire \input_buffer[3][6] ;
 wire \input_buffer[3][7] ;
 wire \input_buffer[3][8] ;
 wire \input_buffer[3][9] ;
 wire \input_buffer[4][0] ;
 wire \input_buffer[4][10] ;
 wire \input_buffer[4][11] ;
 wire \input_buffer[4][12] ;
 wire \input_buffer[4][13] ;
 wire \input_buffer[4][14] ;
 wire \input_buffer[4][15] ;
 wire \input_buffer[4][16] ;
 wire \input_buffer[4][17] ;
 wire \input_buffer[4][18] ;
 wire \input_buffer[4][19] ;
 wire \input_buffer[4][1] ;
 wire \input_buffer[4][20] ;
 wire \input_buffer[4][21] ;
 wire \input_buffer[4][22] ;
 wire \input_buffer[4][23] ;
 wire \input_buffer[4][2] ;
 wire \input_buffer[4][3] ;
 wire \input_buffer[4][4] ;
 wire \input_buffer[4][5] ;
 wire \input_buffer[4][6] ;
 wire \input_buffer[4][7] ;
 wire \input_buffer[4][8] ;
 wire \input_buffer[4][9] ;
 wire \input_buffer_valid[0] ;
 wire \input_buffer_valid[1] ;
 wire \input_buffer_valid[2] ;
 wire \input_buffer_valid[3] ;
 wire \input_buffer_valid[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net344;

 OR4_X2 _1606_ (.A1(\dest_id[4][5] ),
    .A2(\dest_id[4][4] ),
    .A3(\dest_id[4][7] ),
    .A4(\dest_id[4][6] ),
    .ZN(_1274_));
 BUF_X8 _1607_ (.A(_1274_),
    .Z(_1275_));
 INV_X1 _1608_ (.A(_1275_),
    .ZN(_1276_));
 BUF_X4 _1609_ (.A(\dest_id[4][0] ),
    .Z(_1277_));
 INV_X2 _1610_ (.A(_1277_),
    .ZN(_1278_));
 CLKBUF_X3 _1611_ (.A(\dest_id[4][1] ),
    .Z(_1279_));
 CLKBUF_X3 _1612_ (.A(\dest_id[4][2] ),
    .Z(_1280_));
 NOR3_X4 _1613_ (.A1(_1278_),
    .A2(_1279_),
    .A3(_1280_),
    .ZN(_1281_));
 BUF_X4 _1614_ (.A(\dest_id[4][3] ),
    .Z(_1282_));
 INV_X2 _1615_ (.A(_1280_),
    .ZN(_1283_));
 NOR3_X4 _1616_ (.A1(_1277_),
    .A2(_1282_),
    .A3(_1283_),
    .ZN(_1284_));
 OAI21_X4 _1617_ (.A(_1276_),
    .B1(_1281_),
    .B2(_1284_),
    .ZN(_1285_));
 INV_X4 _1618_ (.A(_1285_),
    .ZN(_1603_));
 NOR4_X4 _1619_ (.A1(_1275_),
    .A2(_1282_),
    .A3(_1283_),
    .A4(_1277_),
    .ZN(_1592_));
 INV_X1 _1620_ (.A(_1592_),
    .ZN(_1595_));
 NOR2_X1 _1621_ (.A1(_1279_),
    .A2(_1275_),
    .ZN(_1286_));
 INV_X2 _1622_ (.A(_1282_),
    .ZN(_1287_));
 NOR3_X1 _1623_ (.A1(_1278_),
    .A2(_1287_),
    .A3(_1280_),
    .ZN(_1288_));
 OAI21_X2 _1624_ (.A(_1286_),
    .B1(_1288_),
    .B2(_1284_),
    .ZN(_1591_));
 INV_X1 _1625_ (.A(_1591_),
    .ZN(_1598_));
 BUF_X2 _1626_ (.A(\dest_id[3][5] ),
    .Z(_1289_));
 BUF_X2 _1627_ (.A(\dest_id[3][4] ),
    .Z(_1290_));
 BUF_X2 _1628_ (.A(\dest_id[3][7] ),
    .Z(_1291_));
 BUF_X2 _1629_ (.A(\dest_id[3][6] ),
    .Z(_1292_));
 NOR4_X4 _1630_ (.A1(_1289_),
    .A2(_1290_),
    .A3(_1291_),
    .A4(_1292_),
    .ZN(_1293_));
 INV_X1 _1631_ (.A(\dest_id[3][0] ),
    .ZN(_1294_));
 BUF_X4 _1632_ (.A(\dest_id[3][2] ),
    .Z(_1295_));
 NOR3_X4 _1633_ (.A1(_1294_),
    .A2(\dest_id[3][1] ),
    .A3(_1295_),
    .ZN(_1296_));
 INV_X2 _1634_ (.A(_1295_),
    .ZN(_1297_));
 NOR3_X4 _1635_ (.A1(\dest_id[3][0] ),
    .A2(\dest_id[3][3] ),
    .A3(_1297_),
    .ZN(_1298_));
 OAI21_X4 _1636_ (.A(_1293_),
    .B1(_1296_),
    .B2(_1298_),
    .ZN(_1299_));
 INV_X2 _1637_ (.A(_1299_),
    .ZN(_1588_));
 CLKBUF_X3 _1638_ (.A(\dest_id[3][0] ),
    .Z(_1300_));
 NOR2_X1 _1639_ (.A1(_1300_),
    .A2(_1297_),
    .ZN(_1301_));
 BUF_X4 _1640_ (.A(\dest_id[3][3] ),
    .Z(_1302_));
 OR4_X4 _1641_ (.A1(_1289_),
    .A2(_1290_),
    .A3(_1291_),
    .A4(_1292_),
    .ZN(_1303_));
 NOR2_X2 _1642_ (.A1(_1302_),
    .A2(_1303_),
    .ZN(_1304_));
 NAND2_X2 _1643_ (.A1(_1301_),
    .A2(_1304_),
    .ZN(_1580_));
 CLKBUF_X3 _1644_ (.A(\dest_id[3][1] ),
    .Z(_1305_));
 OR2_X1 _1645_ (.A1(_1305_),
    .A2(_1303_),
    .ZN(_1306_));
 NAND3_X1 _1646_ (.A1(_1300_),
    .A2(_1302_),
    .A3(_1297_),
    .ZN(_1307_));
 OR3_X2 _1647_ (.A1(_1300_),
    .A2(\dest_id[3][3] ),
    .A3(_1297_),
    .ZN(_1308_));
 AOI21_X2 _1648_ (.A(_1306_),
    .B1(_1307_),
    .B2(_1308_),
    .ZN(_1583_));
 BUF_X2 _1649_ (.A(\dest_id[2][5] ),
    .Z(_1309_));
 BUF_X2 _1650_ (.A(\dest_id[2][4] ),
    .Z(_1310_));
 BUF_X2 _1651_ (.A(\dest_id[2][7] ),
    .Z(_1311_));
 BUF_X2 _1652_ (.A(\dest_id[2][6] ),
    .Z(_1312_));
 NOR4_X4 _1653_ (.A1(_1309_),
    .A2(_1310_),
    .A3(_1311_),
    .A4(_1312_),
    .ZN(_1313_));
 BUF_X4 _1654_ (.A(\dest_id[2][0] ),
    .Z(_1314_));
 INV_X2 _1655_ (.A(_1314_),
    .ZN(_1315_));
 BUF_X4 _1656_ (.A(\dest_id[2][1] ),
    .Z(_1316_));
 BUF_X4 _1657_ (.A(\dest_id[2][2] ),
    .Z(_1317_));
 NOR3_X4 _1658_ (.A1(_1315_),
    .A2(_1316_),
    .A3(_1317_),
    .ZN(_1318_));
 BUF_X4 _1659_ (.A(\dest_id[2][3] ),
    .Z(_1319_));
 INV_X2 _1660_ (.A(_1317_),
    .ZN(_1320_));
 NOR3_X4 _1661_ (.A1(_1314_),
    .A2(_1319_),
    .A3(_1320_),
    .ZN(_1321_));
 OAI21_X4 _1662_ (.A(_1313_),
    .B1(_1318_),
    .B2(_1321_),
    .ZN(_1322_));
 INV_X2 _1663_ (.A(_1322_),
    .ZN(_1573_));
 OR4_X4 _1664_ (.A1(_1309_),
    .A2(_1310_),
    .A3(_1311_),
    .A4(_1312_),
    .ZN(_1323_));
 NOR4_X4 _1665_ (.A1(_1323_),
    .A2(_1319_),
    .A3(_1320_),
    .A4(_1314_),
    .ZN(_1562_));
 INV_X1 _1666_ (.A(_1562_),
    .ZN(_1565_));
 OR2_X2 _1667_ (.A1(_1316_),
    .A2(_1323_),
    .ZN(_1324_));
 NAND3_X2 _1668_ (.A1(_1314_),
    .A2(_1319_),
    .A3(_1320_),
    .ZN(_1325_));
 INV_X2 _1669_ (.A(_1319_),
    .ZN(_1326_));
 NAND3_X4 _1670_ (.A1(_1315_),
    .A2(_1326_),
    .A3(_1317_),
    .ZN(_1327_));
 AOI21_X4 _1671_ (.A(_1324_),
    .B1(_1325_),
    .B2(_1327_),
    .ZN(_1568_));
 BUF_X2 _1672_ (.A(\dest_id[1][5] ),
    .Z(_1328_));
 BUF_X2 _1673_ (.A(\dest_id[1][4] ),
    .Z(_1329_));
 BUF_X2 _1674_ (.A(\dest_id[1][7] ),
    .Z(_1330_));
 BUF_X2 _1675_ (.A(\dest_id[1][6] ),
    .Z(_1331_));
 NOR4_X4 _1676_ (.A1(_1328_),
    .A2(_1329_),
    .A3(_1330_),
    .A4(_1331_),
    .ZN(_1332_));
 BUF_X4 _1677_ (.A(\dest_id[1][0] ),
    .Z(_1333_));
 INV_X2 _1678_ (.A(_1333_),
    .ZN(_1334_));
 CLKBUF_X3 _1679_ (.A(\dest_id[1][1] ),
    .Z(_1335_));
 BUF_X4 _1680_ (.A(\dest_id[1][2] ),
    .Z(_1336_));
 NOR3_X4 _1681_ (.A1(_1334_),
    .A2(_1335_),
    .A3(_1336_),
    .ZN(_1337_));
 CLKBUF_X3 _1682_ (.A(\dest_id[1][3] ),
    .Z(_1338_));
 INV_X2 _1683_ (.A(_1336_),
    .ZN(_1339_));
 NOR3_X4 _1684_ (.A1(_1339_),
    .A2(_1338_),
    .A3(_1333_),
    .ZN(_1340_));
 OAI21_X4 _1685_ (.A(_1332_),
    .B1(_1337_),
    .B2(_1340_),
    .ZN(_1341_));
 INV_X4 _1686_ (.A(_1341_),
    .ZN(_1342_));
 BUF_X4 _1687_ (.A(_1342_),
    .Z(_1558_));
 NOR2_X1 _1688_ (.A1(_1333_),
    .A2(_1339_),
    .ZN(_1343_));
 OR4_X4 _1689_ (.A1(_1328_),
    .A2(_1329_),
    .A3(_1330_),
    .A4(_1331_),
    .ZN(_1344_));
 NOR2_X4 _1690_ (.A1(_1338_),
    .A2(_1344_),
    .ZN(_1345_));
 AND2_X4 _1691_ (.A1(_1343_),
    .A2(_1345_),
    .ZN(_1547_));
 INV_X1 _1692_ (.A(_1547_),
    .ZN(_1550_));
 NOR2_X1 _1693_ (.A1(_1335_),
    .A2(_1344_),
    .ZN(_1346_));
 INV_X2 _1694_ (.A(_1338_),
    .ZN(_1347_));
 NOR3_X2 _1695_ (.A1(_1334_),
    .A2(_1347_),
    .A3(_1336_),
    .ZN(_1348_));
 OAI21_X2 _1696_ (.A(_1346_),
    .B1(_1348_),
    .B2(_1340_),
    .ZN(_1546_));
 INV_X1 _1697_ (.A(_1546_),
    .ZN(_1553_));
 BUF_X2 _1698_ (.A(\dest_id[0][3] ),
    .Z(_1349_));
 INV_X1 _1699_ (.A(\dest_id[0][2] ),
    .ZN(_1350_));
 NOR3_X4 _1700_ (.A1(\dest_id[0][0] ),
    .A2(_1349_),
    .A3(_1350_),
    .ZN(_1351_));
 INV_X1 _1701_ (.A(\dest_id[0][0] ),
    .ZN(_1352_));
 INV_X1 _1702_ (.A(_1349_),
    .ZN(_1353_));
 NOR3_X2 _1703_ (.A1(_1352_),
    .A2(_1353_),
    .A3(\dest_id[0][2] ),
    .ZN(_1354_));
 NOR2_X1 _1704_ (.A1(_1351_),
    .A2(_1354_),
    .ZN(_1355_));
 OR4_X1 _1705_ (.A1(\dest_id[0][5] ),
    .A2(\dest_id[0][4] ),
    .A3(\dest_id[0][7] ),
    .A4(\dest_id[0][6] ),
    .ZN(_1356_));
 OR3_X2 _1706_ (.A1(\dest_id[0][1] ),
    .A2(_1355_),
    .A3(_1356_),
    .ZN(_1532_));
 INV_X1 _1707_ (.A(_1532_),
    .ZN(_1535_));
 NOR2_X1 _1708_ (.A1(\dest_id[0][0] ),
    .A2(_1350_),
    .ZN(_1357_));
 NOR2_X1 _1709_ (.A1(_1349_),
    .A2(_1356_),
    .ZN(_1358_));
 AND2_X1 _1710_ (.A1(_1357_),
    .A2(_1358_),
    .ZN(_1531_));
 INV_X1 _1711_ (.A(_1531_),
    .ZN(_1538_));
 INV_X1 _1712_ (.A(_1568_),
    .ZN(_1561_));
 INV_X1 _1713_ (.A(_1583_),
    .ZN(_1576_));
 NOR4_X4 _1714_ (.A1(\dest_id[0][5] ),
    .A2(\dest_id[0][4] ),
    .A3(\dest_id[0][7] ),
    .A4(\dest_id[0][6] ),
    .ZN(_1359_));
 NOR3_X4 _1715_ (.A1(_1352_),
    .A2(\dest_id[0][1] ),
    .A3(\dest_id[0][2] ),
    .ZN(_1360_));
 OAI21_X4 _1716_ (.A(_1359_),
    .B1(_1360_),
    .B2(_1351_),
    .ZN(_1361_));
 INV_X2 _1717_ (.A(_1361_),
    .ZN(_1362_));
 BUF_X4 _1718_ (.A(_1362_),
    .Z(_1543_));
 INV_X1 _1719_ (.A(_1580_),
    .ZN(_1577_));
 BUF_X4 _1720_ (.A(rst_n),
    .Z(_1363_));
 CLKBUF_X3 _1721_ (.A(\input_buffer_valid[0] ),
    .Z(_1364_));
 INV_X4 _1722_ (.A(_1364_),
    .ZN(_1365_));
 BUF_X4 _1723_ (.A(_1365_),
    .Z(_1366_));
 BUF_X8 _1724_ (.A(_1366_),
    .Z(_1367_));
 NAND3_X2 _1725_ (.A1(_1363_),
    .A2(_1367_),
    .A3(net100),
    .ZN(_1368_));
 CLKBUF_X3 _1726_ (.A(_1368_),
    .Z(_1369_));
 MUX2_X1 _1727_ (.A(net68),
    .B(\input_buffer[0][0] ),
    .S(_1369_),
    .Z(_0032_));
 MUX2_X1 _1728_ (.A(net69),
    .B(\input_buffer[0][10] ),
    .S(_1369_),
    .Z(_0033_));
 MUX2_X1 _1729_ (.A(net70),
    .B(\input_buffer[0][11] ),
    .S(_1369_),
    .Z(_0034_));
 MUX2_X1 _1730_ (.A(net71),
    .B(\input_buffer[0][12] ),
    .S(_1369_),
    .Z(_0035_));
 MUX2_X1 _1731_ (.A(net72),
    .B(\input_buffer[0][13] ),
    .S(_1369_),
    .Z(_0036_));
 MUX2_X1 _1732_ (.A(net73),
    .B(\input_buffer[0][14] ),
    .S(_1369_),
    .Z(_0037_));
 MUX2_X1 _1733_ (.A(net74),
    .B(\input_buffer[0][15] ),
    .S(_1369_),
    .Z(_0038_));
 MUX2_X1 _1734_ (.A(net75),
    .B(\input_buffer[0][16] ),
    .S(_1369_),
    .Z(_0039_));
 MUX2_X1 _1735_ (.A(net76),
    .B(\input_buffer[0][17] ),
    .S(_1369_),
    .Z(_0040_));
 MUX2_X1 _1736_ (.A(net77),
    .B(\input_buffer[0][18] ),
    .S(_1369_),
    .Z(_0041_));
 CLKBUF_X3 _1737_ (.A(_1368_),
    .Z(_1370_));
 MUX2_X1 _1738_ (.A(net78),
    .B(\input_buffer[0][19] ),
    .S(_1370_),
    .Z(_0042_));
 MUX2_X1 _1739_ (.A(net79),
    .B(\input_buffer[0][1] ),
    .S(_1370_),
    .Z(_0043_));
 MUX2_X1 _1740_ (.A(net80),
    .B(\input_buffer[0][20] ),
    .S(_1370_),
    .Z(_0044_));
 MUX2_X1 _1741_ (.A(net81),
    .B(\input_buffer[0][21] ),
    .S(_1370_),
    .Z(_0045_));
 MUX2_X1 _1742_ (.A(net82),
    .B(\input_buffer[0][22] ),
    .S(_1370_),
    .Z(_0046_));
 MUX2_X1 _1743_ (.A(net83),
    .B(\input_buffer[0][23] ),
    .S(_1370_),
    .Z(_0047_));
 MUX2_X1 _1744_ (.A(net84),
    .B(\dest_id[0][0] ),
    .S(_1370_),
    .Z(_0048_));
 MUX2_X1 _1745_ (.A(net85),
    .B(\dest_id[0][1] ),
    .S(_1370_),
    .Z(_0049_));
 MUX2_X1 _1746_ (.A(net86),
    .B(\dest_id[0][2] ),
    .S(_1370_),
    .Z(_0050_));
 MUX2_X1 _1747_ (.A(net87),
    .B(_1349_),
    .S(_1370_),
    .Z(_0051_));
 CLKBUF_X3 _1748_ (.A(_1368_),
    .Z(_1371_));
 MUX2_X1 _1749_ (.A(net88),
    .B(\dest_id[0][4] ),
    .S(_1371_),
    .Z(_0052_));
 MUX2_X1 _1750_ (.A(net89),
    .B(\dest_id[0][5] ),
    .S(_1371_),
    .Z(_0053_));
 MUX2_X1 _1751_ (.A(net90),
    .B(\input_buffer[0][2] ),
    .S(_1371_),
    .Z(_0054_));
 MUX2_X1 _1752_ (.A(net91),
    .B(\dest_id[0][6] ),
    .S(_1371_),
    .Z(_0055_));
 MUX2_X1 _1753_ (.A(net92),
    .B(\dest_id[0][7] ),
    .S(_1371_),
    .Z(_0056_));
 MUX2_X1 _1754_ (.A(net93),
    .B(\input_buffer[0][3] ),
    .S(_1371_),
    .Z(_0057_));
 MUX2_X1 _1755_ (.A(net94),
    .B(\input_buffer[0][4] ),
    .S(_1371_),
    .Z(_0058_));
 MUX2_X1 _1756_ (.A(net95),
    .B(\input_buffer[0][5] ),
    .S(_1371_),
    .Z(_0059_));
 MUX2_X1 _1757_ (.A(net96),
    .B(\input_buffer[0][6] ),
    .S(_1371_),
    .Z(_0060_));
 MUX2_X1 _1758_ (.A(net97),
    .B(\input_buffer[0][7] ),
    .S(_1371_),
    .Z(_0061_));
 MUX2_X1 _1759_ (.A(net98),
    .B(\input_buffer[0][8] ),
    .S(_1368_),
    .Z(_0062_));
 MUX2_X1 _1760_ (.A(net99),
    .B(\input_buffer[0][9] ),
    .S(_1368_),
    .Z(_0063_));
 CLKBUF_X3 _1761_ (.A(\input_buffer_valid[1] ),
    .Z(_1372_));
 CLKBUF_X3 _1762_ (.A(_1372_),
    .Z(_1373_));
 INV_X2 _1763_ (.A(_1373_),
    .ZN(_1374_));
 NAND3_X2 _1764_ (.A1(_1363_),
    .A2(_1374_),
    .A3(net33),
    .ZN(_1375_));
 CLKBUF_X3 _1765_ (.A(_1375_),
    .Z(_1376_));
 MUX2_X1 _1766_ (.A(net1),
    .B(\input_buffer[1][0] ),
    .S(_1376_),
    .Z(_0064_));
 MUX2_X1 _1767_ (.A(net2),
    .B(\input_buffer[1][10] ),
    .S(_1376_),
    .Z(_0065_));
 MUX2_X1 _1768_ (.A(net3),
    .B(\input_buffer[1][11] ),
    .S(_1376_),
    .Z(_0066_));
 MUX2_X1 _1769_ (.A(net4),
    .B(\input_buffer[1][12] ),
    .S(_1376_),
    .Z(_0067_));
 MUX2_X1 _1770_ (.A(net5),
    .B(\input_buffer[1][13] ),
    .S(_1376_),
    .Z(_0068_));
 MUX2_X1 _1771_ (.A(net6),
    .B(\input_buffer[1][14] ),
    .S(_1376_),
    .Z(_0069_));
 MUX2_X1 _1772_ (.A(net7),
    .B(\input_buffer[1][15] ),
    .S(_1376_),
    .Z(_0070_));
 MUX2_X1 _1773_ (.A(net8),
    .B(\input_buffer[1][16] ),
    .S(_1376_),
    .Z(_0071_));
 MUX2_X1 _1774_ (.A(net9),
    .B(\input_buffer[1][17] ),
    .S(_1376_),
    .Z(_0072_));
 MUX2_X1 _1775_ (.A(net10),
    .B(\input_buffer[1][18] ),
    .S(_1376_),
    .Z(_0073_));
 CLKBUF_X3 _1776_ (.A(_1375_),
    .Z(_1377_));
 MUX2_X1 _1777_ (.A(net11),
    .B(\input_buffer[1][19] ),
    .S(_1377_),
    .Z(_0074_));
 MUX2_X1 _1778_ (.A(net12),
    .B(\input_buffer[1][1] ),
    .S(_1377_),
    .Z(_0075_));
 MUX2_X1 _1779_ (.A(net13),
    .B(\input_buffer[1][20] ),
    .S(_1377_),
    .Z(_0076_));
 MUX2_X1 _1780_ (.A(net14),
    .B(\input_buffer[1][21] ),
    .S(_1377_),
    .Z(_0077_));
 MUX2_X1 _1781_ (.A(net15),
    .B(\input_buffer[1][22] ),
    .S(_1377_),
    .Z(_0078_));
 MUX2_X1 _1782_ (.A(net16),
    .B(\input_buffer[1][23] ),
    .S(_1377_),
    .Z(_0079_));
 MUX2_X1 _1783_ (.A(net17),
    .B(_1333_),
    .S(_1377_),
    .Z(_0080_));
 MUX2_X1 _1784_ (.A(net18),
    .B(_1335_),
    .S(_1377_),
    .Z(_0081_));
 MUX2_X1 _1785_ (.A(net19),
    .B(_1336_),
    .S(_1377_),
    .Z(_0082_));
 MUX2_X1 _1786_ (.A(net20),
    .B(_1338_),
    .S(_1377_),
    .Z(_0083_));
 CLKBUF_X3 _1787_ (.A(_1375_),
    .Z(_1378_));
 MUX2_X1 _1788_ (.A(net21),
    .B(_1329_),
    .S(_1378_),
    .Z(_0084_));
 MUX2_X1 _1789_ (.A(net22),
    .B(_1328_),
    .S(_1378_),
    .Z(_0085_));
 MUX2_X1 _1790_ (.A(net23),
    .B(\input_buffer[1][2] ),
    .S(_1378_),
    .Z(_0086_));
 MUX2_X1 _1791_ (.A(net24),
    .B(_1331_),
    .S(_1378_),
    .Z(_0087_));
 MUX2_X1 _1792_ (.A(net25),
    .B(_1330_),
    .S(_1378_),
    .Z(_0088_));
 MUX2_X1 _1793_ (.A(net26),
    .B(\input_buffer[1][3] ),
    .S(_1378_),
    .Z(_0089_));
 MUX2_X1 _1794_ (.A(net27),
    .B(\input_buffer[1][4] ),
    .S(_1378_),
    .Z(_0090_));
 MUX2_X1 _1795_ (.A(net28),
    .B(\input_buffer[1][5] ),
    .S(_1378_),
    .Z(_0091_));
 MUX2_X1 _1796_ (.A(net29),
    .B(\input_buffer[1][6] ),
    .S(_1378_),
    .Z(_0092_));
 MUX2_X1 _1797_ (.A(net30),
    .B(\input_buffer[1][7] ),
    .S(_1378_),
    .Z(_0093_));
 MUX2_X1 _1798_ (.A(net31),
    .B(\input_buffer[1][8] ),
    .S(_1375_),
    .Z(_0094_));
 MUX2_X1 _1799_ (.A(net32),
    .B(\input_buffer[1][9] ),
    .S(_1375_),
    .Z(_0095_));
 BUF_X2 _1800_ (.A(\input_buffer[2][0] ),
    .Z(_1379_));
 BUF_X4 _1801_ (.A(\input_buffer_valid[2] ),
    .Z(_1380_));
 INV_X4 _1802_ (.A(_1380_),
    .ZN(_1381_));
 AND2_X1 _1803_ (.A1(_1381_),
    .A2(net133),
    .ZN(_1382_));
 NAND2_X4 _1804_ (.A1(_1363_),
    .A2(_1382_),
    .ZN(_1383_));
 BUF_X4 _1805_ (.A(_1383_),
    .Z(_1384_));
 MUX2_X1 _1806_ (.A(net101),
    .B(_1379_),
    .S(_1384_),
    .Z(_0096_));
 CLKBUF_X2 _1807_ (.A(\input_buffer[2][10] ),
    .Z(_1385_));
 MUX2_X1 _1808_ (.A(net102),
    .B(_1385_),
    .S(_1384_),
    .Z(_0097_));
 CLKBUF_X2 _1809_ (.A(\input_buffer[2][11] ),
    .Z(_1386_));
 MUX2_X1 _1810_ (.A(net103),
    .B(_1386_),
    .S(_1384_),
    .Z(_0098_));
 CLKBUF_X2 _1811_ (.A(\input_buffer[2][12] ),
    .Z(_1387_));
 MUX2_X1 _1812_ (.A(net104),
    .B(_1387_),
    .S(_1384_),
    .Z(_0099_));
 CLKBUF_X2 _1813_ (.A(\input_buffer[2][13] ),
    .Z(_1388_));
 MUX2_X1 _1814_ (.A(net105),
    .B(_1388_),
    .S(_1384_),
    .Z(_0100_));
 CLKBUF_X2 _1815_ (.A(\input_buffer[2][14] ),
    .Z(_1389_));
 MUX2_X1 _1816_ (.A(net106),
    .B(_1389_),
    .S(_1384_),
    .Z(_0101_));
 BUF_X2 _1817_ (.A(\input_buffer[2][15] ),
    .Z(_1390_));
 MUX2_X1 _1818_ (.A(net107),
    .B(_1390_),
    .S(_1384_),
    .Z(_0102_));
 CLKBUF_X2 _1819_ (.A(\input_buffer[2][16] ),
    .Z(_1391_));
 MUX2_X1 _1820_ (.A(net108),
    .B(_1391_),
    .S(_1384_),
    .Z(_0103_));
 CLKBUF_X2 _1821_ (.A(\input_buffer[2][17] ),
    .Z(_1392_));
 MUX2_X1 _1822_ (.A(net109),
    .B(_1392_),
    .S(_1384_),
    .Z(_0104_));
 CLKBUF_X2 _1823_ (.A(\input_buffer[2][18] ),
    .Z(_1393_));
 MUX2_X1 _1824_ (.A(net110),
    .B(_1393_),
    .S(_1384_),
    .Z(_0105_));
 BUF_X2 _1825_ (.A(\input_buffer[2][19] ),
    .Z(_1394_));
 CLKBUF_X3 _1826_ (.A(_1383_),
    .Z(_1395_));
 MUX2_X1 _1827_ (.A(net111),
    .B(_1394_),
    .S(_1395_),
    .Z(_0106_));
 CLKBUF_X2 _1828_ (.A(\input_buffer[2][1] ),
    .Z(_1396_));
 MUX2_X1 _1829_ (.A(net112),
    .B(_1396_),
    .S(_1395_),
    .Z(_0107_));
 BUF_X2 _1830_ (.A(\input_buffer[2][20] ),
    .Z(_1397_));
 MUX2_X1 _1831_ (.A(net113),
    .B(_1397_),
    .S(_1395_),
    .Z(_0108_));
 CLKBUF_X2 _1832_ (.A(\input_buffer[2][21] ),
    .Z(_1398_));
 MUX2_X1 _1833_ (.A(net114),
    .B(_1398_),
    .S(_1395_),
    .Z(_0109_));
 CLKBUF_X2 _1834_ (.A(\input_buffer[2][22] ),
    .Z(_1399_));
 MUX2_X1 _1835_ (.A(net115),
    .B(_1399_),
    .S(_1395_),
    .Z(_0110_));
 BUF_X2 _1836_ (.A(\input_buffer[2][23] ),
    .Z(_1400_));
 MUX2_X1 _1837_ (.A(net116),
    .B(_1400_),
    .S(_1395_),
    .Z(_0111_));
 MUX2_X1 _1838_ (.A(net117),
    .B(_1314_),
    .S(_1395_),
    .Z(_0112_));
 MUX2_X1 _1839_ (.A(net118),
    .B(_1316_),
    .S(_1395_),
    .Z(_0113_));
 MUX2_X1 _1840_ (.A(net119),
    .B(_1317_),
    .S(_1395_),
    .Z(_0114_));
 MUX2_X1 _1841_ (.A(net120),
    .B(_1319_),
    .S(_1395_),
    .Z(_0115_));
 CLKBUF_X3 _1842_ (.A(_1383_),
    .Z(_1401_));
 MUX2_X1 _1843_ (.A(net121),
    .B(_1310_),
    .S(_1401_),
    .Z(_0116_));
 MUX2_X1 _1844_ (.A(net122),
    .B(_1309_),
    .S(_1401_),
    .Z(_0117_));
 BUF_X2 _1845_ (.A(\input_buffer[2][2] ),
    .Z(_1402_));
 MUX2_X1 _1846_ (.A(net123),
    .B(_1402_),
    .S(_1401_),
    .Z(_0118_));
 MUX2_X1 _1847_ (.A(net124),
    .B(_1312_),
    .S(_1401_),
    .Z(_0119_));
 MUX2_X1 _1848_ (.A(net125),
    .B(_1311_),
    .S(_1401_),
    .Z(_0120_));
 BUF_X2 _1849_ (.A(\input_buffer[2][3] ),
    .Z(_0197_));
 MUX2_X1 _1850_ (.A(net126),
    .B(_0197_),
    .S(_1401_),
    .Z(_0121_));
 CLKBUF_X2 _1851_ (.A(\input_buffer[2][4] ),
    .Z(_0198_));
 MUX2_X1 _1852_ (.A(net127),
    .B(_0198_),
    .S(_1401_),
    .Z(_0122_));
 CLKBUF_X2 _1853_ (.A(\input_buffer[2][5] ),
    .Z(_0199_));
 MUX2_X1 _1854_ (.A(net128),
    .B(_0199_),
    .S(_1401_),
    .Z(_0123_));
 CLKBUF_X2 _1855_ (.A(\input_buffer[2][6] ),
    .Z(_0200_));
 MUX2_X1 _1856_ (.A(net129),
    .B(_0200_),
    .S(_1401_),
    .Z(_0124_));
 CLKBUF_X2 _1857_ (.A(\input_buffer[2][7] ),
    .Z(_0201_));
 MUX2_X1 _1858_ (.A(net130),
    .B(_0201_),
    .S(_1401_),
    .Z(_0125_));
 CLKBUF_X2 _1859_ (.A(\input_buffer[2][8] ),
    .Z(_0202_));
 MUX2_X1 _1860_ (.A(net131),
    .B(_0202_),
    .S(_1383_),
    .Z(_0126_));
 BUF_X2 _1861_ (.A(\input_buffer[2][9] ),
    .Z(_0203_));
 MUX2_X1 _1862_ (.A(net132),
    .B(_0203_),
    .S(_1383_),
    .Z(_0127_));
 BUF_X2 _1863_ (.A(\input_buffer[3][0] ),
    .Z(_0204_));
 BUF_X4 _1864_ (.A(\input_buffer_valid[3] ),
    .Z(_0205_));
 INV_X4 _1865_ (.A(_0205_),
    .ZN(_0206_));
 NAND3_X4 _1866_ (.A1(_1363_),
    .A2(_0206_),
    .A3(net167),
    .ZN(_0207_));
 BUF_X4 _1867_ (.A(_0207_),
    .Z(_0208_));
 MUX2_X1 _1868_ (.A(net135),
    .B(_0204_),
    .S(_0208_),
    .Z(_0128_));
 BUF_X2 _1869_ (.A(\input_buffer[3][10] ),
    .Z(_0209_));
 MUX2_X1 _1870_ (.A(net136),
    .B(_0209_),
    .S(_0208_),
    .Z(_0129_));
 BUF_X2 _1871_ (.A(\input_buffer[3][11] ),
    .Z(_0210_));
 MUX2_X1 _1872_ (.A(net137),
    .B(_0210_),
    .S(_0208_),
    .Z(_0130_));
 BUF_X2 _1873_ (.A(\input_buffer[3][12] ),
    .Z(_0211_));
 MUX2_X1 _1874_ (.A(net138),
    .B(_0211_),
    .S(_0208_),
    .Z(_0131_));
 BUF_X2 _1875_ (.A(\input_buffer[3][13] ),
    .Z(_0212_));
 MUX2_X1 _1876_ (.A(net139),
    .B(_0212_),
    .S(_0208_),
    .Z(_0132_));
 BUF_X2 _1877_ (.A(\input_buffer[3][14] ),
    .Z(_0213_));
 MUX2_X1 _1878_ (.A(net140),
    .B(_0213_),
    .S(_0208_),
    .Z(_0133_));
 BUF_X2 _1879_ (.A(\input_buffer[3][15] ),
    .Z(_0214_));
 MUX2_X1 _1880_ (.A(net141),
    .B(_0214_),
    .S(_0208_),
    .Z(_0134_));
 BUF_X2 _1881_ (.A(\input_buffer[3][16] ),
    .Z(_0215_));
 MUX2_X1 _1882_ (.A(net142),
    .B(_0215_),
    .S(_0208_),
    .Z(_0135_));
 BUF_X2 _1883_ (.A(\input_buffer[3][17] ),
    .Z(_0216_));
 MUX2_X1 _1884_ (.A(net143),
    .B(_0216_),
    .S(_0208_),
    .Z(_0136_));
 BUF_X2 _1885_ (.A(\input_buffer[3][18] ),
    .Z(_0217_));
 MUX2_X1 _1886_ (.A(net144),
    .B(_0217_),
    .S(_0208_),
    .Z(_0137_));
 BUF_X2 _1887_ (.A(\input_buffer[3][19] ),
    .Z(_0218_));
 CLKBUF_X3 _1888_ (.A(_0207_),
    .Z(_0219_));
 MUX2_X1 _1889_ (.A(net145),
    .B(_0218_),
    .S(_0219_),
    .Z(_0138_));
 BUF_X2 _1890_ (.A(\input_buffer[3][1] ),
    .Z(_0220_));
 MUX2_X1 _1891_ (.A(net146),
    .B(_0220_),
    .S(_0219_),
    .Z(_0139_));
 BUF_X2 _1892_ (.A(\input_buffer[3][20] ),
    .Z(_0221_));
 MUX2_X1 _1893_ (.A(net147),
    .B(_0221_),
    .S(_0219_),
    .Z(_0140_));
 BUF_X2 _1894_ (.A(\input_buffer[3][21] ),
    .Z(_0222_));
 MUX2_X1 _1895_ (.A(net148),
    .B(_0222_),
    .S(_0219_),
    .Z(_0141_));
 BUF_X2 _1896_ (.A(\input_buffer[3][22] ),
    .Z(_0223_));
 MUX2_X1 _1897_ (.A(net149),
    .B(_0223_),
    .S(_0219_),
    .Z(_0142_));
 BUF_X2 _1898_ (.A(\input_buffer[3][23] ),
    .Z(_0224_));
 MUX2_X1 _1899_ (.A(net150),
    .B(_0224_),
    .S(_0219_),
    .Z(_0143_));
 MUX2_X1 _1900_ (.A(net151),
    .B(_1300_),
    .S(_0219_),
    .Z(_0144_));
 MUX2_X1 _1901_ (.A(net152),
    .B(_1305_),
    .S(_0219_),
    .Z(_0145_));
 MUX2_X1 _1902_ (.A(net153),
    .B(_1295_),
    .S(_0219_),
    .Z(_0146_));
 MUX2_X1 _1903_ (.A(net154),
    .B(_1302_),
    .S(_0219_),
    .Z(_0147_));
 CLKBUF_X3 _1904_ (.A(_0207_),
    .Z(_0225_));
 MUX2_X1 _1905_ (.A(net155),
    .B(_1290_),
    .S(_0225_),
    .Z(_0148_));
 MUX2_X1 _1906_ (.A(net156),
    .B(_1289_),
    .S(_0225_),
    .Z(_0149_));
 BUF_X2 _1907_ (.A(\input_buffer[3][2] ),
    .Z(_0226_));
 MUX2_X1 _1908_ (.A(net157),
    .B(_0226_),
    .S(_0225_),
    .Z(_0150_));
 MUX2_X1 _1909_ (.A(net158),
    .B(_1292_),
    .S(_0225_),
    .Z(_0151_));
 MUX2_X1 _1910_ (.A(net159),
    .B(_1291_),
    .S(_0225_),
    .Z(_0152_));
 BUF_X2 _1911_ (.A(\input_buffer[3][3] ),
    .Z(_0227_));
 MUX2_X1 _1912_ (.A(net160),
    .B(_0227_),
    .S(_0225_),
    .Z(_0153_));
 BUF_X2 _1913_ (.A(\input_buffer[3][4] ),
    .Z(_0228_));
 MUX2_X1 _1914_ (.A(net161),
    .B(_0228_),
    .S(_0225_),
    .Z(_0154_));
 BUF_X2 _1915_ (.A(\input_buffer[3][5] ),
    .Z(_0229_));
 MUX2_X1 _1916_ (.A(net162),
    .B(_0229_),
    .S(_0225_),
    .Z(_0155_));
 BUF_X2 _1917_ (.A(\input_buffer[3][6] ),
    .Z(_0230_));
 MUX2_X1 _1918_ (.A(net163),
    .B(_0230_),
    .S(_0225_),
    .Z(_0156_));
 BUF_X2 _1919_ (.A(\input_buffer[3][7] ),
    .Z(_0231_));
 MUX2_X1 _1920_ (.A(net164),
    .B(_0231_),
    .S(_0225_),
    .Z(_0157_));
 BUF_X2 _1921_ (.A(\input_buffer[3][8] ),
    .Z(_0232_));
 MUX2_X1 _1922_ (.A(net165),
    .B(_0232_),
    .S(_0207_),
    .Z(_0158_));
 CLKBUF_X2 _1923_ (.A(\input_buffer[3][9] ),
    .Z(_0233_));
 MUX2_X1 _1924_ (.A(net166),
    .B(_0233_),
    .S(_0207_),
    .Z(_0159_));
 BUF_X2 _1925_ (.A(\input_buffer[4][0] ),
    .Z(_0234_));
 BUF_X2 _1926_ (.A(\input_buffer_valid[4] ),
    .Z(_0235_));
 INV_X2 _1927_ (.A(_0235_),
    .ZN(_0236_));
 NAND3_X4 _1928_ (.A1(_0236_),
    .A2(net67),
    .A3(_1363_),
    .ZN(_0237_));
 CLKBUF_X3 _1929_ (.A(_0237_),
    .Z(_0238_));
 MUX2_X1 _1930_ (.A(net35),
    .B(_0234_),
    .S(_0238_),
    .Z(_0160_));
 BUF_X2 _1931_ (.A(\input_buffer[4][10] ),
    .Z(_0239_));
 MUX2_X1 _1932_ (.A(net36),
    .B(_0239_),
    .S(_0238_),
    .Z(_0161_));
 BUF_X2 _1933_ (.A(\input_buffer[4][11] ),
    .Z(_0240_));
 MUX2_X1 _1934_ (.A(net37),
    .B(_0240_),
    .S(_0238_),
    .Z(_0162_));
 BUF_X2 _1935_ (.A(\input_buffer[4][12] ),
    .Z(_0241_));
 MUX2_X1 _1936_ (.A(net38),
    .B(_0241_),
    .S(_0238_),
    .Z(_0163_));
 BUF_X2 _1937_ (.A(\input_buffer[4][13] ),
    .Z(_0242_));
 MUX2_X1 _1938_ (.A(net39),
    .B(_0242_),
    .S(_0238_),
    .Z(_0164_));
 BUF_X2 _1939_ (.A(\input_buffer[4][14] ),
    .Z(_0243_));
 MUX2_X1 _1940_ (.A(net40),
    .B(_0243_),
    .S(_0238_),
    .Z(_0165_));
 BUF_X2 _1941_ (.A(\input_buffer[4][15] ),
    .Z(_0244_));
 MUX2_X1 _1942_ (.A(net41),
    .B(_0244_),
    .S(_0238_),
    .Z(_0166_));
 BUF_X2 _1943_ (.A(\input_buffer[4][16] ),
    .Z(_0245_));
 MUX2_X1 _1944_ (.A(net42),
    .B(_0245_),
    .S(_0238_),
    .Z(_0167_));
 CLKBUF_X2 _1945_ (.A(\input_buffer[4][17] ),
    .Z(_0246_));
 MUX2_X1 _1946_ (.A(net43),
    .B(_0246_),
    .S(_0238_),
    .Z(_0168_));
 CLKBUF_X2 _1947_ (.A(\input_buffer[4][18] ),
    .Z(_0247_));
 MUX2_X1 _1948_ (.A(net44),
    .B(_0247_),
    .S(_0238_),
    .Z(_0169_));
 CLKBUF_X2 _1949_ (.A(\input_buffer[4][19] ),
    .Z(_0248_));
 CLKBUF_X3 _1950_ (.A(_0237_),
    .Z(_0249_));
 MUX2_X1 _1951_ (.A(net45),
    .B(_0248_),
    .S(_0249_),
    .Z(_0170_));
 CLKBUF_X2 _1952_ (.A(\input_buffer[4][1] ),
    .Z(_0250_));
 MUX2_X1 _1953_ (.A(net46),
    .B(_0250_),
    .S(_0249_),
    .Z(_0171_));
 BUF_X2 _1954_ (.A(\input_buffer[4][20] ),
    .Z(_0251_));
 MUX2_X1 _1955_ (.A(net47),
    .B(_0251_),
    .S(_0249_),
    .Z(_0172_));
 CLKBUF_X2 _1956_ (.A(\input_buffer[4][21] ),
    .Z(_0252_));
 MUX2_X1 _1957_ (.A(net48),
    .B(_0252_),
    .S(_0249_),
    .Z(_0173_));
 CLKBUF_X2 _1958_ (.A(\input_buffer[4][22] ),
    .Z(_0253_));
 MUX2_X1 _1959_ (.A(net49),
    .B(_0253_),
    .S(_0249_),
    .Z(_0174_));
 CLKBUF_X2 _1960_ (.A(\input_buffer[4][23] ),
    .Z(_0254_));
 MUX2_X1 _1961_ (.A(net50),
    .B(_0254_),
    .S(_0249_),
    .Z(_0175_));
 MUX2_X1 _1962_ (.A(net51),
    .B(_1277_),
    .S(_0249_),
    .Z(_0176_));
 MUX2_X1 _1963_ (.A(net52),
    .B(_1279_),
    .S(_0249_),
    .Z(_0177_));
 MUX2_X1 _1964_ (.A(net53),
    .B(_1280_),
    .S(_0249_),
    .Z(_0178_));
 MUX2_X1 _1965_ (.A(net54),
    .B(_1282_),
    .S(_0249_),
    .Z(_0179_));
 CLKBUF_X3 _1966_ (.A(_0237_),
    .Z(_0255_));
 MUX2_X1 _1967_ (.A(net55),
    .B(\dest_id[4][4] ),
    .S(_0255_),
    .Z(_0180_));
 MUX2_X1 _1968_ (.A(net56),
    .B(\dest_id[4][5] ),
    .S(_0255_),
    .Z(_0181_));
 BUF_X2 _1969_ (.A(\input_buffer[4][2] ),
    .Z(_0256_));
 MUX2_X1 _1970_ (.A(net57),
    .B(_0256_),
    .S(_0255_),
    .Z(_0182_));
 MUX2_X1 _1971_ (.A(net58),
    .B(\dest_id[4][6] ),
    .S(_0255_),
    .Z(_0183_));
 MUX2_X1 _1972_ (.A(net59),
    .B(\dest_id[4][7] ),
    .S(_0255_),
    .Z(_0184_));
 BUF_X2 _1973_ (.A(\input_buffer[4][3] ),
    .Z(_0257_));
 MUX2_X1 _1974_ (.A(net60),
    .B(_0257_),
    .S(_0255_),
    .Z(_0185_));
 BUF_X2 _1975_ (.A(\input_buffer[4][4] ),
    .Z(_0258_));
 MUX2_X1 _1976_ (.A(net61),
    .B(_0258_),
    .S(_0255_),
    .Z(_0186_));
 BUF_X2 _1977_ (.A(\input_buffer[4][5] ),
    .Z(_0259_));
 MUX2_X1 _1978_ (.A(net62),
    .B(_0259_),
    .S(_0255_),
    .Z(_0187_));
 BUF_X2 _1979_ (.A(\input_buffer[4][6] ),
    .Z(_0260_));
 MUX2_X1 _1980_ (.A(net63),
    .B(_0260_),
    .S(_0255_),
    .Z(_0188_));
 BUF_X2 _1981_ (.A(\input_buffer[4][7] ),
    .Z(_0261_));
 MUX2_X1 _1982_ (.A(net64),
    .B(_0261_),
    .S(_0255_),
    .Z(_0189_));
 CLKBUF_X2 _1983_ (.A(\input_buffer[4][8] ),
    .Z(_0262_));
 MUX2_X1 _1984_ (.A(net65),
    .B(_0262_),
    .S(_0237_),
    .Z(_0190_));
 BUF_X2 _1985_ (.A(\input_buffer[4][9] ),
    .Z(_0263_));
 MUX2_X1 _1986_ (.A(net66),
    .B(_0263_),
    .S(_0237_),
    .Z(_0191_));
 CLKBUF_X3 _1987_ (.A(_1364_),
    .Z(_0264_));
 OAI21_X1 _1988_ (.A(_1363_),
    .B1(_0264_),
    .B2(net100),
    .ZN(_0265_));
 CLKBUF_X2 _1989_ (.A(local_out_ready),
    .Z(_0266_));
 NOR2_X1 _1990_ (.A1(_0266_),
    .A2(_1543_),
    .ZN(_0267_));
 BUF_X2 _1991_ (.A(_1536_),
    .Z(_0268_));
 CLKBUF_X3 _1992_ (.A(_1544_),
    .Z(_0269_));
 BUF_X4 _1993_ (.A(_0269_),
    .Z(_0270_));
 NOR4_X2 _1994_ (.A1(_1533_),
    .A2(_0268_),
    .A3(_1541_),
    .A4(_0270_),
    .ZN(_0271_));
 CLKBUF_X2 _1995_ (.A(north_out_ready),
    .Z(_0272_));
 INV_X1 _1996_ (.A(_0272_),
    .ZN(_0273_));
 INV_X1 _1997_ (.A(net34),
    .ZN(_0274_));
 AND2_X1 _1998_ (.A1(_0274_),
    .A2(\dest_id[0][1] ),
    .ZN(_0275_));
 AOI22_X2 _1999_ (.A1(_0273_),
    .A2(_1360_),
    .B1(_0275_),
    .B2(_1357_),
    .ZN(_0276_));
 INV_X1 _2000_ (.A(net168),
    .ZN(_0277_));
 INV_X1 _2001_ (.A(net134),
    .ZN(_0278_));
 AOI22_X2 _2002_ (.A1(_0277_),
    .A2(_1351_),
    .B1(_1354_),
    .B2(_0278_),
    .ZN(_0279_));
 OAI22_X2 _2003_ (.A1(_1349_),
    .A2(_0276_),
    .B1(_0279_),
    .B2(\dest_id[0][1] ),
    .ZN(_0280_));
 AOI221_X2 _2004_ (.A(_0267_),
    .B1(_0271_),
    .B2(_1543_),
    .C1(_1359_),
    .C2(_0280_),
    .ZN(_0281_));
 NOR2_X1 _2005_ (.A1(_1367_),
    .A2(net237),
    .ZN(_0282_));
 AOI21_X1 _2006_ (.A(_0265_),
    .B1(_0281_),
    .B2(_0282_),
    .ZN(_0192_));
 CLKBUF_X3 _2007_ (.A(_1373_),
    .Z(_0283_));
 BUF_X4 _2008_ (.A(_0283_),
    .Z(_0284_));
 OAI21_X1 _2009_ (.A(_1363_),
    .B1(_0284_),
    .B2(net33),
    .ZN(_0285_));
 NOR2_X1 _2010_ (.A1(_0266_),
    .A2(_1558_),
    .ZN(_0286_));
 CLKBUF_X3 _2011_ (.A(_1554_),
    .Z(_0287_));
 BUF_X2 _2012_ (.A(_1556_),
    .Z(_0288_));
 NOR4_X1 _2013_ (.A1(_1559_),
    .A2(_1548_),
    .A3(_0287_),
    .A4(_0288_),
    .ZN(_0289_));
 AND2_X1 _2014_ (.A1(_1558_),
    .A2(_0289_),
    .ZN(_0290_));
 NOR4_X1 _2015_ (.A1(_1374_),
    .A2(net169),
    .A3(_0286_),
    .A4(_0290_),
    .ZN(_0291_));
 NAND3_X1 _2016_ (.A1(_0274_),
    .A2(_1335_),
    .A3(_1343_),
    .ZN(_0292_));
 OR3_X4 _2017_ (.A1(_1334_),
    .A2(_1335_),
    .A3(_1336_),
    .ZN(_0293_));
 OAI21_X1 _2018_ (.A(_0292_),
    .B1(_0293_),
    .B2(_0272_),
    .ZN(_0294_));
 NAND2_X1 _2019_ (.A1(_0278_),
    .A2(_1348_),
    .ZN(_0295_));
 NAND3_X4 _2020_ (.A1(_1334_),
    .A2(_1347_),
    .A3(_1336_),
    .ZN(_0296_));
 OAI21_X1 _2021_ (.A(_0295_),
    .B1(_0296_),
    .B2(net168),
    .ZN(_0297_));
 AOI22_X1 _2022_ (.A1(_1345_),
    .A2(_0294_),
    .B1(_0297_),
    .B2(_1346_),
    .ZN(_0298_));
 AOI21_X1 _2023_ (.A(_0285_),
    .B1(_0291_),
    .B2(_0298_),
    .ZN(_0193_));
 INV_X1 _2024_ (.A(_1363_),
    .ZN(_0299_));
 AOI21_X1 _2025_ (.A(_1381_),
    .B1(_0266_),
    .B2(_1322_),
    .ZN(_0300_));
 MUX2_X1 _2026_ (.A(net134),
    .B(net168),
    .S(_1562_),
    .Z(_0301_));
 BUF_X2 _2027_ (.A(_1563_),
    .Z(_0302_));
 BUF_X2 _2028_ (.A(_1569_),
    .Z(_0303_));
 BUF_X2 _2029_ (.A(_1571_),
    .Z(_0304_));
 OR4_X1 _2030_ (.A1(_1574_),
    .A2(_0302_),
    .A3(_0303_),
    .A4(_0304_),
    .ZN(_0305_));
 NAND3_X1 _2031_ (.A1(_1568_),
    .A2(_0301_),
    .A3(_0305_),
    .ZN(_0306_));
 MUX2_X1 _2032_ (.A(_0272_),
    .B(net34),
    .S(_1321_),
    .Z(_0307_));
 OR3_X4 _2033_ (.A1(_1315_),
    .A2(_1316_),
    .A3(_1317_),
    .ZN(_0308_));
 NAND3_X1 _2034_ (.A1(_1315_),
    .A2(_1316_),
    .A3(_1317_),
    .ZN(_0309_));
 AOI21_X2 _2035_ (.A(_1319_),
    .B1(_0308_),
    .B2(_0309_),
    .ZN(_0310_));
 NAND4_X1 _2036_ (.A1(_1313_),
    .A2(_0305_),
    .A3(_0307_),
    .A4(_0310_),
    .ZN(_0311_));
 NAND3_X1 _2037_ (.A1(_0300_),
    .A2(_0306_),
    .A3(_0311_),
    .ZN(_0312_));
 AOI21_X1 _2038_ (.A(_1382_),
    .B1(net271),
    .B2(_1380_),
    .ZN(_0313_));
 AOI21_X1 _2039_ (.A(_0299_),
    .B1(_0312_),
    .B2(_0313_),
    .ZN(_0194_));
 CLKBUF_X3 _2040_ (.A(_0205_),
    .Z(_0314_));
 OAI21_X1 _2041_ (.A(_1363_),
    .B1(_0314_),
    .B2(net167),
    .ZN(_0315_));
 OR2_X1 _2042_ (.A1(_0206_),
    .A2(net305),
    .ZN(_0316_));
 NAND2_X1 _2043_ (.A1(net134),
    .A2(_1580_),
    .ZN(_0317_));
 NAND2_X1 _2044_ (.A1(_0277_),
    .A2(_1298_),
    .ZN(_0318_));
 AOI21_X1 _2045_ (.A(_1306_),
    .B1(_1307_),
    .B2(_0318_),
    .ZN(_0319_));
 NAND3_X1 _2046_ (.A1(_0274_),
    .A2(_1305_),
    .A3(_1301_),
    .ZN(_0320_));
 OR3_X2 _2047_ (.A1(_1294_),
    .A2(_1305_),
    .A3(_1295_),
    .ZN(_0321_));
 OAI21_X1 _2048_ (.A(_0320_),
    .B1(_0321_),
    .B2(_0272_),
    .ZN(_0322_));
 AOI221_X2 _2049_ (.A(_0316_),
    .B1(_0317_),
    .B2(_0319_),
    .C1(_0322_),
    .C2(_1304_),
    .ZN(_0323_));
 NAND2_X1 _2050_ (.A1(_0266_),
    .A2(_1299_),
    .ZN(_0324_));
 CLKBUF_X3 _2051_ (.A(_1589_),
    .Z(_0325_));
 BUF_X4 _2052_ (.A(_0325_),
    .Z(_0326_));
 BUF_X2 _2053_ (.A(_1584_),
    .Z(_0327_));
 NOR4_X1 _2054_ (.A1(_0326_),
    .A2(_1578_),
    .A3(_0327_),
    .A4(_1586_),
    .ZN(_0328_));
 OAI21_X1 _2055_ (.A(_0324_),
    .B1(_0328_),
    .B2(_1299_),
    .ZN(_0329_));
 AOI21_X1 _2056_ (.A(_0315_),
    .B1(_0323_),
    .B2(_0329_),
    .ZN(_0195_));
 BUF_X4 _2057_ (.A(_0235_),
    .Z(_0330_));
 MUX2_X1 _2058_ (.A(_0272_),
    .B(net34),
    .S(_1592_),
    .Z(_0331_));
 NOR2_X1 _2059_ (.A1(_1282_),
    .A2(_1275_),
    .ZN(_0332_));
 AND3_X1 _2060_ (.A1(_1278_),
    .A2(_1279_),
    .A3(_1280_),
    .ZN(_0333_));
 OAI21_X2 _2061_ (.A(_0332_),
    .B1(_0333_),
    .B2(_1281_),
    .ZN(_0334_));
 OAI221_X1 _2062_ (.A(_0330_),
    .B1(_0266_),
    .B2(_1603_),
    .C1(_0331_),
    .C2(_0334_),
    .ZN(_0335_));
 MUX2_X1 _2063_ (.A(net134),
    .B(net168),
    .S(_1592_),
    .Z(_0336_));
 NOR2_X1 _2064_ (.A1(_1591_),
    .A2(_0336_),
    .ZN(_0337_));
 OAI221_X1 _2065_ (.A(_1363_),
    .B1(_0335_),
    .B2(_0337_),
    .C1(net67),
    .C2(_0330_),
    .ZN(_0338_));
 INV_X1 _2066_ (.A(_0338_),
    .ZN(_0196_));
 NAND2_X1 _2067_ (.A1(_0235_),
    .A2(_1593_),
    .ZN(_0339_));
 NAND3_X1 _2068_ (.A1(_1278_),
    .A2(_1287_),
    .A3(_1280_),
    .ZN(_0340_));
 OR3_X1 _2069_ (.A1(_1278_),
    .A2(_1279_),
    .A3(_1280_),
    .ZN(_0341_));
 AOI211_X4 _2070_ (.A(_1275_),
    .B(_0339_),
    .C1(_0340_),
    .C2(_0341_),
    .ZN(_0342_));
 CLKBUF_X3 _2071_ (.A(_0342_),
    .Z(_0343_));
 BUF_X4 _2072_ (.A(_0343_),
    .Z(_0344_));
 INV_X2 _2073_ (.A(_1578_),
    .ZN(_0345_));
 NOR2_X4 _2074_ (.A1(_0206_),
    .A2(_1303_),
    .ZN(_0346_));
 OAI21_X2 _2075_ (.A(_0346_),
    .B1(_1298_),
    .B2(_1296_),
    .ZN(_0347_));
 NOR3_X4 _2076_ (.A1(_0345_),
    .A2(_0347_),
    .A3(_0342_),
    .ZN(_0348_));
 BUF_X4 _2077_ (.A(_0348_),
    .Z(_0349_));
 AOI22_X1 _2078_ (.A1(_0234_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0204_),
    .ZN(_0350_));
 OR2_X1 _2079_ (.A1(_1285_),
    .A2(_0339_),
    .ZN(_0351_));
 NAND2_X2 _2080_ (.A1(_0308_),
    .A2(_1327_),
    .ZN(_0352_));
 NAND4_X4 _2081_ (.A1(_1380_),
    .A2(_0302_),
    .A3(_1313_),
    .A4(_0352_),
    .ZN(_0353_));
 OAI221_X2 _2082_ (.A(_0351_),
    .B1(_0347_),
    .B2(_0345_),
    .C1(_1379_),
    .C2(_0353_),
    .ZN(_0354_));
 NAND3_X1 _2083_ (.A1(_1380_),
    .A2(_0302_),
    .A3(_1313_),
    .ZN(_0355_));
 AOI21_X4 _2084_ (.A(_0355_),
    .B1(_1327_),
    .B2(_0308_),
    .ZN(_0356_));
 INV_X2 _2085_ (.A(_1533_),
    .ZN(_0357_));
 NAND3_X2 _2086_ (.A1(_1372_),
    .A2(_1548_),
    .A3(net339),
    .ZN(_0358_));
 AOI21_X4 _2087_ (.A(_0358_),
    .B1(_0296_),
    .B2(_0293_),
    .ZN(_0359_));
 NOR2_X4 _2088_ (.A1(_0357_),
    .A2(_0359_),
    .ZN(_0360_));
 BUF_X4 _2089_ (.A(_0360_),
    .Z(_0361_));
 NOR2_X1 _2090_ (.A1(_1366_),
    .A2(_0005_),
    .ZN(_0362_));
 AND2_X1 _2091_ (.A1(_1543_),
    .A2(_0362_),
    .ZN(_0363_));
 INV_X2 _2092_ (.A(_1548_),
    .ZN(_0364_));
 NAND2_X1 _2093_ (.A1(_0283_),
    .A2(\input_buffer[1][0] ),
    .ZN(_0365_));
 NOR2_X1 _2094_ (.A1(_0364_),
    .A2(_0365_),
    .ZN(_0366_));
 AOI221_X1 _2095_ (.A(_0356_),
    .B1(_0361_),
    .B2(_0363_),
    .C1(_0366_),
    .C2(_1558_),
    .ZN(_0367_));
 OAI21_X1 _2096_ (.A(_0350_),
    .B1(_0354_),
    .B2(_0367_),
    .ZN(net170));
 AOI22_X1 _2097_ (.A1(_0239_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0209_),
    .ZN(_0368_));
 NAND2_X2 _2098_ (.A1(_0205_),
    .A2(_1293_),
    .ZN(_0369_));
 AOI211_X2 _2099_ (.A(_0345_),
    .B(_0369_),
    .C1(_1308_),
    .C2(_0321_),
    .ZN(_0370_));
 NOR2_X4 _2100_ (.A1(_0370_),
    .A2(_0342_),
    .ZN(_0371_));
 CLKBUF_X3 _2101_ (.A(_0371_),
    .Z(_0372_));
 CLKBUF_X3 _2102_ (.A(_0353_),
    .Z(_0373_));
 OAI21_X1 _2103_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1385_),
    .ZN(_0374_));
 INV_X1 _2104_ (.A(_0302_),
    .ZN(_0375_));
 NOR2_X4 _2105_ (.A1(_1381_),
    .A2(_1323_),
    .ZN(_0376_));
 OAI21_X4 _2106_ (.A(_0376_),
    .B1(_1321_),
    .B2(_1318_),
    .ZN(_0377_));
 NOR2_X4 _2107_ (.A1(_0375_),
    .A2(_0377_),
    .ZN(_0378_));
 BUF_X4 _2108_ (.A(_0378_),
    .Z(_0379_));
 CLKBUF_X3 _2109_ (.A(_1361_),
    .Z(_0380_));
 INV_X1 _2110_ (.A(_0015_),
    .ZN(_0381_));
 NAND2_X1 _2111_ (.A1(_1364_),
    .A2(_0381_),
    .ZN(_0382_));
 NOR2_X1 _2112_ (.A1(_0380_),
    .A2(_0382_),
    .ZN(_0383_));
 AND2_X1 _2113_ (.A1(_0283_),
    .A2(\input_buffer[1][10] ),
    .ZN(_0384_));
 NOR2_X4 _2114_ (.A1(_0364_),
    .A2(_1341_),
    .ZN(_0385_));
 BUF_X4 _2115_ (.A(_0385_),
    .Z(_0386_));
 AOI221_X1 _2116_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0383_),
    .C1(_0384_),
    .C2(_0386_),
    .ZN(_0387_));
 OAI21_X1 _2117_ (.A(_0368_),
    .B1(_0374_),
    .B2(_0387_),
    .ZN(net171));
 AOI22_X1 _2118_ (.A1(_0240_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0210_),
    .ZN(_0388_));
 OAI21_X1 _2119_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1386_),
    .ZN(_0389_));
 NOR2_X1 _2120_ (.A1(_1366_),
    .A2(_0016_),
    .ZN(_0390_));
 AND2_X1 _2121_ (.A1(_1543_),
    .A2(_0390_),
    .ZN(_0391_));
 NAND2_X1 _2122_ (.A1(_1373_),
    .A2(\input_buffer[1][11] ),
    .ZN(_0392_));
 NOR2_X1 _2123_ (.A1(_0364_),
    .A2(_0392_),
    .ZN(_0393_));
 AOI221_X2 _2124_ (.A(_0356_),
    .B1(_0361_),
    .B2(_0391_),
    .C1(_0393_),
    .C2(_1558_),
    .ZN(_0394_));
 OAI21_X1 _2125_ (.A(_0388_),
    .B1(_0389_),
    .B2(_0394_),
    .ZN(net172));
 AOI22_X1 _2126_ (.A1(_0241_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0211_),
    .ZN(_0395_));
 OAI21_X1 _2127_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1387_),
    .ZN(_0396_));
 BUF_X8 _2128_ (.A(_1361_),
    .Z(_0397_));
 NOR3_X4 _2129_ (.A1(_1367_),
    .A2(_0017_),
    .A3(_0397_),
    .ZN(_0398_));
 AND2_X2 _2130_ (.A1(_0283_),
    .A2(\input_buffer[1][12] ),
    .ZN(_0399_));
 AOI221_X2 _2131_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0398_),
    .C1(_0399_),
    .C2(_0386_),
    .ZN(_0400_));
 OAI21_X1 _2132_ (.A(_0395_),
    .B1(_0396_),
    .B2(_0400_),
    .ZN(net173));
 AOI22_X1 _2133_ (.A1(_0242_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0212_),
    .ZN(_0401_));
 OAI21_X1 _2134_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1388_),
    .ZN(_0402_));
 BUF_X8 _2135_ (.A(_1366_),
    .Z(_0403_));
 NOR3_X4 _2136_ (.A1(_0403_),
    .A2(_0018_),
    .A3(_0397_),
    .ZN(_0404_));
 AND2_X2 _2137_ (.A1(_0283_),
    .A2(\input_buffer[1][13] ),
    .ZN(_0405_));
 AOI221_X2 _2138_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0404_),
    .C1(_0405_),
    .C2(_0386_),
    .ZN(_0406_));
 OAI21_X1 _2139_ (.A(_0401_),
    .B1(_0402_),
    .B2(_0406_),
    .ZN(net174));
 AOI22_X1 _2140_ (.A1(_0243_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0213_),
    .ZN(_0407_));
 OAI21_X1 _2141_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1389_),
    .ZN(_0408_));
 NOR3_X4 _2142_ (.A1(_0403_),
    .A2(_0019_),
    .A3(_0397_),
    .ZN(_0409_));
 AND2_X2 _2143_ (.A1(_0283_),
    .A2(\input_buffer[1][14] ),
    .ZN(_0410_));
 AOI221_X2 _2144_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0409_),
    .C1(_0410_),
    .C2(_0386_),
    .ZN(_0411_));
 OAI21_X1 _2145_ (.A(_0407_),
    .B1(_0408_),
    .B2(_0411_),
    .ZN(net175));
 AOI22_X1 _2146_ (.A1(_0244_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0214_),
    .ZN(_0412_));
 OAI21_X1 _2147_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1390_),
    .ZN(_0413_));
 NOR3_X4 _2148_ (.A1(_0403_),
    .A2(_0020_),
    .A3(_0397_),
    .ZN(_0414_));
 AND2_X2 _2149_ (.A1(_0283_),
    .A2(\input_buffer[1][15] ),
    .ZN(_0415_));
 AOI221_X2 _2150_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0414_),
    .C1(_0415_),
    .C2(_0386_),
    .ZN(_0416_));
 OAI21_X1 _2151_ (.A(_0412_),
    .B1(_0413_),
    .B2(_0416_),
    .ZN(net176));
 AOI22_X1 _2152_ (.A1(_0245_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0215_),
    .ZN(_0417_));
 OAI21_X1 _2153_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1391_),
    .ZN(_0418_));
 BUF_X4 _2154_ (.A(_1361_),
    .Z(_0419_));
 NOR3_X4 _2155_ (.A1(_0403_),
    .A2(_0021_),
    .A3(_0419_),
    .ZN(_0420_));
 AND2_X2 _2156_ (.A1(_0283_),
    .A2(\input_buffer[1][16] ),
    .ZN(_0421_));
 AOI221_X2 _2157_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0420_),
    .C1(_0421_),
    .C2(_0386_),
    .ZN(_0422_));
 OAI21_X1 _2158_ (.A(_0417_),
    .B1(_0418_),
    .B2(_0422_),
    .ZN(net177));
 AOI22_X1 _2159_ (.A1(_0246_),
    .A2(_0344_),
    .B1(_0349_),
    .B2(_0216_),
    .ZN(_0423_));
 OAI21_X1 _2160_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1392_),
    .ZN(_0424_));
 NOR3_X2 _2161_ (.A1(_0403_),
    .A2(_0022_),
    .A3(_0419_),
    .ZN(_0425_));
 BUF_X2 _2162_ (.A(_1372_),
    .Z(_0426_));
 AND2_X1 _2163_ (.A1(_0426_),
    .A2(\input_buffer[1][17] ),
    .ZN(_0427_));
 AOI221_X1 _2164_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0425_),
    .C1(_0427_),
    .C2(_0386_),
    .ZN(_0428_));
 OAI21_X1 _2165_ (.A(_0423_),
    .B1(_0424_),
    .B2(_0428_),
    .ZN(net178));
 CLKBUF_X3 _2166_ (.A(_0342_),
    .Z(_0429_));
 AOI22_X1 _2167_ (.A1(_0247_),
    .A2(_0429_),
    .B1(_0349_),
    .B2(_0217_),
    .ZN(_0430_));
 OAI21_X1 _2168_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1393_),
    .ZN(_0431_));
 NOR3_X2 _2169_ (.A1(_0403_),
    .A2(_0023_),
    .A3(_0419_),
    .ZN(_0432_));
 AND2_X1 _2170_ (.A1(_0426_),
    .A2(\input_buffer[1][18] ),
    .ZN(_0433_));
 AOI221_X1 _2171_ (.A(_0379_),
    .B1(_0361_),
    .B2(_0432_),
    .C1(_0433_),
    .C2(_0386_),
    .ZN(_0434_));
 OAI21_X1 _2172_ (.A(_0430_),
    .B1(_0431_),
    .B2(_0434_),
    .ZN(net179));
 BUF_X4 _2173_ (.A(_0348_),
    .Z(_0435_));
 AOI22_X1 _2174_ (.A1(_0248_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0218_),
    .ZN(_0436_));
 OAI21_X1 _2175_ (.A(_0372_),
    .B1(_0373_),
    .B2(_1394_),
    .ZN(_0437_));
 BUF_X4 _2176_ (.A(_0378_),
    .Z(_0438_));
 BUF_X4 _2177_ (.A(_0360_),
    .Z(_0439_));
 NOR3_X4 _2178_ (.A1(_1367_),
    .A2(_0024_),
    .A3(_0397_),
    .ZN(_0440_));
 AND2_X1 _2179_ (.A1(_1373_),
    .A2(\input_buffer[1][19] ),
    .ZN(_0441_));
 AOI221_X2 _2180_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0440_),
    .C1(_0441_),
    .C2(_0386_),
    .ZN(_0442_));
 OAI21_X1 _2181_ (.A(_0436_),
    .B1(_0437_),
    .B2(_0442_),
    .ZN(net180));
 AOI22_X1 _2182_ (.A1(_0250_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0220_),
    .ZN(_0443_));
 CLKBUF_X3 _2183_ (.A(_0371_),
    .Z(_0444_));
 CLKBUF_X3 _2184_ (.A(_0353_),
    .Z(_0445_));
 OAI21_X1 _2185_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1396_),
    .ZN(_0446_));
 NOR3_X4 _2186_ (.A1(_0403_),
    .A2(_0006_),
    .A3(_0419_),
    .ZN(_0447_));
 AND2_X1 _2187_ (.A1(_0426_),
    .A2(\input_buffer[1][1] ),
    .ZN(_0448_));
 AOI221_X2 _2188_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0447_),
    .C1(_0448_),
    .C2(_0386_),
    .ZN(_0449_));
 OAI21_X1 _2189_ (.A(_0443_),
    .B1(_0446_),
    .B2(_0449_),
    .ZN(net181));
 AOI22_X1 _2190_ (.A1(_0251_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0221_),
    .ZN(_0450_));
 OAI21_X1 _2191_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1397_),
    .ZN(_0451_));
 INV_X1 _2192_ (.A(_0025_),
    .ZN(_0452_));
 NAND2_X1 _2193_ (.A1(_1364_),
    .A2(_0452_),
    .ZN(_0453_));
 NOR2_X2 _2194_ (.A1(_0397_),
    .A2(_0453_),
    .ZN(_0454_));
 AND2_X1 _2195_ (.A1(_0283_),
    .A2(\input_buffer[1][20] ),
    .ZN(_0455_));
 BUF_X4 _2196_ (.A(_0385_),
    .Z(_0456_));
 AOI221_X2 _2197_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0454_),
    .C1(_0455_),
    .C2(_0456_),
    .ZN(_0457_));
 OAI21_X1 _2198_ (.A(_0450_),
    .B1(_0451_),
    .B2(_0457_),
    .ZN(net182));
 AOI22_X1 _2199_ (.A1(_0252_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0222_),
    .ZN(_0458_));
 OAI21_X1 _2200_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1398_),
    .ZN(_0459_));
 NOR3_X2 _2201_ (.A1(_0403_),
    .A2(_0026_),
    .A3(_0419_),
    .ZN(_0460_));
 AND2_X1 _2202_ (.A1(_0426_),
    .A2(\input_buffer[1][21] ),
    .ZN(_0461_));
 AOI221_X2 _2203_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0460_),
    .C1(_0461_),
    .C2(_0456_),
    .ZN(_0462_));
 OAI21_X1 _2204_ (.A(_0458_),
    .B1(_0459_),
    .B2(_0462_),
    .ZN(net183));
 AOI22_X1 _2205_ (.A1(_0253_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0223_),
    .ZN(_0463_));
 OAI21_X1 _2206_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1399_),
    .ZN(_0464_));
 NOR3_X2 _2207_ (.A1(_0403_),
    .A2(_0027_),
    .A3(_0419_),
    .ZN(_0465_));
 AND2_X1 _2208_ (.A1(_0426_),
    .A2(\input_buffer[1][22] ),
    .ZN(_0466_));
 AOI221_X2 _2209_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0465_),
    .C1(_0466_),
    .C2(_0456_),
    .ZN(_0467_));
 OAI21_X1 _2210_ (.A(_0463_),
    .B1(_0464_),
    .B2(_0467_),
    .ZN(net184));
 AOI22_X1 _2211_ (.A1(_0254_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_0224_),
    .ZN(_0468_));
 OAI21_X1 _2212_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1400_),
    .ZN(_0469_));
 NOR3_X4 _2213_ (.A1(_0403_),
    .A2(_0028_),
    .A3(_0419_),
    .ZN(_0470_));
 AND2_X2 _2214_ (.A1(_0426_),
    .A2(\input_buffer[1][23] ),
    .ZN(_0471_));
 AOI221_X2 _2215_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0470_),
    .C1(_0471_),
    .C2(_0456_),
    .ZN(_0472_));
 OAI21_X1 _2216_ (.A(_0468_),
    .B1(_0469_),
    .B2(_0472_),
    .ZN(net185));
 AOI22_X1 _2217_ (.A1(_1277_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_1300_),
    .ZN(_0473_));
 OAI21_X1 _2218_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1314_),
    .ZN(_0474_));
 NOR2_X1 _2219_ (.A1(_0357_),
    .A2(_0380_),
    .ZN(_0475_));
 INV_X1 _2220_ (.A(_0029_),
    .ZN(_0476_));
 NAND2_X1 _2221_ (.A1(_1364_),
    .A2(_0476_),
    .ZN(_0477_));
 NOR2_X1 _2222_ (.A1(_0359_),
    .A2(_0477_),
    .ZN(_0478_));
 AOI221_X2 _2223_ (.A(_0356_),
    .B1(_0475_),
    .B2(_0478_),
    .C1(_0359_),
    .C2(_1333_),
    .ZN(_0479_));
 OAI21_X1 _2224_ (.A(_0473_),
    .B1(_0474_),
    .B2(_0479_),
    .ZN(net186));
 AOI22_X1 _2225_ (.A1(_1279_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_1305_),
    .ZN(_0480_));
 OAI21_X1 _2226_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1316_),
    .ZN(_0481_));
 NOR3_X2 _2227_ (.A1(_1366_),
    .A2(_0030_),
    .A3(_0419_),
    .ZN(_0482_));
 AND2_X1 _2228_ (.A1(_0426_),
    .A2(_1335_),
    .ZN(_0483_));
 AOI221_X2 _2229_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0482_),
    .C1(_0483_),
    .C2(_0456_),
    .ZN(_0484_));
 OAI21_X1 _2230_ (.A(_0480_),
    .B1(_0481_),
    .B2(_0484_),
    .ZN(net187));
 AOI22_X1 _2231_ (.A1(_1278_),
    .A2(_0429_),
    .B1(_0435_),
    .B2(_1295_),
    .ZN(_0485_));
 OAI21_X1 _2232_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1317_),
    .ZN(_0486_));
 INV_X1 _2233_ (.A(_0031_),
    .ZN(_0487_));
 NAND2_X1 _2234_ (.A1(_1364_),
    .A2(_0487_),
    .ZN(_0488_));
 NOR4_X1 _2235_ (.A1(_0357_),
    .A2(_0380_),
    .A3(_0359_),
    .A4(_0488_),
    .ZN(_0489_));
 NOR3_X1 _2236_ (.A1(_1339_),
    .A2(_0296_),
    .A3(_0358_),
    .ZN(_0490_));
 NOR3_X1 _2237_ (.A1(_0379_),
    .A2(_0489_),
    .A3(_0490_),
    .ZN(_0491_));
 OAI21_X1 _2238_ (.A(_0485_),
    .B1(_0486_),
    .B2(_0491_),
    .ZN(net188));
 AOI21_X1 _2239_ (.A(_0370_),
    .B1(_0356_),
    .B2(_1326_),
    .ZN(_0492_));
 NOR2_X2 _2240_ (.A1(_1366_),
    .A2(_0000_),
    .ZN(_0493_));
 OAI211_X2 _2241_ (.A(_1359_),
    .B(_0493_),
    .C1(_1360_),
    .C2(_1351_),
    .ZN(_0494_));
 NAND2_X1 _2242_ (.A1(_0283_),
    .A2(_1338_),
    .ZN(_0495_));
 BUF_X4 _2243_ (.A(_1341_),
    .Z(_0496_));
 OAI33_X1 _2244_ (.A1(_0357_),
    .A2(_0359_),
    .A3(_0494_),
    .B1(_0495_),
    .B2(_0496_),
    .B3(_0364_),
    .ZN(_0497_));
 OAI21_X1 _2245_ (.A(_0492_),
    .B1(_0497_),
    .B2(_0379_),
    .ZN(_0498_));
 AOI21_X1 _2246_ (.A(_0343_),
    .B1(_0370_),
    .B2(_1302_),
    .ZN(_0499_));
 AOI22_X2 _2247_ (.A1(_1287_),
    .A2(_0344_),
    .B1(_0498_),
    .B2(_0499_),
    .ZN(net189));
 CLKBUF_X3 _2248_ (.A(_1365_),
    .Z(_0500_));
 OR2_X1 _2249_ (.A1(_0500_),
    .A2(_0001_),
    .ZN(_0501_));
 NOR3_X1 _2250_ (.A1(_0370_),
    .A2(_0356_),
    .A3(_0359_),
    .ZN(_0502_));
 NAND3_X2 _2251_ (.A1(_0351_),
    .A2(_0475_),
    .A3(_0502_),
    .ZN(_0503_));
 NOR2_X1 _2252_ (.A1(_0501_),
    .A2(_0503_),
    .ZN(net190));
 OR2_X1 _2253_ (.A1(_0500_),
    .A2(_0002_),
    .ZN(_0504_));
 NOR2_X1 _2254_ (.A1(_0503_),
    .A2(_0504_),
    .ZN(net191));
 AOI22_X1 _2255_ (.A1(_0256_),
    .A2(_0343_),
    .B1(_0435_),
    .B2(_0226_),
    .ZN(_0505_));
 OAI21_X1 _2256_ (.A(_0444_),
    .B1(_0445_),
    .B2(_1402_),
    .ZN(_0506_));
 NOR3_X2 _2257_ (.A1(_1366_),
    .A2(_0007_),
    .A3(_0419_),
    .ZN(_0507_));
 AND2_X1 _2258_ (.A1(_0426_),
    .A2(\input_buffer[1][2] ),
    .ZN(_0508_));
 AOI221_X2 _2259_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0507_),
    .C1(_0508_),
    .C2(_0456_),
    .ZN(_0509_));
 OAI21_X1 _2260_ (.A(_0505_),
    .B1(_0506_),
    .B2(_0509_),
    .ZN(net192));
 OR2_X1 _2261_ (.A1(_0500_),
    .A2(_0003_),
    .ZN(_0510_));
 NOR2_X1 _2262_ (.A1(_0503_),
    .A2(_0510_),
    .ZN(net193));
 OR2_X1 _2263_ (.A1(_0500_),
    .A2(_0004_),
    .ZN(_0511_));
 NOR2_X1 _2264_ (.A1(_0503_),
    .A2(_0511_),
    .ZN(net194));
 AOI22_X1 _2265_ (.A1(_0257_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0227_),
    .ZN(_0512_));
 OAI21_X1 _2266_ (.A(_0444_),
    .B1(_0445_),
    .B2(_0197_),
    .ZN(_0513_));
 NOR3_X4 _2267_ (.A1(_1367_),
    .A2(_0008_),
    .A3(_0397_),
    .ZN(_0514_));
 AND2_X1 _2268_ (.A1(_1373_),
    .A2(\input_buffer[1][3] ),
    .ZN(_0515_));
 AOI221_X2 _2269_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0514_),
    .C1(_0515_),
    .C2(_0456_),
    .ZN(_0516_));
 OAI21_X1 _2270_ (.A(_0512_),
    .B1(_0513_),
    .B2(_0516_),
    .ZN(net195));
 AOI22_X1 _2271_ (.A1(_0258_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0228_),
    .ZN(_0517_));
 OAI21_X1 _2272_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0198_),
    .ZN(_0518_));
 NOR3_X2 _2273_ (.A1(_1366_),
    .A2(_0009_),
    .A3(_0419_),
    .ZN(_0519_));
 AND2_X1 _2274_ (.A1(_0426_),
    .A2(\input_buffer[1][4] ),
    .ZN(_0520_));
 AOI221_X2 _2275_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0519_),
    .C1(_0520_),
    .C2(_0456_),
    .ZN(_0521_));
 OAI21_X1 _2276_ (.A(_0517_),
    .B1(_0518_),
    .B2(_0521_),
    .ZN(net196));
 AOI22_X1 _2277_ (.A1(_0259_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0229_),
    .ZN(_0522_));
 OAI21_X1 _2278_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0199_),
    .ZN(_0523_));
 NOR3_X4 _2279_ (.A1(_1367_),
    .A2(_0010_),
    .A3(_0397_),
    .ZN(_0524_));
 AND2_X1 _2280_ (.A1(_1373_),
    .A2(\input_buffer[1][5] ),
    .ZN(_0525_));
 AOI221_X2 _2281_ (.A(_0378_),
    .B1(_0360_),
    .B2(_0524_),
    .C1(_0525_),
    .C2(_0456_),
    .ZN(_0526_));
 OAI21_X1 _2282_ (.A(_0522_),
    .B1(_0523_),
    .B2(_0526_),
    .ZN(net197));
 AOI22_X1 _2283_ (.A1(_0260_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0230_),
    .ZN(_0527_));
 OAI21_X1 _2284_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0200_),
    .ZN(_0528_));
 NOR3_X4 _2285_ (.A1(_1366_),
    .A2(_0011_),
    .A3(_1361_),
    .ZN(_0529_));
 AND2_X2 _2286_ (.A1(_0426_),
    .A2(\input_buffer[1][6] ),
    .ZN(_0530_));
 AOI221_X2 _2287_ (.A(_0378_),
    .B1(_0360_),
    .B2(_0529_),
    .C1(_0530_),
    .C2(_0456_),
    .ZN(_0531_));
 OAI21_X1 _2288_ (.A(_0527_),
    .B1(_0528_),
    .B2(_0531_),
    .ZN(net198));
 AOI22_X1 _2289_ (.A1(_0261_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0231_),
    .ZN(_0532_));
 OAI21_X1 _2290_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0201_),
    .ZN(_0533_));
 NOR3_X2 _2291_ (.A1(_1367_),
    .A2(_0012_),
    .A3(_0397_),
    .ZN(_0534_));
 AND2_X1 _2292_ (.A1(_1373_),
    .A2(\input_buffer[1][7] ),
    .ZN(_0535_));
 AOI221_X1 _2293_ (.A(_0378_),
    .B1(_0360_),
    .B2(_0534_),
    .C1(_0535_),
    .C2(_0385_),
    .ZN(_0536_));
 OAI21_X1 _2294_ (.A(_0532_),
    .B1(_0533_),
    .B2(_0536_),
    .ZN(net199));
 AOI22_X1 _2295_ (.A1(_0262_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0232_),
    .ZN(_0537_));
 OAI21_X1 _2296_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0202_),
    .ZN(_0538_));
 NOR3_X2 _2297_ (.A1(_1367_),
    .A2(_0013_),
    .A3(_0397_),
    .ZN(_0539_));
 AND2_X1 _2298_ (.A1(_1373_),
    .A2(\input_buffer[1][8] ),
    .ZN(_0540_));
 AOI221_X2 _2299_ (.A(_0378_),
    .B1(_0360_),
    .B2(_0539_),
    .C1(_0540_),
    .C2(_0385_),
    .ZN(_0541_));
 OAI21_X1 _2300_ (.A(_0537_),
    .B1(_0538_),
    .B2(_0541_),
    .ZN(net200));
 AOI22_X1 _2301_ (.A1(_0263_),
    .A2(_0343_),
    .B1(_0348_),
    .B2(_0233_),
    .ZN(_0542_));
 OAI21_X1 _2302_ (.A(_0371_),
    .B1(_0353_),
    .B2(_0203_),
    .ZN(_0543_));
 NOR2_X1 _2303_ (.A1(_1366_),
    .A2(_0014_),
    .ZN(_0544_));
 AND2_X1 _2304_ (.A1(_1543_),
    .A2(_0544_),
    .ZN(_0545_));
 AND2_X1 _2305_ (.A1(_1373_),
    .A2(\input_buffer[1][9] ),
    .ZN(_0546_));
 AOI221_X1 _2306_ (.A(_0378_),
    .B1(_0360_),
    .B2(_0545_),
    .C1(_0546_),
    .C2(_0385_),
    .ZN(_0547_));
 OAI21_X1 _2307_ (.A(_0542_),
    .B1(_0543_),
    .B2(_0547_),
    .ZN(net201));
 AND2_X1 _2308_ (.A1(_0330_),
    .A2(_1605_),
    .ZN(_0548_));
 AND2_X1 _2309_ (.A1(_1380_),
    .A2(_1575_),
    .ZN(_0549_));
 AOI22_X1 _2310_ (.A1(_1593_),
    .A2(_0548_),
    .B1(_0549_),
    .B2(_0302_),
    .ZN(_0550_));
 NAND3_X1 _2311_ (.A1(_0284_),
    .A2(_1560_),
    .A3(_1548_),
    .ZN(_0551_));
 NAND3_X1 _2312_ (.A1(_0264_),
    .A2(_1545_),
    .A3(_1533_),
    .ZN(_0552_));
 NAND3_X1 _2313_ (.A1(_0314_),
    .A2(_1590_),
    .A3(_1578_),
    .ZN(_0553_));
 NAND4_X1 _2314_ (.A1(_0550_),
    .A2(_0551_),
    .A3(_0552_),
    .A4(_0553_),
    .ZN(net202));
 OAI22_X4 _2315_ (.A1(_0236_),
    .A2(_1603_),
    .B1(_1573_),
    .B2(_1381_),
    .ZN(_0554_));
 BUF_X4 _2316_ (.A(_0554_),
    .Z(_0555_));
 AOI21_X4 _2317_ (.A(_1362_),
    .B1(_1341_),
    .B2(_1372_),
    .ZN(_0556_));
 BUF_X4 _2318_ (.A(_0556_),
    .Z(_0557_));
 BUF_X4 _2319_ (.A(_0557_),
    .Z(_0558_));
 AOI21_X1 _2320_ (.A(_0555_),
    .B1(_0558_),
    .B2(_0362_),
    .ZN(_0559_));
 BUF_X4 _2321_ (.A(_0496_),
    .Z(_0560_));
 INV_X1 _2322_ (.A(_0365_),
    .ZN(_0561_));
 NOR2_X2 _2323_ (.A1(_0206_),
    .A2(_1588_),
    .ZN(_0562_));
 BUF_X4 _2324_ (.A(_0562_),
    .Z(_0563_));
 AOI22_X2 _2325_ (.A1(_0560_),
    .A2(_0561_),
    .B1(_0563_),
    .B2(_0204_),
    .ZN(_0564_));
 NAND2_X1 _2326_ (.A1(_0235_),
    .A2(_1285_),
    .ZN(_0565_));
 BUF_X4 _2327_ (.A(_0565_),
    .Z(_0566_));
 BUF_X4 _2328_ (.A(_0566_),
    .Z(_0567_));
 NAND2_X4 _2329_ (.A1(_0205_),
    .A2(_1299_),
    .ZN(_0568_));
 CLKBUF_X3 _2330_ (.A(_0568_),
    .Z(_0569_));
 OAI211_X4 _2331_ (.A(_1380_),
    .B(_1322_),
    .C1(_1588_),
    .C2(_0206_),
    .ZN(_0570_));
 CLKBUF_X3 _2332_ (.A(_0570_),
    .Z(_0571_));
 OAI221_X2 _2333_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0204_),
    .C1(_0571_),
    .C2(_1379_),
    .ZN(_0572_));
 NOR2_X2 _2334_ (.A1(_0236_),
    .A2(_1603_),
    .ZN(_0573_));
 CLKBUF_X3 _2335_ (.A(_0573_),
    .Z(_0574_));
 NAND2_X1 _2336_ (.A1(_0234_),
    .A2(_0574_),
    .ZN(_0575_));
 AOI22_X2 _2337_ (.A1(_0559_),
    .A2(_0564_),
    .B1(_0572_),
    .B2(_0575_),
    .ZN(net204));
 CLKBUF_X3 _2338_ (.A(_0264_),
    .Z(_0576_));
 NAND3_X1 _2339_ (.A1(_0576_),
    .A2(_0381_),
    .A3(_0558_),
    .ZN(_0577_));
 AOI221_X1 _2340_ (.A(_0555_),
    .B1(_0563_),
    .B2(_0209_),
    .C1(_0560_),
    .C2(_0384_),
    .ZN(_0578_));
 OAI221_X1 _2341_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0209_),
    .C1(_0571_),
    .C2(_1385_),
    .ZN(_0579_));
 NAND2_X1 _2342_ (.A1(_0239_),
    .A2(_0574_),
    .ZN(_0580_));
 AOI22_X1 _2343_ (.A1(_0577_),
    .A2(_0578_),
    .B1(_0579_),
    .B2(_0580_),
    .ZN(net205));
 AOI21_X1 _2344_ (.A(_0555_),
    .B1(_0558_),
    .B2(_0390_),
    .ZN(_0581_));
 NOR2_X1 _2345_ (.A1(_1558_),
    .A2(_0392_),
    .ZN(_0582_));
 AOI21_X1 _2346_ (.A(_0582_),
    .B1(_0563_),
    .B2(_0210_),
    .ZN(_0583_));
 OAI221_X1 _2347_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0210_),
    .C1(_0571_),
    .C2(_1386_),
    .ZN(_0584_));
 NAND2_X1 _2348_ (.A1(_0240_),
    .A2(_0574_),
    .ZN(_0585_));
 AOI22_X1 _2349_ (.A1(_0581_),
    .A2(_0583_),
    .B1(_0584_),
    .B2(_0585_),
    .ZN(net206));
 INV_X1 _2350_ (.A(_0017_),
    .ZN(_0586_));
 NAND3_X1 _2351_ (.A1(_0576_),
    .A2(_0586_),
    .A3(_0558_),
    .ZN(_0587_));
 AOI221_X1 _2352_ (.A(_0555_),
    .B1(_0563_),
    .B2(_0211_),
    .C1(_0560_),
    .C2(_0399_),
    .ZN(_0588_));
 OAI221_X1 _2353_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0211_),
    .C1(_0571_),
    .C2(_1387_),
    .ZN(_0589_));
 NAND2_X1 _2354_ (.A1(_0241_),
    .A2(_0574_),
    .ZN(_0590_));
 AOI22_X1 _2355_ (.A1(_0587_),
    .A2(_0588_),
    .B1(_0589_),
    .B2(_0590_),
    .ZN(net207));
 INV_X1 _2356_ (.A(_0018_),
    .ZN(_0591_));
 NAND3_X1 _2357_ (.A1(_0576_),
    .A2(_0591_),
    .A3(_0558_),
    .ZN(_0592_));
 AOI221_X1 _2358_ (.A(_0555_),
    .B1(_0563_),
    .B2(_0212_),
    .C1(_0560_),
    .C2(_0405_),
    .ZN(_0593_));
 OAI221_X1 _2359_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0212_),
    .C1(_0571_),
    .C2(_1388_),
    .ZN(_0594_));
 NAND2_X1 _2360_ (.A1(_0242_),
    .A2(_0574_),
    .ZN(_0595_));
 AOI22_X1 _2361_ (.A1(_0592_),
    .A2(_0593_),
    .B1(_0594_),
    .B2(_0595_),
    .ZN(net208));
 INV_X1 _2362_ (.A(_0019_),
    .ZN(_0596_));
 NAND3_X1 _2363_ (.A1(_0576_),
    .A2(_0596_),
    .A3(_0558_),
    .ZN(_0597_));
 AOI221_X2 _2364_ (.A(_0555_),
    .B1(_0563_),
    .B2(_0213_),
    .C1(_0560_),
    .C2(_0410_),
    .ZN(_0598_));
 OAI221_X1 _2365_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0213_),
    .C1(_0571_),
    .C2(_1389_),
    .ZN(_0599_));
 NAND2_X1 _2366_ (.A1(_0243_),
    .A2(_0574_),
    .ZN(_0600_));
 AOI22_X1 _2367_ (.A1(_0597_),
    .A2(_0598_),
    .B1(_0599_),
    .B2(_0600_),
    .ZN(net209));
 INV_X1 _2368_ (.A(_0020_),
    .ZN(_0601_));
 NAND3_X1 _2369_ (.A1(_0576_),
    .A2(_0601_),
    .A3(_0558_),
    .ZN(_0602_));
 AOI221_X2 _2370_ (.A(_0555_),
    .B1(_0563_),
    .B2(_0214_),
    .C1(_0560_),
    .C2(_0415_),
    .ZN(_0603_));
 OAI221_X2 _2371_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0214_),
    .C1(_0571_),
    .C2(_1390_),
    .ZN(_0604_));
 CLKBUF_X3 _2372_ (.A(_0573_),
    .Z(_0605_));
 NAND2_X1 _2373_ (.A1(_0244_),
    .A2(_0605_),
    .ZN(_0606_));
 AOI22_X2 _2374_ (.A1(_0602_),
    .A2(_0603_),
    .B1(_0604_),
    .B2(_0606_),
    .ZN(net210));
 INV_X1 _2375_ (.A(_0021_),
    .ZN(_0607_));
 NAND3_X1 _2376_ (.A1(_0576_),
    .A2(_0607_),
    .A3(_0558_),
    .ZN(_0608_));
 BUF_X4 _2377_ (.A(_0562_),
    .Z(_0609_));
 BUF_X4 _2378_ (.A(_0609_),
    .Z(_0610_));
 AOI221_X1 _2379_ (.A(_0555_),
    .B1(_0610_),
    .B2(_0215_),
    .C1(_0560_),
    .C2(_0421_),
    .ZN(_0611_));
 OAI221_X1 _2380_ (.A(_0567_),
    .B1(_0569_),
    .B2(_0215_),
    .C1(_0571_),
    .C2(_1391_),
    .ZN(_0612_));
 NAND2_X1 _2381_ (.A1(_0245_),
    .A2(_0605_),
    .ZN(_0613_));
 AOI22_X1 _2382_ (.A1(_0608_),
    .A2(_0611_),
    .B1(_0612_),
    .B2(_0613_),
    .ZN(net211));
 INV_X1 _2383_ (.A(_0022_),
    .ZN(_0614_));
 NAND3_X1 _2384_ (.A1(_0576_),
    .A2(_0614_),
    .A3(_0558_),
    .ZN(_0615_));
 BUF_X4 _2385_ (.A(_0554_),
    .Z(_0616_));
 AOI221_X1 _2386_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0216_),
    .C1(_0560_),
    .C2(_0427_),
    .ZN(_0617_));
 BUF_X4 _2387_ (.A(_0565_),
    .Z(_0618_));
 OAI221_X1 _2388_ (.A(_0618_),
    .B1(_0569_),
    .B2(_0216_),
    .C1(_0571_),
    .C2(_1392_),
    .ZN(_0619_));
 NAND2_X1 _2389_ (.A1(_0246_),
    .A2(_0605_),
    .ZN(_0620_));
 AOI22_X1 _2390_ (.A1(_0615_),
    .A2(_0617_),
    .B1(_0619_),
    .B2(_0620_),
    .ZN(net212));
 INV_X1 _2391_ (.A(_0023_),
    .ZN(_0621_));
 NAND3_X1 _2392_ (.A1(_0576_),
    .A2(_0621_),
    .A3(_0558_),
    .ZN(_0622_));
 BUF_X4 _2393_ (.A(_0496_),
    .Z(_0623_));
 AOI221_X2 _2394_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0217_),
    .C1(_0623_),
    .C2(_0433_),
    .ZN(_0624_));
 OAI221_X1 _2395_ (.A(_0618_),
    .B1(_0569_),
    .B2(_0217_),
    .C1(_0571_),
    .C2(_1393_),
    .ZN(_0625_));
 NAND2_X1 _2396_ (.A1(_0247_),
    .A2(_0605_),
    .ZN(_0626_));
 AOI22_X1 _2397_ (.A1(_0622_),
    .A2(_0624_),
    .B1(_0625_),
    .B2(_0626_),
    .ZN(net213));
 INV_X1 _2398_ (.A(_0024_),
    .ZN(_0627_));
 BUF_X4 _2399_ (.A(_0557_),
    .Z(_0628_));
 NAND3_X1 _2400_ (.A1(_0576_),
    .A2(_0627_),
    .A3(_0628_),
    .ZN(_0629_));
 AOI221_X2 _2401_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0218_),
    .C1(_0623_),
    .C2(_0441_),
    .ZN(_0630_));
 BUF_X4 _2402_ (.A(_0568_),
    .Z(_0631_));
 BUF_X4 _2403_ (.A(_0570_),
    .Z(_0632_));
 OAI221_X2 _2404_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0218_),
    .C1(_0632_),
    .C2(_1394_),
    .ZN(_0633_));
 NAND2_X1 _2405_ (.A1(_0248_),
    .A2(_0605_),
    .ZN(_0634_));
 AOI22_X2 _2406_ (.A1(_0629_),
    .A2(_0630_),
    .B1(_0633_),
    .B2(_0634_),
    .ZN(net214));
 CLKBUF_X3 _2407_ (.A(_0264_),
    .Z(_0635_));
 INV_X1 _2408_ (.A(_0006_),
    .ZN(_0636_));
 NAND3_X1 _2409_ (.A1(_0635_),
    .A2(_0636_),
    .A3(_0628_),
    .ZN(_0637_));
 AOI221_X1 _2410_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0220_),
    .C1(_0623_),
    .C2(_0448_),
    .ZN(_0638_));
 OAI221_X1 _2411_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0220_),
    .C1(_0632_),
    .C2(_1396_),
    .ZN(_0639_));
 NAND2_X1 _2412_ (.A1(_0250_),
    .A2(_0605_),
    .ZN(_0640_));
 AOI22_X1 _2413_ (.A1(_0637_),
    .A2(_0638_),
    .B1(_0639_),
    .B2(_0640_),
    .ZN(net215));
 NAND3_X1 _2414_ (.A1(_0635_),
    .A2(_0452_),
    .A3(_0628_),
    .ZN(_0641_));
 AOI221_X1 _2415_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0221_),
    .C1(_0623_),
    .C2(_0455_),
    .ZN(_0642_));
 OAI221_X1 _2416_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0221_),
    .C1(_0632_),
    .C2(_1397_),
    .ZN(_0643_));
 NAND2_X1 _2417_ (.A1(_0251_),
    .A2(_0605_),
    .ZN(_0644_));
 AOI22_X1 _2418_ (.A1(_0641_),
    .A2(_0642_),
    .B1(_0643_),
    .B2(_0644_),
    .ZN(net216));
 INV_X1 _2419_ (.A(_0026_),
    .ZN(_0645_));
 NAND3_X1 _2420_ (.A1(_0635_),
    .A2(_0645_),
    .A3(_0628_),
    .ZN(_0646_));
 AOI221_X1 _2421_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0222_),
    .C1(_0623_),
    .C2(_0461_),
    .ZN(_0647_));
 OAI221_X1 _2422_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0222_),
    .C1(_0632_),
    .C2(_1398_),
    .ZN(_0648_));
 NAND2_X1 _2423_ (.A1(_0252_),
    .A2(_0605_),
    .ZN(_0649_));
 AOI22_X1 _2424_ (.A1(_0646_),
    .A2(_0647_),
    .B1(_0648_),
    .B2(_0649_),
    .ZN(net217));
 INV_X1 _2425_ (.A(_0027_),
    .ZN(_0650_));
 NAND3_X1 _2426_ (.A1(_0635_),
    .A2(_0650_),
    .A3(_0628_),
    .ZN(_0651_));
 AOI221_X1 _2427_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0223_),
    .C1(_0623_),
    .C2(_0466_),
    .ZN(_0652_));
 OAI221_X1 _2428_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0223_),
    .C1(_0632_),
    .C2(_1399_),
    .ZN(_0653_));
 NAND2_X1 _2429_ (.A1(_0253_),
    .A2(_0605_),
    .ZN(_0654_));
 AOI22_X1 _2430_ (.A1(_0651_),
    .A2(_0652_),
    .B1(_0653_),
    .B2(_0654_),
    .ZN(net218));
 INV_X1 _2431_ (.A(_0028_),
    .ZN(_0655_));
 NAND3_X1 _2432_ (.A1(_0635_),
    .A2(_0655_),
    .A3(_0628_),
    .ZN(_0656_));
 AOI221_X2 _2433_ (.A(_0616_),
    .B1(_0610_),
    .B2(_0224_),
    .C1(_0623_),
    .C2(_0471_),
    .ZN(_0657_));
 OAI221_X2 _2434_ (.A(_0618_),
    .B1(_0631_),
    .B2(_0224_),
    .C1(_0632_),
    .C2(_1400_),
    .ZN(_0658_));
 NAND2_X1 _2435_ (.A1(_0254_),
    .A2(_0605_),
    .ZN(_0659_));
 AOI22_X2 _2436_ (.A1(_0656_),
    .A2(_0657_),
    .B1(_0658_),
    .B2(_0659_),
    .ZN(net219));
 NAND3_X1 _2437_ (.A1(_0635_),
    .A2(_0476_),
    .A3(_0628_),
    .ZN(_0660_));
 NOR2_X2 _2438_ (.A1(_1374_),
    .A2(_1342_),
    .ZN(_0661_));
 AOI221_X2 _2439_ (.A(_0616_),
    .B1(_0610_),
    .B2(_1300_),
    .C1(_1333_),
    .C2(_0661_),
    .ZN(_0662_));
 OAI221_X2 _2440_ (.A(_0618_),
    .B1(_0631_),
    .B2(_1300_),
    .C1(_0632_),
    .C2(_1314_),
    .ZN(_0663_));
 CLKBUF_X3 _2441_ (.A(_0573_),
    .Z(_0664_));
 NAND2_X1 _2442_ (.A1(_1277_),
    .A2(_0664_),
    .ZN(_0665_));
 AOI22_X2 _2443_ (.A1(_0660_),
    .A2(_0662_),
    .B1(_0663_),
    .B2(_0665_),
    .ZN(net220));
 INV_X1 _2444_ (.A(_0030_),
    .ZN(_0666_));
 NAND3_X1 _2445_ (.A1(_0635_),
    .A2(_0666_),
    .A3(_0628_),
    .ZN(_0667_));
 AOI221_X2 _2446_ (.A(_0616_),
    .B1(_0609_),
    .B2(_1305_),
    .C1(_0623_),
    .C2(_0483_),
    .ZN(_0668_));
 OAI221_X2 _2447_ (.A(_0618_),
    .B1(_0631_),
    .B2(_1305_),
    .C1(_0632_),
    .C2(_1316_),
    .ZN(_0669_));
 NAND2_X1 _2448_ (.A1(_1279_),
    .A2(_0664_),
    .ZN(_0670_));
 AOI22_X2 _2449_ (.A1(_0667_),
    .A2(_0668_),
    .B1(_0669_),
    .B2(_0670_),
    .ZN(net221));
 NAND3_X1 _2450_ (.A1(_0635_),
    .A2(_0487_),
    .A3(_0628_),
    .ZN(_0671_));
 AOI221_X2 _2451_ (.A(_0554_),
    .B1(_0609_),
    .B2(_1295_),
    .C1(_1336_),
    .C2(_0661_),
    .ZN(_0672_));
 OAI221_X2 _2452_ (.A(_0566_),
    .B1(_0631_),
    .B2(_1295_),
    .C1(_0632_),
    .C2(_1317_),
    .ZN(_0673_));
 NAND2_X1 _2453_ (.A1(_1280_),
    .A2(_0664_),
    .ZN(_0674_));
 AOI22_X2 _2454_ (.A1(_0671_),
    .A2(_0672_),
    .B1(_0673_),
    .B2(_0674_),
    .ZN(net222));
 NOR2_X1 _2455_ (.A1(_1374_),
    .A2(_1347_),
    .ZN(_0675_));
 AOI21_X1 _2456_ (.A(_0555_),
    .B1(_0675_),
    .B2(_0560_),
    .ZN(_0676_));
 AOI22_X2 _2457_ (.A1(_0493_),
    .A2(_0557_),
    .B1(_0563_),
    .B2(_1302_),
    .ZN(_0677_));
 OAI221_X2 _2458_ (.A(_0566_),
    .B1(_0631_),
    .B2(_1302_),
    .C1(_0632_),
    .C2(_1319_),
    .ZN(_0678_));
 NAND2_X1 _2459_ (.A1(_1282_),
    .A2(_0664_),
    .ZN(_0679_));
 AOI22_X2 _2460_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0678_),
    .B2(_0679_),
    .ZN(net223));
 NAND2_X1 _2461_ (.A1(_0330_),
    .A2(\dest_id[4][4] ),
    .ZN(_0680_));
 NOR2_X4 _2462_ (.A1(_1381_),
    .A2(_1573_),
    .ZN(_0681_));
 INV_X1 _2463_ (.A(_0501_),
    .ZN(_0682_));
 AOI221_X2 _2464_ (.A(_0681_),
    .B1(_0557_),
    .B2(_0682_),
    .C1(_0284_),
    .C2(_1329_),
    .ZN(_0683_));
 BUF_X4 _2465_ (.A(_0205_),
    .Z(_0684_));
 AOI22_X4 _2466_ (.A1(_0330_),
    .A2(_1285_),
    .B1(_1299_),
    .B2(_0684_),
    .ZN(_0685_));
 NAND2_X2 _2467_ (.A1(_1380_),
    .A2(_1322_),
    .ZN(_0686_));
 OAI21_X1 _2468_ (.A(_0685_),
    .B1(_0686_),
    .B2(_1310_),
    .ZN(_0687_));
 NAND2_X1 _2469_ (.A1(_0314_),
    .A2(_1290_),
    .ZN(_0688_));
 OAI221_X1 _2470_ (.A(_0680_),
    .B1(_0683_),
    .B2(_0687_),
    .C1(_0688_),
    .C2(_0574_),
    .ZN(net224));
 NAND2_X1 _2471_ (.A1(_0330_),
    .A2(\dest_id[4][5] ),
    .ZN(_0689_));
 INV_X1 _2472_ (.A(_0504_),
    .ZN(_0690_));
 AOI221_X2 _2473_ (.A(_0681_),
    .B1(_0556_),
    .B2(_0690_),
    .C1(_0284_),
    .C2(_1328_),
    .ZN(_0691_));
 OAI21_X1 _2474_ (.A(_0685_),
    .B1(_0686_),
    .B2(_1309_),
    .ZN(_0692_));
 NAND2_X1 _2475_ (.A1(_0314_),
    .A2(_1289_),
    .ZN(_0693_));
 OAI221_X1 _2476_ (.A(_0689_),
    .B1(_0691_),
    .B2(_0692_),
    .C1(_0693_),
    .C2(_0574_),
    .ZN(net225));
 INV_X1 _2477_ (.A(_0007_),
    .ZN(_0694_));
 NAND3_X1 _2478_ (.A1(_0635_),
    .A2(_0694_),
    .A3(_0628_),
    .ZN(_0695_));
 AOI221_X1 _2479_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0226_),
    .C1(_0623_),
    .C2(_0508_),
    .ZN(_0696_));
 OAI221_X1 _2480_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0226_),
    .C1(_0570_),
    .C2(_1402_),
    .ZN(_0697_));
 NAND2_X1 _2481_ (.A1(_0256_),
    .A2(_0664_),
    .ZN(_0698_));
 AOI22_X1 _2482_ (.A1(_0695_),
    .A2(_0696_),
    .B1(_0697_),
    .B2(_0698_),
    .ZN(net226));
 NAND2_X1 _2483_ (.A1(_0330_),
    .A2(\dest_id[4][6] ),
    .ZN(_0699_));
 INV_X1 _2484_ (.A(_0510_),
    .ZN(_0700_));
 AOI221_X2 _2485_ (.A(_0681_),
    .B1(_0556_),
    .B2(_0700_),
    .C1(_0284_),
    .C2(_1331_),
    .ZN(_0701_));
 OAI21_X1 _2486_ (.A(_0685_),
    .B1(_0686_),
    .B2(_1312_),
    .ZN(_0702_));
 NAND2_X1 _2487_ (.A1(_0314_),
    .A2(_1292_),
    .ZN(_0703_));
 OAI221_X1 _2488_ (.A(_0699_),
    .B1(_0701_),
    .B2(_0702_),
    .C1(_0703_),
    .C2(_0574_),
    .ZN(net227));
 NAND2_X1 _2489_ (.A1(_0330_),
    .A2(\dest_id[4][7] ),
    .ZN(_0704_));
 INV_X1 _2490_ (.A(_0511_),
    .ZN(_0705_));
 AOI221_X2 _2491_ (.A(_0681_),
    .B1(_0556_),
    .B2(_0705_),
    .C1(_0284_),
    .C2(_1330_),
    .ZN(_0706_));
 OAI21_X1 _2492_ (.A(_0685_),
    .B1(_0686_),
    .B2(_1311_),
    .ZN(_0707_));
 NAND2_X1 _2493_ (.A1(_0314_),
    .A2(_1291_),
    .ZN(_0708_));
 OAI221_X1 _2494_ (.A(_0704_),
    .B1(_0706_),
    .B2(_0707_),
    .C1(_0708_),
    .C2(_0574_),
    .ZN(net228));
 INV_X1 _2495_ (.A(_0008_),
    .ZN(_0709_));
 NAND3_X1 _2496_ (.A1(_0635_),
    .A2(_0709_),
    .A3(_0557_),
    .ZN(_0710_));
 AOI221_X1 _2497_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0227_),
    .C1(_0623_),
    .C2(_0515_),
    .ZN(_0711_));
 OAI221_X1 _2498_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0227_),
    .C1(_0570_),
    .C2(_0197_),
    .ZN(_0712_));
 NAND2_X1 _2499_ (.A1(_0257_),
    .A2(_0664_),
    .ZN(_0713_));
 AOI22_X1 _2500_ (.A1(_0710_),
    .A2(_0711_),
    .B1(_0712_),
    .B2(_0713_),
    .ZN(net229));
 INV_X1 _2501_ (.A(_0009_),
    .ZN(_0714_));
 NAND3_X1 _2502_ (.A1(_0264_),
    .A2(_0714_),
    .A3(_0557_),
    .ZN(_0715_));
 AOI221_X2 _2503_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0228_),
    .C1(_0496_),
    .C2(_0520_),
    .ZN(_0716_));
 OAI221_X1 _2504_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0228_),
    .C1(_0570_),
    .C2(_0198_),
    .ZN(_0717_));
 NAND2_X1 _2505_ (.A1(_0258_),
    .A2(_0664_),
    .ZN(_0718_));
 AOI22_X1 _2506_ (.A1(_0715_),
    .A2(_0716_),
    .B1(_0717_),
    .B2(_0718_),
    .ZN(net230));
 INV_X1 _2507_ (.A(_0010_),
    .ZN(_0719_));
 NAND3_X1 _2508_ (.A1(_0264_),
    .A2(_0719_),
    .A3(_0557_),
    .ZN(_0720_));
 AOI221_X1 _2509_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0229_),
    .C1(_0496_),
    .C2(_0525_),
    .ZN(_0721_));
 OAI221_X1 _2510_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0229_),
    .C1(_0570_),
    .C2(_0199_),
    .ZN(_0722_));
 NAND2_X1 _2511_ (.A1(_0259_),
    .A2(_0664_),
    .ZN(_0723_));
 AOI22_X1 _2512_ (.A1(_0720_),
    .A2(_0721_),
    .B1(_0722_),
    .B2(_0723_),
    .ZN(net231));
 INV_X1 _2513_ (.A(_0011_),
    .ZN(_0724_));
 NAND3_X1 _2514_ (.A1(_0264_),
    .A2(_0724_),
    .A3(_0557_),
    .ZN(_0725_));
 AOI221_X2 _2515_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0230_),
    .C1(_0496_),
    .C2(_0530_),
    .ZN(_0726_));
 OAI221_X1 _2516_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0230_),
    .C1(_0570_),
    .C2(_0200_),
    .ZN(_0727_));
 NAND2_X1 _2517_ (.A1(_0260_),
    .A2(_0664_),
    .ZN(_0728_));
 AOI22_X1 _2518_ (.A1(_0725_),
    .A2(_0726_),
    .B1(_0727_),
    .B2(_0728_),
    .ZN(net232));
 INV_X1 _2519_ (.A(_0012_),
    .ZN(_0729_));
 NAND3_X1 _2520_ (.A1(_0264_),
    .A2(_0729_),
    .A3(_0557_),
    .ZN(_0730_));
 AOI221_X1 _2521_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0231_),
    .C1(_0496_),
    .C2(_0535_),
    .ZN(_0731_));
 OAI221_X1 _2522_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0231_),
    .C1(_0570_),
    .C2(_0201_),
    .ZN(_0732_));
 NAND2_X1 _2523_ (.A1(_0261_),
    .A2(_0664_),
    .ZN(_0733_));
 AOI22_X1 _2524_ (.A1(_0730_),
    .A2(_0731_),
    .B1(_0732_),
    .B2(_0733_),
    .ZN(net233));
 INV_X1 _2525_ (.A(_0013_),
    .ZN(_0734_));
 NAND3_X1 _2526_ (.A1(_0264_),
    .A2(_0734_),
    .A3(_0557_),
    .ZN(_0735_));
 AOI221_X1 _2527_ (.A(_0554_),
    .B1(_0609_),
    .B2(_0232_),
    .C1(_0496_),
    .C2(_0540_),
    .ZN(_0736_));
 OAI221_X1 _2528_ (.A(_0566_),
    .B1(_0568_),
    .B2(_0232_),
    .C1(_0570_),
    .C2(_0202_),
    .ZN(_0737_));
 NAND2_X1 _2529_ (.A1(_0262_),
    .A2(_0573_),
    .ZN(_0738_));
 AOI22_X1 _2530_ (.A1(_0735_),
    .A2(_0736_),
    .B1(_0737_),
    .B2(_0738_),
    .ZN(net234));
 NAND3_X1 _2531_ (.A1(_0233_),
    .A2(_0567_),
    .A3(_0563_),
    .ZN(_0739_));
 OAI21_X1 _2532_ (.A(_0685_),
    .B1(_0686_),
    .B2(_0203_),
    .ZN(_0740_));
 AOI221_X1 _2533_ (.A(_0681_),
    .B1(_0556_),
    .B2(_0544_),
    .C1(_0496_),
    .C2(_0546_),
    .ZN(_0741_));
 INV_X1 _2534_ (.A(_0263_),
    .ZN(_0742_));
 OAI221_X1 _2535_ (.A(_0739_),
    .B1(_0740_),
    .B2(_0741_),
    .C1(_0742_),
    .C2(_0567_),
    .ZN(net235));
 NOR3_X1 _2536_ (.A1(_0661_),
    .A2(_0555_),
    .A3(_0563_),
    .ZN(_0743_));
 OAI21_X1 _2537_ (.A(_0743_),
    .B1(_1543_),
    .B2(_1367_),
    .ZN(net236));
 NAND2_X1 _2538_ (.A1(_0235_),
    .A2(_1604_),
    .ZN(_0744_));
 CLKBUF_X3 _2539_ (.A(_0744_),
    .Z(_0745_));
 CLKBUF_X3 _2540_ (.A(_0745_),
    .Z(_0746_));
 NOR2_X1 _2541_ (.A1(_0234_),
    .A2(_0746_),
    .ZN(_0747_));
 NAND2_X1 _2542_ (.A1(_1380_),
    .A2(_1574_),
    .ZN(_0748_));
 BUF_X8 _2543_ (.A(_0748_),
    .Z(_0749_));
 BUF_X4 _2544_ (.A(_0749_),
    .Z(_0750_));
 NOR2_X1 _2545_ (.A1(_1379_),
    .A2(_0750_),
    .ZN(_0751_));
 AND2_X4 _2546_ (.A1(_1372_),
    .A2(_1559_),
    .ZN(_0752_));
 BUF_X1 rebuffer5 (.A(_1599_),
    .Z(net343));
 BUF_X4 _2548_ (.A(_0752_),
    .Z(_0754_));
 BUF_X4 _2549_ (.A(_0754_),
    .Z(_0755_));
 NOR3_X1 _2550_ (.A1(_0500_),
    .A2(_0005_),
    .A3(_0754_),
    .ZN(_0756_));
 AOI22_X1 _2551_ (.A1(\input_buffer[1][0] ),
    .A2(_0755_),
    .B1(_0756_),
    .B2(_0270_),
    .ZN(_0757_));
 BUF_X4 _2552_ (.A(_0749_),
    .Z(_0758_));
 AOI221_X1 _2553_ (.A(_0751_),
    .B1(_0757_),
    .B2(_0758_),
    .C1(_0314_),
    .C2(_0326_),
    .ZN(_0759_));
 AND2_X1 _2554_ (.A1(_0205_),
    .A2(_0325_),
    .ZN(_0760_));
 CLKBUF_X2 _2555_ (.A(_0760_),
    .Z(_0761_));
 CLKBUF_X3 _2556_ (.A(_0761_),
    .Z(_0762_));
 AOI21_X1 _2557_ (.A(_0759_),
    .B1(_0762_),
    .B2(_0204_),
    .ZN(_0763_));
 CLKBUF_X3 _2558_ (.A(_0745_),
    .Z(_0764_));
 AOI21_X1 _2559_ (.A(_0747_),
    .B1(_0763_),
    .B2(_0764_),
    .ZN(net238));
 NOR2_X1 _2560_ (.A1(_0239_),
    .A2(_0746_),
    .ZN(_0765_));
 NOR2_X1 _2561_ (.A1(_1385_),
    .A2(_0750_),
    .ZN(_0766_));
 NOR3_X1 _2562_ (.A1(_0500_),
    .A2(_0015_),
    .A3(_0754_),
    .ZN(_0767_));
 AOI22_X1 _2563_ (.A1(\input_buffer[1][10] ),
    .A2(_0755_),
    .B1(_0767_),
    .B2(_0270_),
    .ZN(_0768_));
 AOI221_X1 _2564_ (.A(_0766_),
    .B1(_0768_),
    .B2(_0758_),
    .C1(_0314_),
    .C2(_0326_),
    .ZN(_0769_));
 AOI21_X1 _2565_ (.A(_0769_),
    .B1(_0762_),
    .B2(_0209_),
    .ZN(_0770_));
 AOI21_X1 _2566_ (.A(_0765_),
    .B1(_0770_),
    .B2(_0764_),
    .ZN(net239));
 NOR2_X1 _2567_ (.A1(_0240_),
    .A2(_0746_),
    .ZN(_0771_));
 NOR2_X1 _2568_ (.A1(_1386_),
    .A2(_0750_),
    .ZN(_0772_));
 NOR3_X2 _2569_ (.A1(_0500_),
    .A2(_0016_),
    .A3(_0754_),
    .ZN(_0773_));
 AOI22_X2 _2570_ (.A1(\input_buffer[1][11] ),
    .A2(_0755_),
    .B1(_0773_),
    .B2(_0270_),
    .ZN(_0774_));
 AOI221_X2 _2571_ (.A(_0772_),
    .B1(_0774_),
    .B2(_0758_),
    .C1(_0314_),
    .C2(_0326_),
    .ZN(_0775_));
 AOI21_X1 _2572_ (.A(_0775_),
    .B1(_0762_),
    .B2(_0210_),
    .ZN(_0776_));
 AOI21_X1 _2573_ (.A(_0771_),
    .B1(_0776_),
    .B2(_0764_),
    .ZN(net240));
 NOR2_X1 _2574_ (.A1(_0241_),
    .A2(_0746_),
    .ZN(_0777_));
 NOR2_X1 _2575_ (.A1(_1387_),
    .A2(_0750_),
    .ZN(_0778_));
 NOR3_X1 _2576_ (.A1(_0500_),
    .A2(_0017_),
    .A3(_0754_),
    .ZN(_0779_));
 AOI22_X2 _2577_ (.A1(\input_buffer[1][12] ),
    .A2(_0755_),
    .B1(_0779_),
    .B2(_0270_),
    .ZN(_0780_));
 BUF_X4 _2578_ (.A(_0205_),
    .Z(_0781_));
 AOI221_X2 _2579_ (.A(_0778_),
    .B1(_0780_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0782_));
 AOI21_X1 _2580_ (.A(_0782_),
    .B1(_0762_),
    .B2(_0211_),
    .ZN(_0783_));
 AOI21_X1 _2581_ (.A(_0777_),
    .B1(_0783_),
    .B2(_0764_),
    .ZN(net241));
 NOR2_X1 _2582_ (.A1(_0242_),
    .A2(_0746_),
    .ZN(_0784_));
 NOR2_X1 _2583_ (.A1(_1388_),
    .A2(_0750_),
    .ZN(_0785_));
 NOR3_X1 _2584_ (.A1(_0500_),
    .A2(_0018_),
    .A3(_0754_),
    .ZN(_0786_));
 AOI22_X2 _2585_ (.A1(\input_buffer[1][13] ),
    .A2(_0755_),
    .B1(_0786_),
    .B2(_0270_),
    .ZN(_0787_));
 AOI221_X2 _2586_ (.A(_0785_),
    .B1(_0787_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0788_));
 AOI21_X1 _2587_ (.A(_0788_),
    .B1(_0762_),
    .B2(_0212_),
    .ZN(_0789_));
 AOI21_X1 _2588_ (.A(_0784_),
    .B1(_0789_),
    .B2(_0764_),
    .ZN(net242));
 NOR2_X1 _2589_ (.A1(_0243_),
    .A2(_0746_),
    .ZN(_0790_));
 NOR2_X1 _2590_ (.A1(_1389_),
    .A2(_0750_),
    .ZN(_0791_));
 BUF_X4 _2591_ (.A(_0752_),
    .Z(_0792_));
 NOR3_X1 _2592_ (.A1(_0500_),
    .A2(_0019_),
    .A3(_0792_),
    .ZN(_0793_));
 AOI22_X2 _2593_ (.A1(\input_buffer[1][14] ),
    .A2(_0755_),
    .B1(_0793_),
    .B2(_0270_),
    .ZN(_0794_));
 AOI221_X2 _2594_ (.A(_0791_),
    .B1(_0794_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0795_));
 AOI21_X1 _2595_ (.A(_0795_),
    .B1(_0762_),
    .B2(_0213_),
    .ZN(_0796_));
 AOI21_X1 _2596_ (.A(_0790_),
    .B1(_0796_),
    .B2(_0764_),
    .ZN(net243));
 NOR2_X1 _2597_ (.A1(_0244_),
    .A2(_0746_),
    .ZN(_0797_));
 NOR2_X1 _2598_ (.A1(_1390_),
    .A2(_0750_),
    .ZN(_0798_));
 CLKBUF_X3 _2599_ (.A(_1365_),
    .Z(_0799_));
 NOR3_X1 _2600_ (.A1(_0799_),
    .A2(_0020_),
    .A3(_0792_),
    .ZN(_0800_));
 AOI22_X2 _2601_ (.A1(\input_buffer[1][15] ),
    .A2(_0755_),
    .B1(_0800_),
    .B2(_0270_),
    .ZN(_0801_));
 AOI221_X2 _2602_ (.A(_0798_),
    .B1(_0801_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0802_));
 AOI21_X1 _2603_ (.A(_0802_),
    .B1(_0762_),
    .B2(_0214_),
    .ZN(_0803_));
 AOI21_X1 _2604_ (.A(_0797_),
    .B1(_0803_),
    .B2(_0764_),
    .ZN(net244));
 NOR2_X1 _2605_ (.A1(_0245_),
    .A2(_0746_),
    .ZN(_0804_));
 NOR2_X1 _2606_ (.A1(_1391_),
    .A2(_0750_),
    .ZN(_0805_));
 NOR3_X1 _2607_ (.A1(_0799_),
    .A2(_0021_),
    .A3(_0792_),
    .ZN(_0806_));
 AOI22_X2 _2608_ (.A1(\input_buffer[1][16] ),
    .A2(_0755_),
    .B1(_0806_),
    .B2(_0270_),
    .ZN(_0807_));
 AOI221_X2 _2609_ (.A(_0805_),
    .B1(_0807_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0808_));
 AOI21_X1 _2610_ (.A(_0808_),
    .B1(_0762_),
    .B2(_0215_),
    .ZN(_0809_));
 AOI21_X1 _2611_ (.A(_0804_),
    .B1(_0809_),
    .B2(_0764_),
    .ZN(net245));
 CLKBUF_X3 _2612_ (.A(_0745_),
    .Z(_0810_));
 NOR2_X1 _2613_ (.A1(_0246_),
    .A2(_0810_),
    .ZN(_0811_));
 BUF_X4 _2614_ (.A(_0749_),
    .Z(_0812_));
 NOR2_X1 _2615_ (.A1(_1392_),
    .A2(_0812_),
    .ZN(_0813_));
 NOR3_X1 _2616_ (.A1(_0799_),
    .A2(_0022_),
    .A3(_0792_),
    .ZN(_0814_));
 AOI22_X1 _2617_ (.A1(\input_buffer[1][17] ),
    .A2(_0755_),
    .B1(_0814_),
    .B2(_0270_),
    .ZN(_0815_));
 AOI221_X1 _2618_ (.A(_0813_),
    .B1(_0815_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0326_),
    .ZN(_0816_));
 AOI21_X1 _2619_ (.A(_0816_),
    .B1(_0762_),
    .B2(_0216_),
    .ZN(_0817_));
 AOI21_X1 _2620_ (.A(_0811_),
    .B1(_0817_),
    .B2(_0764_),
    .ZN(net246));
 NOR2_X1 _2621_ (.A1(_0247_),
    .A2(_0810_),
    .ZN(_0818_));
 NOR2_X1 _2622_ (.A1(_1393_),
    .A2(_0812_),
    .ZN(_0819_));
 NOR3_X1 _2623_ (.A1(_0799_),
    .A2(_0023_),
    .A3(_0792_),
    .ZN(_0820_));
 BUF_X4 _2624_ (.A(_0269_),
    .Z(_0821_));
 AOI22_X1 _2625_ (.A1(\input_buffer[1][18] ),
    .A2(_0755_),
    .B1(_0820_),
    .B2(_0821_),
    .ZN(_0822_));
 BUF_X4 _2626_ (.A(_0325_),
    .Z(_0823_));
 AOI221_X1 _2627_ (.A(_0819_),
    .B1(_0822_),
    .B2(_0758_),
    .C1(_0781_),
    .C2(_0823_),
    .ZN(_0824_));
 AOI21_X1 _2628_ (.A(_0824_),
    .B1(_0762_),
    .B2(_0217_),
    .ZN(_0825_));
 AOI21_X1 _2629_ (.A(_0818_),
    .B1(_0825_),
    .B2(_0764_),
    .ZN(net247));
 NOR2_X1 _2630_ (.A1(_0248_),
    .A2(_0810_),
    .ZN(_0826_));
 NOR2_X1 _2631_ (.A1(_1394_),
    .A2(_0812_),
    .ZN(_0827_));
 BUF_X4 _2632_ (.A(_0754_),
    .Z(_0828_));
 NOR3_X1 _2633_ (.A1(_0799_),
    .A2(_0024_),
    .A3(_0792_),
    .ZN(_0829_));
 AOI22_X1 _2634_ (.A1(\input_buffer[1][19] ),
    .A2(_0828_),
    .B1(_0829_),
    .B2(_0821_),
    .ZN(_0830_));
 BUF_X4 _2635_ (.A(_0749_),
    .Z(_0831_));
 AOI221_X1 _2636_ (.A(_0827_),
    .B1(_0830_),
    .B2(_0831_),
    .C1(_0781_),
    .C2(_0823_),
    .ZN(_0832_));
 CLKBUF_X3 _2637_ (.A(_0761_),
    .Z(_0833_));
 AOI21_X1 _2638_ (.A(_0832_),
    .B1(_0833_),
    .B2(_0218_),
    .ZN(_0834_));
 CLKBUF_X3 _2639_ (.A(_0745_),
    .Z(_0835_));
 AOI21_X1 _2640_ (.A(_0826_),
    .B1(_0834_),
    .B2(_0835_),
    .ZN(net248));
 NOR2_X1 _2641_ (.A1(_0250_),
    .A2(_0810_),
    .ZN(_0836_));
 NOR2_X1 _2642_ (.A1(_1396_),
    .A2(_0812_),
    .ZN(_0837_));
 NOR3_X1 _2643_ (.A1(_0799_),
    .A2(_0006_),
    .A3(_0792_),
    .ZN(_0838_));
 AOI22_X1 _2644_ (.A1(\input_buffer[1][1] ),
    .A2(_0828_),
    .B1(_0838_),
    .B2(_0821_),
    .ZN(_0839_));
 AOI221_X1 _2645_ (.A(_0837_),
    .B1(_0839_),
    .B2(_0831_),
    .C1(_0781_),
    .C2(_0823_),
    .ZN(_0840_));
 AOI21_X1 _2646_ (.A(_0840_),
    .B1(_0833_),
    .B2(_0220_),
    .ZN(_0841_));
 AOI21_X1 _2647_ (.A(_0836_),
    .B1(_0841_),
    .B2(_0835_),
    .ZN(net249));
 NOR2_X1 _2648_ (.A1(_0251_),
    .A2(_0810_),
    .ZN(_0842_));
 NOR2_X1 _2649_ (.A1(_1397_),
    .A2(_0812_),
    .ZN(_0843_));
 NOR3_X1 _2650_ (.A1(_0799_),
    .A2(_0025_),
    .A3(_0792_),
    .ZN(_0844_));
 AOI22_X1 _2651_ (.A1(\input_buffer[1][20] ),
    .A2(_0828_),
    .B1(_0844_),
    .B2(_0821_),
    .ZN(_0845_));
 AOI221_X1 _2652_ (.A(_0843_),
    .B1(_0845_),
    .B2(_0831_),
    .C1(_0781_),
    .C2(_0823_),
    .ZN(_0846_));
 AOI21_X1 _2653_ (.A(_0846_),
    .B1(_0833_),
    .B2(_0221_),
    .ZN(_0847_));
 AOI21_X1 _2654_ (.A(_0842_),
    .B1(_0847_),
    .B2(_0835_),
    .ZN(net250));
 NOR2_X1 _2655_ (.A1(_0252_),
    .A2(_0810_),
    .ZN(_0848_));
 NOR2_X1 _2656_ (.A1(_1398_),
    .A2(_0812_),
    .ZN(_0849_));
 NOR3_X1 _2657_ (.A1(_0799_),
    .A2(_0026_),
    .A3(_0792_),
    .ZN(_0850_));
 AOI22_X2 _2658_ (.A1(\input_buffer[1][21] ),
    .A2(_0828_),
    .B1(_0850_),
    .B2(_0821_),
    .ZN(_0851_));
 BUF_X4 _2659_ (.A(_0205_),
    .Z(_0852_));
 AOI221_X2 _2660_ (.A(_0849_),
    .B1(_0851_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0853_));
 AOI21_X1 _2661_ (.A(_0853_),
    .B1(_0833_),
    .B2(_0222_),
    .ZN(_0854_));
 AOI21_X1 _2662_ (.A(_0848_),
    .B1(_0854_),
    .B2(_0835_),
    .ZN(net251));
 NOR2_X1 _2663_ (.A1(_0253_),
    .A2(_0810_),
    .ZN(_0855_));
 NOR2_X1 _2664_ (.A1(_1399_),
    .A2(_0812_),
    .ZN(_0856_));
 NOR3_X1 _2665_ (.A1(_0799_),
    .A2(_0027_),
    .A3(_0792_),
    .ZN(_0857_));
 AOI22_X2 _2666_ (.A1(\input_buffer[1][22] ),
    .A2(_0828_),
    .B1(_0857_),
    .B2(_0821_),
    .ZN(_0858_));
 AOI221_X2 _2667_ (.A(_0856_),
    .B1(_0858_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0859_));
 AOI21_X1 _2668_ (.A(_0859_),
    .B1(_0833_),
    .B2(_0223_),
    .ZN(_0860_));
 AOI21_X1 _2669_ (.A(_0855_),
    .B1(_0860_),
    .B2(_0835_),
    .ZN(net252));
 NOR2_X1 _2670_ (.A1(_0254_),
    .A2(_0810_),
    .ZN(_0861_));
 NOR2_X1 _2671_ (.A1(_1400_),
    .A2(_0812_),
    .ZN(_0862_));
 BUF_X4 _2672_ (.A(_0752_),
    .Z(_0863_));
 NOR3_X2 _2673_ (.A1(_0799_),
    .A2(_0028_),
    .A3(_0863_),
    .ZN(_0864_));
 AOI22_X2 _2674_ (.A1(\input_buffer[1][23] ),
    .A2(_0828_),
    .B1(_0864_),
    .B2(_0821_),
    .ZN(_0865_));
 AOI221_X2 _2675_ (.A(_0862_),
    .B1(_0865_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0866_));
 AOI21_X1 _2676_ (.A(_0866_),
    .B1(_0833_),
    .B2(_0224_),
    .ZN(_0867_));
 AOI21_X1 _2677_ (.A(_0861_),
    .B1(_0867_),
    .B2(_0835_),
    .ZN(net253));
 NOR2_X1 _2678_ (.A1(_1277_),
    .A2(_0810_),
    .ZN(_0868_));
 NOR2_X1 _2679_ (.A1(_1314_),
    .A2(_0812_),
    .ZN(_0869_));
 CLKBUF_X3 _2680_ (.A(_1365_),
    .Z(_0870_));
 NOR3_X1 _2681_ (.A1(_0870_),
    .A2(_0029_),
    .A3(_0863_),
    .ZN(_0871_));
 AOI22_X1 _2682_ (.A1(_1333_),
    .A2(_0828_),
    .B1(_0871_),
    .B2(_0821_),
    .ZN(_0872_));
 AOI221_X1 _2683_ (.A(_0869_),
    .B1(_0872_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0873_));
 AOI21_X1 _2684_ (.A(_0873_),
    .B1(_0833_),
    .B2(_1300_),
    .ZN(_0874_));
 AOI21_X2 _2685_ (.A(_0868_),
    .B1(_0874_),
    .B2(_0835_),
    .ZN(net254));
 NOR2_X1 _2686_ (.A1(_1279_),
    .A2(_0810_),
    .ZN(_0875_));
 NOR2_X1 _2687_ (.A1(_1316_),
    .A2(_0812_),
    .ZN(_0876_));
 NOR3_X1 _2688_ (.A1(_0870_),
    .A2(_0030_),
    .A3(_0863_),
    .ZN(_0877_));
 AOI22_X2 _2689_ (.A1(_1335_),
    .A2(_0828_),
    .B1(_0877_),
    .B2(_0821_),
    .ZN(_0878_));
 AOI221_X2 _2690_ (.A(_0876_),
    .B1(_0878_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0879_));
 AOI21_X1 _2691_ (.A(_0879_),
    .B1(_0833_),
    .B2(_1305_),
    .ZN(_0880_));
 AOI21_X1 _2692_ (.A(_0875_),
    .B1(_0880_),
    .B2(_0835_),
    .ZN(net255));
 CLKBUF_X3 _2693_ (.A(_0745_),
    .Z(_0881_));
 NOR2_X1 _2694_ (.A1(_1280_),
    .A2(_0881_),
    .ZN(_0882_));
 BUF_X4 _2695_ (.A(_0749_),
    .Z(_0883_));
 NOR2_X1 _2696_ (.A1(_1317_),
    .A2(_0883_),
    .ZN(_0884_));
 NOR3_X1 _2697_ (.A1(_0870_),
    .A2(_0031_),
    .A3(_0863_),
    .ZN(_0885_));
 AOI22_X1 _2698_ (.A1(_1336_),
    .A2(_0828_),
    .B1(_0885_),
    .B2(_0821_),
    .ZN(_0886_));
 AOI221_X2 _2699_ (.A(_0884_),
    .B1(_0831_),
    .B2(_0886_),
    .C1(_0852_),
    .C2(_0823_),
    .ZN(_0887_));
 AOI21_X1 _2700_ (.A(_0887_),
    .B1(_0833_),
    .B2(_1295_),
    .ZN(_0888_));
 AOI21_X2 _2701_ (.A(_0882_),
    .B1(_0888_),
    .B2(_0835_),
    .ZN(net256));
 NOR2_X1 _2702_ (.A1(_1282_),
    .A2(_0881_),
    .ZN(_0889_));
 NOR2_X1 _2703_ (.A1(_1319_),
    .A2(_0883_),
    .ZN(_0890_));
 NOR3_X1 _2704_ (.A1(_0870_),
    .A2(_0000_),
    .A3(_0863_),
    .ZN(_0891_));
 BUF_X4 _2705_ (.A(_0269_),
    .Z(_0892_));
 AOI22_X1 _2706_ (.A1(_1338_),
    .A2(_0828_),
    .B1(_0891_),
    .B2(_0892_),
    .ZN(_0893_));
 BUF_X4 _2707_ (.A(_0325_),
    .Z(_0894_));
 AOI221_X1 _2708_ (.A(_0890_),
    .B1(_0893_),
    .B2(_0831_),
    .C1(_0852_),
    .C2(_0894_),
    .ZN(_0895_));
 AOI21_X1 _2709_ (.A(_0895_),
    .B1(_0833_),
    .B2(_1302_),
    .ZN(_0896_));
 AOI21_X1 _2710_ (.A(_0889_),
    .B1(_0896_),
    .B2(_0835_),
    .ZN(net257));
 NOR2_X1 _2711_ (.A1(\dest_id[4][4] ),
    .A2(_0881_),
    .ZN(_0897_));
 NOR2_X1 _2712_ (.A1(_1310_),
    .A2(_0883_),
    .ZN(_0898_));
 BUF_X4 _2713_ (.A(_0754_),
    .Z(_0899_));
 NOR3_X1 _2714_ (.A1(_0870_),
    .A2(_0001_),
    .A3(_0863_),
    .ZN(_0900_));
 AOI22_X2 _2715_ (.A1(_1329_),
    .A2(_0899_),
    .B1(_0900_),
    .B2(_0892_),
    .ZN(_0901_));
 BUF_X4 _2716_ (.A(_0749_),
    .Z(_0902_));
 AOI221_X2 _2717_ (.A(_0898_),
    .B1(_0901_),
    .B2(_0902_),
    .C1(_0852_),
    .C2(_0894_),
    .ZN(_0903_));
 CLKBUF_X3 _2718_ (.A(_0761_),
    .Z(_0904_));
 AOI21_X1 _2719_ (.A(_0903_),
    .B1(_0904_),
    .B2(_1290_),
    .ZN(_0905_));
 CLKBUF_X3 _2720_ (.A(_0745_),
    .Z(_0906_));
 AOI21_X1 _2721_ (.A(_0897_),
    .B1(_0905_),
    .B2(_0906_),
    .ZN(net258));
 NOR2_X1 _2722_ (.A1(\dest_id[4][5] ),
    .A2(_0881_),
    .ZN(_0907_));
 NOR2_X1 _2723_ (.A1(_1309_),
    .A2(_0883_),
    .ZN(_0908_));
 NOR3_X1 _2724_ (.A1(_0870_),
    .A2(_0002_),
    .A3(_0863_),
    .ZN(_0909_));
 AOI22_X2 _2725_ (.A1(_1328_),
    .A2(_0899_),
    .B1(_0909_),
    .B2(_0892_),
    .ZN(_0910_));
 AOI221_X2 _2726_ (.A(_0908_),
    .B1(_0910_),
    .B2(_0902_),
    .C1(_0852_),
    .C2(_0894_),
    .ZN(_0911_));
 AOI21_X1 _2727_ (.A(_0911_),
    .B1(_0904_),
    .B2(_1289_),
    .ZN(_0912_));
 AOI21_X1 _2728_ (.A(_0907_),
    .B1(_0912_),
    .B2(_0906_),
    .ZN(net259));
 NOR2_X1 _2729_ (.A1(_0256_),
    .A2(_0881_),
    .ZN(_0913_));
 NOR2_X1 _2730_ (.A1(_1402_),
    .A2(_0883_),
    .ZN(_0914_));
 NOR3_X1 _2731_ (.A1(_0870_),
    .A2(_0007_),
    .A3(_0863_),
    .ZN(_0915_));
 AOI22_X2 _2732_ (.A1(\input_buffer[1][2] ),
    .A2(_0899_),
    .B1(_0915_),
    .B2(_0892_),
    .ZN(_0916_));
 AOI221_X2 _2733_ (.A(_0914_),
    .B1(_0916_),
    .B2(_0902_),
    .C1(_0852_),
    .C2(_0894_),
    .ZN(_0917_));
 AOI21_X1 _2734_ (.A(_0917_),
    .B1(_0904_),
    .B2(_0226_),
    .ZN(_0918_));
 AOI21_X1 _2735_ (.A(_0913_),
    .B1(_0918_),
    .B2(_0906_),
    .ZN(net260));
 NOR2_X1 _2736_ (.A1(\dest_id[4][6] ),
    .A2(_0881_),
    .ZN(_0919_));
 NOR2_X1 _2737_ (.A1(_1312_),
    .A2(_0883_),
    .ZN(_0920_));
 NOR3_X1 _2738_ (.A1(_0870_),
    .A2(_0003_),
    .A3(_0863_),
    .ZN(_0921_));
 AOI22_X2 _2739_ (.A1(_1331_),
    .A2(_0899_),
    .B1(_0921_),
    .B2(_0892_),
    .ZN(_0922_));
 AOI221_X2 _2740_ (.A(_0920_),
    .B1(_0922_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0923_));
 AOI21_X1 _2741_ (.A(_0923_),
    .B1(_0904_),
    .B2(_1292_),
    .ZN(_0924_));
 AOI21_X1 _2742_ (.A(_0919_),
    .B1(_0924_),
    .B2(_0906_),
    .ZN(net261));
 NOR2_X1 _2743_ (.A1(\dest_id[4][7] ),
    .A2(_0881_),
    .ZN(_0925_));
 NOR2_X1 _2744_ (.A1(_1311_),
    .A2(_0883_),
    .ZN(_0926_));
 NOR3_X1 _2745_ (.A1(_0870_),
    .A2(_0004_),
    .A3(_0863_),
    .ZN(_0927_));
 AOI22_X2 _2746_ (.A1(_1330_),
    .A2(_0899_),
    .B1(_0927_),
    .B2(_0892_),
    .ZN(_0928_));
 AOI221_X2 _2747_ (.A(_0926_),
    .B1(_0928_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0929_));
 AOI21_X1 _2748_ (.A(_0929_),
    .B1(_0904_),
    .B2(_1291_),
    .ZN(_0930_));
 AOI21_X1 _2749_ (.A(_0925_),
    .B1(_0930_),
    .B2(_0906_),
    .ZN(net262));
 NOR2_X1 _2750_ (.A1(_0257_),
    .A2(_0881_),
    .ZN(_0931_));
 NOR2_X1 _2751_ (.A1(_0197_),
    .A2(_0883_),
    .ZN(_0932_));
 NOR3_X1 _2752_ (.A1(_0870_),
    .A2(_0008_),
    .A3(_0752_),
    .ZN(_0933_));
 AOI22_X1 _2753_ (.A1(\input_buffer[1][3] ),
    .A2(_0899_),
    .B1(_0933_),
    .B2(_0892_),
    .ZN(_0934_));
 AOI221_X1 _2754_ (.A(_0932_),
    .B1(_0934_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0935_));
 AOI21_X1 _2755_ (.A(_0935_),
    .B1(_0904_),
    .B2(_0227_),
    .ZN(_0936_));
 AOI21_X1 _2756_ (.A(_0931_),
    .B1(_0936_),
    .B2(_0906_),
    .ZN(net263));
 NOR2_X1 _2757_ (.A1(_0258_),
    .A2(_0881_),
    .ZN(_0937_));
 NOR2_X1 _2758_ (.A1(_0198_),
    .A2(_0883_),
    .ZN(_0938_));
 NOR3_X1 _2759_ (.A1(_1365_),
    .A2(_0009_),
    .A3(_0752_),
    .ZN(_0939_));
 AOI22_X1 _2760_ (.A1(\input_buffer[1][4] ),
    .A2(_0899_),
    .B1(_0939_),
    .B2(_0892_),
    .ZN(_0940_));
 AOI221_X1 _2761_ (.A(_0938_),
    .B1(_0940_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0941_));
 AOI21_X1 _2762_ (.A(_0941_),
    .B1(_0904_),
    .B2(_0228_),
    .ZN(_0942_));
 AOI21_X1 _2763_ (.A(_0937_),
    .B1(_0942_),
    .B2(_0906_),
    .ZN(net264));
 NOR2_X1 _2764_ (.A1(_0259_),
    .A2(_0881_),
    .ZN(_0943_));
 NOR2_X1 _2765_ (.A1(_0199_),
    .A2(_0883_),
    .ZN(_0944_));
 NOR3_X1 _2766_ (.A1(_1365_),
    .A2(_0010_),
    .A3(_0752_),
    .ZN(_0945_));
 AOI22_X1 _2767_ (.A1(\input_buffer[1][5] ),
    .A2(_0899_),
    .B1(_0945_),
    .B2(_0892_),
    .ZN(_0946_));
 AOI221_X1 _2768_ (.A(_0944_),
    .B1(_0946_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0947_));
 AOI21_X1 _2769_ (.A(_0947_),
    .B1(_0904_),
    .B2(_0229_),
    .ZN(_0948_));
 AOI21_X1 _2770_ (.A(_0943_),
    .B1(_0948_),
    .B2(_0906_),
    .ZN(net265));
 NOR2_X1 _2771_ (.A1(_0260_),
    .A2(_0745_),
    .ZN(_0949_));
 NOR2_X1 _2772_ (.A1(_0200_),
    .A2(_0749_),
    .ZN(_0950_));
 NOR3_X1 _2773_ (.A1(_1365_),
    .A2(_0011_),
    .A3(_0752_),
    .ZN(_0951_));
 AOI22_X1 _2774_ (.A1(\input_buffer[1][6] ),
    .A2(_0899_),
    .B1(_0951_),
    .B2(_0892_),
    .ZN(_0952_));
 AOI221_X1 _2775_ (.A(_0950_),
    .B1(_0952_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0894_),
    .ZN(_0953_));
 AOI21_X1 _2776_ (.A(_0953_),
    .B1(_0904_),
    .B2(_0230_),
    .ZN(_0954_));
 AOI21_X1 _2777_ (.A(_0949_),
    .B1(_0954_),
    .B2(_0906_),
    .ZN(net266));
 NOR2_X1 _2778_ (.A1(_0261_),
    .A2(_0745_),
    .ZN(_0955_));
 NOR2_X1 _2779_ (.A1(_0201_),
    .A2(_0749_),
    .ZN(_0956_));
 NOR3_X1 _2780_ (.A1(_1365_),
    .A2(_0012_),
    .A3(_0752_),
    .ZN(_0957_));
 AOI22_X1 _2781_ (.A1(\input_buffer[1][7] ),
    .A2(_0899_),
    .B1(_0957_),
    .B2(_0269_),
    .ZN(_0958_));
 AOI221_X1 _2782_ (.A(_0956_),
    .B1(_0958_),
    .B2(_0902_),
    .C1(_0684_),
    .C2(_0325_),
    .ZN(_0959_));
 AOI21_X1 _2783_ (.A(_0959_),
    .B1(_0904_),
    .B2(_0231_),
    .ZN(_0960_));
 AOI21_X1 _2784_ (.A(_0955_),
    .B1(_0960_),
    .B2(_0906_),
    .ZN(net267));
 NOR2_X1 _2785_ (.A1(_0262_),
    .A2(_0745_),
    .ZN(_0961_));
 NOR2_X1 _2786_ (.A1(_0202_),
    .A2(_0749_),
    .ZN(_0962_));
 NOR3_X1 _2787_ (.A1(_1365_),
    .A2(_0013_),
    .A3(_0752_),
    .ZN(_0963_));
 AOI22_X1 _2788_ (.A1(\input_buffer[1][8] ),
    .A2(_0754_),
    .B1(_0963_),
    .B2(_0269_),
    .ZN(_0964_));
 AOI221_X1 _2789_ (.A(_0962_),
    .B1(_0964_),
    .B2(_0750_),
    .C1(_0684_),
    .C2(_0325_),
    .ZN(_0965_));
 AOI21_X1 _2790_ (.A(_0965_),
    .B1(_0761_),
    .B2(_0232_),
    .ZN(_0966_));
 AOI21_X1 _2791_ (.A(_0961_),
    .B1(_0966_),
    .B2(_0746_),
    .ZN(net268));
 NOR2_X1 _2792_ (.A1(_0263_),
    .A2(_0745_),
    .ZN(_0967_));
 NOR2_X1 _2793_ (.A1(_0203_),
    .A2(_0749_),
    .ZN(_0968_));
 NOR3_X1 _2794_ (.A1(_1365_),
    .A2(_0014_),
    .A3(_0752_),
    .ZN(_0969_));
 AOI22_X1 _2795_ (.A1(\input_buffer[1][9] ),
    .A2(_0754_),
    .B1(_0969_),
    .B2(_0269_),
    .ZN(_0970_));
 AOI221_X1 _2796_ (.A(_0968_),
    .B1(_0970_),
    .B2(_0750_),
    .C1(_0684_),
    .C2(_0325_),
    .ZN(_0971_));
 AOI21_X1 _2797_ (.A(_0971_),
    .B1(_0761_),
    .B2(_0233_),
    .ZN(_0972_));
 AOI21_X1 _2798_ (.A(_0967_),
    .B1(_0972_),
    .B2(_0746_),
    .ZN(net269));
 NOR2_X1 _2799_ (.A1(_1302_),
    .A2(_1590_),
    .ZN(_0973_));
 NAND4_X1 _2800_ (.A1(_1579_),
    .A2(_1296_),
    .A3(_0346_),
    .A4(_0973_),
    .ZN(_0974_));
 INV_X1 _2801_ (.A(_1560_),
    .ZN(_0975_));
 AND4_X1 _2802_ (.A1(_0284_),
    .A2(_0975_),
    .A3(_1549_),
    .A4(_1337_),
    .ZN(_0976_));
 INV_X1 _2803_ (.A(_1545_),
    .ZN(_0977_));
 AND4_X1 _2804_ (.A1(_0264_),
    .A2(_1534_),
    .A3(_0977_),
    .A4(_1360_),
    .ZN(_0978_));
 AOI22_X1 _2805_ (.A1(_1345_),
    .A2(_0976_),
    .B1(_0978_),
    .B2(_1358_),
    .ZN(_0979_));
 INV_X1 _2806_ (.A(_1564_),
    .ZN(_0980_));
 NOR3_X1 _2807_ (.A1(_1575_),
    .A2(_0980_),
    .A3(_1321_),
    .ZN(_0981_));
 NAND3_X1 _2808_ (.A1(_0376_),
    .A2(_0310_),
    .A3(_0981_),
    .ZN(_0982_));
 NAND2_X1 _2809_ (.A1(_0330_),
    .A2(_1594_),
    .ZN(_0983_));
 OR4_X1 _2810_ (.A1(_1605_),
    .A2(_1592_),
    .A3(_0334_),
    .A4(_0983_),
    .ZN(_0984_));
 NAND4_X1 _2811_ (.A1(_0974_),
    .A2(_0979_),
    .A3(_0982_),
    .A4(_0984_),
    .ZN(net270));
 NAND2_X1 _2812_ (.A1(_0235_),
    .A2(_1601_),
    .ZN(_0985_));
 AOI211_X4 _2813_ (.A(_1275_),
    .B(_0985_),
    .C1(_0340_),
    .C2(_0341_),
    .ZN(_0986_));
 BUF_X4 _2814_ (.A(_0986_),
    .Z(_0987_));
 CLKBUF_X3 _2815_ (.A(_0987_),
    .Z(_0988_));
 OAI211_X4 _2816_ (.A(_1586_),
    .B(_0346_),
    .C1(_1298_),
    .C2(_1296_),
    .ZN(_0989_));
 NOR2_X4 _2817_ (.A1(_0989_),
    .A2(_0986_),
    .ZN(_0990_));
 CLKBUF_X3 _2818_ (.A(_0990_),
    .Z(_0991_));
 AOI22_X1 _2819_ (.A1(_0234_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0204_),
    .ZN(_0992_));
 NAND4_X4 _2820_ (.A1(_1380_),
    .A2(_0304_),
    .A3(_1313_),
    .A4(_0352_),
    .ZN(_0993_));
 OAI221_X2 _2821_ (.A(_0989_),
    .B1(_0985_),
    .B2(_1285_),
    .C1(_0993_),
    .C2(_1379_),
    .ZN(_0994_));
 NAND3_X2 _2822_ (.A1(_1380_),
    .A2(_0304_),
    .A3(_1313_),
    .ZN(_0995_));
 AOI21_X4 _2823_ (.A(_0995_),
    .B1(_1327_),
    .B2(_0308_),
    .ZN(_0996_));
 INV_X2 _2824_ (.A(_1541_),
    .ZN(_0997_));
 NAND3_X2 _2825_ (.A1(_1372_),
    .A2(_0288_),
    .A3(net342),
    .ZN(_0998_));
 AOI21_X4 _2826_ (.A(_0998_),
    .B1(_0296_),
    .B2(_0293_),
    .ZN(_0999_));
 NOR2_X4 _2827_ (.A1(_0997_),
    .A2(_0999_),
    .ZN(_1000_));
 INV_X1 _2828_ (.A(_0288_),
    .ZN(_1001_));
 NOR2_X1 _2829_ (.A1(_1001_),
    .A2(_0365_),
    .ZN(_1002_));
 AOI221_X1 _2830_ (.A(_0996_),
    .B1(_1000_),
    .B2(_0363_),
    .C1(_1558_),
    .C2(_1002_),
    .ZN(_1003_));
 OAI21_X1 _2831_ (.A(_0992_),
    .B1(_0994_),
    .B2(_1003_),
    .ZN(net272));
 AOI22_X1 _2832_ (.A1(_0239_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0209_),
    .ZN(_1004_));
 INV_X1 _2833_ (.A(_1586_),
    .ZN(_1005_));
 AOI211_X2 _2834_ (.A(_1005_),
    .B(_0369_),
    .C1(_1308_),
    .C2(_0321_),
    .ZN(_1006_));
 NOR2_X4 _2835_ (.A1(_1006_),
    .A2(_0986_),
    .ZN(_1007_));
 CLKBUF_X3 _2836_ (.A(_1007_),
    .Z(_1008_));
 CLKBUF_X3 _2837_ (.A(_0993_),
    .Z(_1009_));
 OAI21_X1 _2838_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1385_),
    .ZN(_1010_));
 INV_X1 _2839_ (.A(_0304_),
    .ZN(_1011_));
 NOR2_X4 _2840_ (.A1(_1011_),
    .A2(_0377_),
    .ZN(_1012_));
 BUF_X4 _2841_ (.A(_1012_),
    .Z(_1013_));
 NOR2_X2 _2842_ (.A1(_1001_),
    .A2(_1341_),
    .ZN(_1014_));
 BUF_X4 _2843_ (.A(_1014_),
    .Z(_1015_));
 BUF_X4 _2844_ (.A(_1000_),
    .Z(_1016_));
 AOI221_X1 _2845_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0384_),
    .C1(_1016_),
    .C2(_0383_),
    .ZN(_1017_));
 OAI21_X1 _2846_ (.A(_1004_),
    .B1(_1010_),
    .B2(_1017_),
    .ZN(net273));
 AOI22_X1 _2847_ (.A1(_0240_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0210_),
    .ZN(_1018_));
 OAI21_X1 _2848_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1386_),
    .ZN(_1019_));
 NOR2_X1 _2849_ (.A1(_1001_),
    .A2(_0392_),
    .ZN(_1020_));
 AOI221_X2 _2850_ (.A(_0996_),
    .B1(_1020_),
    .B2(_1558_),
    .C1(_0391_),
    .C2(_1000_),
    .ZN(_1021_));
 OAI21_X1 _2851_ (.A(_1018_),
    .B1(_1019_),
    .B2(_1021_),
    .ZN(net274));
 AOI22_X1 _2852_ (.A1(_0241_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0211_),
    .ZN(_1022_));
 OAI21_X1 _2853_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1387_),
    .ZN(_1023_));
 AOI221_X2 _2854_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0399_),
    .C1(_1016_),
    .C2(_0398_),
    .ZN(_1024_));
 OAI21_X1 _2855_ (.A(_1022_),
    .B1(_1023_),
    .B2(_1024_),
    .ZN(net275));
 AOI22_X1 _2856_ (.A1(_0242_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0212_),
    .ZN(_1025_));
 OAI21_X1 _2857_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1388_),
    .ZN(_1026_));
 AOI221_X2 _2858_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0405_),
    .C1(_1016_),
    .C2(_0404_),
    .ZN(_1027_));
 OAI21_X1 _2859_ (.A(_1025_),
    .B1(_1026_),
    .B2(_1027_),
    .ZN(net276));
 AOI22_X1 _2860_ (.A1(_0243_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0213_),
    .ZN(_1028_));
 OAI21_X1 _2861_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1389_),
    .ZN(_1029_));
 AOI221_X2 _2862_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0410_),
    .C1(_1016_),
    .C2(_0409_),
    .ZN(_1030_));
 OAI21_X1 _2863_ (.A(_1028_),
    .B1(_1029_),
    .B2(_1030_),
    .ZN(net277));
 AOI22_X1 _2864_ (.A1(_0244_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0214_),
    .ZN(_1031_));
 OAI21_X1 _2865_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1390_),
    .ZN(_1032_));
 AOI221_X2 _2866_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0415_),
    .C1(_1016_),
    .C2(_0414_),
    .ZN(_1033_));
 OAI21_X1 _2867_ (.A(_1031_),
    .B1(_1032_),
    .B2(_1033_),
    .ZN(net278));
 AOI22_X1 _2868_ (.A1(_0245_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0215_),
    .ZN(_1034_));
 OAI21_X1 _2869_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1391_),
    .ZN(_1035_));
 AOI221_X2 _2870_ (.A(_1013_),
    .B1(_1015_),
    .B2(_0421_),
    .C1(_1016_),
    .C2(_0420_),
    .ZN(_1036_));
 OAI21_X1 _2871_ (.A(_1034_),
    .B1(_1035_),
    .B2(_1036_),
    .ZN(net279));
 AOI22_X1 _2872_ (.A1(_0246_),
    .A2(_0988_),
    .B1(_0991_),
    .B2(_0216_),
    .ZN(_1037_));
 OAI21_X1 _2873_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1392_),
    .ZN(_1038_));
 BUF_X4 _2874_ (.A(_1012_),
    .Z(_1039_));
 AOI221_X1 _2875_ (.A(_1039_),
    .B1(_1015_),
    .B2(_0427_),
    .C1(_1016_),
    .C2(_0425_),
    .ZN(_1040_));
 OAI21_X1 _2876_ (.A(_1037_),
    .B1(_1038_),
    .B2(_1040_),
    .ZN(net280));
 CLKBUF_X3 _2877_ (.A(_0986_),
    .Z(_1041_));
 AOI22_X1 _2878_ (.A1(_0247_),
    .A2(_1041_),
    .B1(_0991_),
    .B2(_0217_),
    .ZN(_1042_));
 OAI21_X1 _2879_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1393_),
    .ZN(_1043_));
 AOI221_X1 _2880_ (.A(_1039_),
    .B1(_1015_),
    .B2(_0433_),
    .C1(_1016_),
    .C2(_0432_),
    .ZN(_1044_));
 OAI21_X1 _2881_ (.A(_1042_),
    .B1(_1043_),
    .B2(_1044_),
    .ZN(net281));
 CLKBUF_X3 _2882_ (.A(_0990_),
    .Z(_1045_));
 AOI22_X1 _2883_ (.A1(_0248_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0218_),
    .ZN(_1046_));
 OAI21_X1 _2884_ (.A(_1008_),
    .B1(_1009_),
    .B2(_1394_),
    .ZN(_1047_));
 AND2_X1 _2885_ (.A1(_0288_),
    .A2(_0441_),
    .ZN(_1048_));
 AOI221_X2 _2886_ (.A(_0996_),
    .B1(_1048_),
    .B2(_1558_),
    .C1(_0440_),
    .C2(_1000_),
    .ZN(_1049_));
 OAI21_X1 _2887_ (.A(_1046_),
    .B1(_1047_),
    .B2(_1049_),
    .ZN(net282));
 AOI22_X1 _2888_ (.A1(_0250_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0220_),
    .ZN(_1050_));
 CLKBUF_X3 _2889_ (.A(_1007_),
    .Z(_1051_));
 CLKBUF_X3 _2890_ (.A(_0993_),
    .Z(_1052_));
 OAI21_X1 _2891_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1396_),
    .ZN(_1053_));
 AOI221_X2 _2892_ (.A(_1039_),
    .B1(_1015_),
    .B2(_0448_),
    .C1(_1016_),
    .C2(_0447_),
    .ZN(_1054_));
 OAI21_X1 _2893_ (.A(_1050_),
    .B1(_1053_),
    .B2(_1054_),
    .ZN(net283));
 AOI22_X1 _2894_ (.A1(_0251_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0221_),
    .ZN(_1055_));
 OAI21_X1 _2895_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1397_),
    .ZN(_1056_));
 AOI221_X2 _2896_ (.A(_1039_),
    .B1(_1015_),
    .B2(_0455_),
    .C1(_1016_),
    .C2(_0454_),
    .ZN(_1057_));
 OAI21_X1 _2897_ (.A(_1055_),
    .B1(_1056_),
    .B2(_1057_),
    .ZN(net284));
 AOI22_X1 _2898_ (.A1(_0252_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0222_),
    .ZN(_1058_));
 OAI21_X1 _2899_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1398_),
    .ZN(_1059_));
 BUF_X4 _2900_ (.A(_1014_),
    .Z(_1060_));
 BUF_X4 _2901_ (.A(_1000_),
    .Z(_1061_));
 AOI221_X1 _2902_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0461_),
    .C1(_1061_),
    .C2(_0460_),
    .ZN(_1062_));
 OAI21_X1 _2903_ (.A(_1058_),
    .B1(_1059_),
    .B2(_1062_),
    .ZN(net285));
 AOI22_X1 _2904_ (.A1(_0253_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0223_),
    .ZN(_1063_));
 OAI21_X1 _2905_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1399_),
    .ZN(_1064_));
 AOI221_X1 _2906_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0466_),
    .C1(_1061_),
    .C2(_0465_),
    .ZN(_1065_));
 OAI21_X1 _2907_ (.A(_1063_),
    .B1(_1064_),
    .B2(_1065_),
    .ZN(net286));
 AOI22_X1 _2908_ (.A1(_0254_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_0224_),
    .ZN(_1066_));
 OAI21_X1 _2909_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1400_),
    .ZN(_1067_));
 AOI221_X2 _2910_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0471_),
    .C1(_1061_),
    .C2(_0470_),
    .ZN(_1068_));
 OAI21_X1 _2911_ (.A(_1066_),
    .B1(_1067_),
    .B2(_1068_),
    .ZN(net287));
 AOI22_X1 _2912_ (.A1(_1277_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_1300_),
    .ZN(_1069_));
 OAI21_X1 _2913_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1314_),
    .ZN(_1070_));
 NOR4_X1 _2914_ (.A1(_0997_),
    .A2(_0380_),
    .A3(_0477_),
    .A4(_0999_),
    .ZN(_1071_));
 AND2_X1 _2915_ (.A1(_1333_),
    .A2(_0999_),
    .ZN(_1072_));
 NOR3_X1 _2916_ (.A1(_1013_),
    .A2(_1071_),
    .A3(_1072_),
    .ZN(_1073_));
 OAI21_X1 _2917_ (.A(_1069_),
    .B1(_1070_),
    .B2(_1073_),
    .ZN(net288));
 AOI22_X1 _2918_ (.A1(_1279_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_1305_),
    .ZN(_1074_));
 OAI21_X1 _2919_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1316_),
    .ZN(_1075_));
 AOI221_X1 _2920_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0483_),
    .C1(_1061_),
    .C2(_0482_),
    .ZN(_1076_));
 OAI21_X1 _2921_ (.A(_1074_),
    .B1(_1075_),
    .B2(_1076_),
    .ZN(net289));
 AOI22_X1 _2922_ (.A1(_1278_),
    .A2(_1041_),
    .B1(_1045_),
    .B2(_1295_),
    .ZN(_1077_));
 OAI21_X1 _2923_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1317_),
    .ZN(_1078_));
 NOR4_X1 _2924_ (.A1(_0997_),
    .A2(_0380_),
    .A3(_0488_),
    .A4(_0999_),
    .ZN(_1079_));
 NOR3_X1 _2925_ (.A1(_1339_),
    .A2(_0296_),
    .A3(_0998_),
    .ZN(_1080_));
 NOR3_X1 _2926_ (.A1(_1013_),
    .A2(_1079_),
    .A3(_1080_),
    .ZN(_1081_));
 OAI21_X1 _2927_ (.A(_1077_),
    .B1(_1078_),
    .B2(_1081_),
    .ZN(net290));
 AOI21_X1 _2928_ (.A(_1006_),
    .B1(_0996_),
    .B2(_1326_),
    .ZN(_1082_));
 OAI33_X1 _2929_ (.A1(_1001_),
    .A2(_0560_),
    .A3(_0495_),
    .B1(_0999_),
    .B2(_0494_),
    .B3(_0997_),
    .ZN(_1083_));
 OAI21_X1 _2930_ (.A(_1082_),
    .B1(_1083_),
    .B2(_1013_),
    .ZN(_1084_));
 AOI21_X1 _2931_ (.A(_0987_),
    .B1(_1006_),
    .B2(_1302_),
    .ZN(_1085_));
 AOI22_X2 _2932_ (.A1(_1287_),
    .A2(_0988_),
    .B1(_1084_),
    .B2(_1085_),
    .ZN(net291));
 NAND3_X1 _2933_ (.A1(_1541_),
    .A2(_1543_),
    .A3(_0989_),
    .ZN(_1086_));
 OR4_X2 _2934_ (.A1(_0999_),
    .A2(_1013_),
    .A3(_0986_),
    .A4(_1086_),
    .ZN(_1087_));
 NOR2_X1 _2935_ (.A1(_0501_),
    .A2(_1087_),
    .ZN(net292));
 NOR2_X1 _2936_ (.A1(_0504_),
    .A2(_1087_),
    .ZN(net293));
 AOI22_X1 _2937_ (.A1(_0256_),
    .A2(_0987_),
    .B1(_1045_),
    .B2(_0226_),
    .ZN(_1088_));
 OAI21_X1 _2938_ (.A(_1051_),
    .B1(_1052_),
    .B2(_1402_),
    .ZN(_1089_));
 AOI221_X1 _2939_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0508_),
    .C1(_1061_),
    .C2(_0507_),
    .ZN(_1090_));
 OAI21_X1 _2940_ (.A(_1088_),
    .B1(_1089_),
    .B2(_1090_),
    .ZN(net294));
 NOR2_X1 _2941_ (.A1(_0510_),
    .A2(_1087_),
    .ZN(net295));
 NOR2_X1 _2942_ (.A1(_0511_),
    .A2(_1087_),
    .ZN(net296));
 AOI22_X1 _2943_ (.A1(_0257_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0227_),
    .ZN(_1091_));
 OAI21_X1 _2944_ (.A(_1051_),
    .B1(_1052_),
    .B2(_0197_),
    .ZN(_1092_));
 AND2_X1 _2945_ (.A1(_0288_),
    .A2(_0515_),
    .ZN(_1093_));
 AOI221_X2 _2946_ (.A(_0996_),
    .B1(_1093_),
    .B2(_1558_),
    .C1(_0514_),
    .C2(_1000_),
    .ZN(_1094_));
 OAI21_X1 _2947_ (.A(_1091_),
    .B1(_1092_),
    .B2(_1094_),
    .ZN(net297));
 AOI22_X1 _2948_ (.A1(_0258_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0228_),
    .ZN(_1095_));
 OAI21_X1 _2949_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0198_),
    .ZN(_1096_));
 AOI221_X1 _2950_ (.A(_1039_),
    .B1(_1060_),
    .B2(_0520_),
    .C1(_1061_),
    .C2(_0519_),
    .ZN(_1097_));
 OAI21_X1 _2951_ (.A(_1095_),
    .B1(_1096_),
    .B2(_1097_),
    .ZN(net298));
 AOI22_X1 _2952_ (.A1(_0259_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0229_),
    .ZN(_1098_));
 OAI21_X1 _2953_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0199_),
    .ZN(_1099_));
 AOI221_X2 _2954_ (.A(_1012_),
    .B1(_1060_),
    .B2(_0525_),
    .C1(_1061_),
    .C2(_0524_),
    .ZN(_1100_));
 OAI21_X1 _2955_ (.A(_1098_),
    .B1(_1099_),
    .B2(_1100_),
    .ZN(net299));
 AOI22_X1 _2956_ (.A1(_0260_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0230_),
    .ZN(_1101_));
 OAI21_X1 _2957_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0200_),
    .ZN(_1102_));
 AOI221_X2 _2958_ (.A(_1012_),
    .B1(_1060_),
    .B2(_0530_),
    .C1(_1061_),
    .C2(_0529_),
    .ZN(_1103_));
 OAI21_X1 _2959_ (.A(_1101_),
    .B1(_1102_),
    .B2(_1103_),
    .ZN(net300));
 AOI22_X1 _2960_ (.A1(_0261_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0231_),
    .ZN(_1104_));
 OAI21_X1 _2961_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0201_),
    .ZN(_1105_));
 AOI221_X1 _2962_ (.A(_1012_),
    .B1(_1060_),
    .B2(_0535_),
    .C1(_1061_),
    .C2(_0534_),
    .ZN(_1106_));
 OAI21_X1 _2963_ (.A(_1104_),
    .B1(_1105_),
    .B2(_1106_),
    .ZN(net301));
 AOI22_X1 _2964_ (.A1(_0262_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0232_),
    .ZN(_1107_));
 OAI21_X1 _2965_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0202_),
    .ZN(_1108_));
 AND2_X1 _2966_ (.A1(_0288_),
    .A2(_0540_),
    .ZN(_1109_));
 AOI221_X1 _2967_ (.A(_0996_),
    .B1(_1109_),
    .B2(_1342_),
    .C1(_0539_),
    .C2(_1000_),
    .ZN(_1110_));
 OAI21_X1 _2968_ (.A(_1107_),
    .B1(_1108_),
    .B2(_1110_),
    .ZN(net302));
 AOI22_X1 _2969_ (.A1(_0263_),
    .A2(_0987_),
    .B1(_0990_),
    .B2(_0233_),
    .ZN(_1111_));
 OAI21_X1 _2970_ (.A(_1007_),
    .B1(_0993_),
    .B2(_0203_),
    .ZN(_1112_));
 AOI221_X1 _2971_ (.A(_1012_),
    .B1(_1060_),
    .B2(_0546_),
    .C1(_1061_),
    .C2(_0545_),
    .ZN(_1113_));
 OAI21_X1 _2972_ (.A(_1111_),
    .B1(_1112_),
    .B2(_1113_),
    .ZN(net303));
 OAI21_X1 _2973_ (.A(_1358_),
    .B1(_1360_),
    .B2(_1357_),
    .ZN(_1114_));
 NOR3_X1 _2974_ (.A1(_1367_),
    .A2(_1534_),
    .A3(_0977_),
    .ZN(_1115_));
 OAI21_X1 _2975_ (.A(_1304_),
    .B1(_1301_),
    .B2(_1296_),
    .ZN(_1116_));
 INV_X1 _2976_ (.A(_1590_),
    .ZN(_1117_));
 NOR3_X1 _2977_ (.A1(_0206_),
    .A2(_1117_),
    .A3(_1579_),
    .ZN(_1118_));
 OAI21_X1 _2978_ (.A(_1345_),
    .B1(_1343_),
    .B2(_1337_),
    .ZN(_1119_));
 NOR3_X1 _2979_ (.A1(_1374_),
    .A2(_0975_),
    .A3(_1549_),
    .ZN(_1120_));
 AOI222_X2 _2980_ (.A1(_1114_),
    .A2(_1115_),
    .B1(_1116_),
    .B2(_1118_),
    .C1(_1119_),
    .C2(_1120_),
    .ZN(_1121_));
 OAI21_X1 _2981_ (.A(_1313_),
    .B1(_1321_),
    .B2(_0310_),
    .ZN(_1122_));
 INV_X1 _2982_ (.A(_1122_),
    .ZN(_1123_));
 NAND2_X1 _2983_ (.A1(_0980_),
    .A2(_0549_),
    .ZN(_1124_));
 INV_X1 _2984_ (.A(_1594_),
    .ZN(_1125_));
 NAND3_X1 _2985_ (.A1(_1125_),
    .A2(_0334_),
    .A3(_0548_),
    .ZN(_1126_));
 OAI221_X1 _2986_ (.A(_1121_),
    .B1(_1123_),
    .B2(_1124_),
    .C1(_1126_),
    .C2(_1592_),
    .ZN(net304));
 NAND3_X4 _2987_ (.A1(_0330_),
    .A2(net343),
    .A3(_1603_),
    .ZN(_1127_));
 NOR2_X1 _2988_ (.A1(_0234_),
    .A2(_1127_),
    .ZN(_1128_));
 AND3_X1 _2989_ (.A1(_0235_),
    .A2(net343),
    .A3(_1603_),
    .ZN(_1129_));
 CLKBUF_X3 _2990_ (.A(_1129_),
    .Z(_1130_));
 INV_X1 _2991_ (.A(_0327_),
    .ZN(_1131_));
 AOI211_X4 _2992_ (.A(_1131_),
    .B(_0369_),
    .C1(_1308_),
    .C2(_0321_),
    .ZN(_1132_));
 AOI21_X1 _2993_ (.A(_1130_),
    .B1(_1132_),
    .B2(_0204_),
    .ZN(_1133_));
 OAI211_X4 _2994_ (.A(_0327_),
    .B(_0346_),
    .C1(_1298_),
    .C2(_1296_),
    .ZN(_1134_));
 OAI211_X4 _2995_ (.A(_0303_),
    .B(_0376_),
    .C1(_1321_),
    .C2(_1318_),
    .ZN(_1135_));
 CLKBUF_X3 _2996_ (.A(_1135_),
    .Z(_1136_));
 OAI211_X2 _2997_ (.A(_0287_),
    .B(net341),
    .C1(_1337_),
    .C2(_1340_),
    .ZN(_1137_));
 OAI21_X1 _2998_ (.A(_1136_),
    .B1(_1137_),
    .B2(_0365_),
    .ZN(_1138_));
 AND3_X1 _2999_ (.A1(_1373_),
    .A2(_0287_),
    .A3(net340),
    .ZN(_1139_));
 OAI21_X4 _3000_ (.A(_1139_),
    .B1(_1340_),
    .B2(_1337_),
    .ZN(_1140_));
 AND4_X1 _3001_ (.A1(_0268_),
    .A2(_1543_),
    .A3(_0362_),
    .A4(_1140_),
    .ZN(_1141_));
 OAI221_X1 _3002_ (.A(_1134_),
    .B1(_1138_),
    .B2(_1141_),
    .C1(_1379_),
    .C2(_1136_),
    .ZN(_1142_));
 AOI21_X1 _3003_ (.A(_1128_),
    .B1(_1133_),
    .B2(_1142_),
    .ZN(net306));
 NOR2_X1 _3004_ (.A1(_0239_),
    .A2(_1127_),
    .ZN(_1143_));
 AOI21_X1 _3005_ (.A(_1130_),
    .B1(_1132_),
    .B2(_0209_),
    .ZN(_1144_));
 INV_X2 _3006_ (.A(_0268_),
    .ZN(_1145_));
 NAND3_X1 _3007_ (.A1(_1372_),
    .A2(_0287_),
    .A3(_1332_),
    .ZN(_1146_));
 AOI21_X4 _3008_ (.A(_1146_),
    .B1(_0296_),
    .B2(_0293_),
    .ZN(_1147_));
 NOR4_X1 _3009_ (.A1(_1145_),
    .A2(_0380_),
    .A3(_0382_),
    .A4(_1147_),
    .ZN(_1148_));
 NAND2_X1 _3010_ (.A1(_0284_),
    .A2(\input_buffer[1][10] ),
    .ZN(_1149_));
 OAI21_X1 _3011_ (.A(_1136_),
    .B1(_1137_),
    .B2(_1149_),
    .ZN(_1150_));
 OAI221_X1 _3012_ (.A(_1134_),
    .B1(_1148_),
    .B2(_1150_),
    .C1(_1136_),
    .C2(_1385_),
    .ZN(_1151_));
 AOI21_X1 _3013_ (.A(_1143_),
    .B1(_1144_),
    .B2(_1151_),
    .ZN(net307));
 NOR2_X1 _3014_ (.A1(_0240_),
    .A2(_1127_),
    .ZN(_1152_));
 AOI21_X1 _3015_ (.A(_1130_),
    .B1(_1132_),
    .B2(_0210_),
    .ZN(_1153_));
 AND4_X1 _3016_ (.A1(_0268_),
    .A2(_1543_),
    .A3(_0390_),
    .A4(_1140_),
    .ZN(_1154_));
 OAI21_X1 _3017_ (.A(_1136_),
    .B1(_1137_),
    .B2(_0392_),
    .ZN(_1155_));
 OAI221_X1 _3018_ (.A(_1134_),
    .B1(_1154_),
    .B2(_1155_),
    .C1(_1136_),
    .C2(_1386_),
    .ZN(_1156_));
 AOI21_X1 _3019_ (.A(_1152_),
    .B1(_1153_),
    .B2(_1156_),
    .ZN(net308));
 NAND2_X1 _3020_ (.A1(_0235_),
    .A2(_1599_),
    .ZN(_1157_));
 AOI211_X4 _3021_ (.A(_1275_),
    .B(_1157_),
    .C1(_0340_),
    .C2(_0341_),
    .ZN(_1158_));
 CLKBUF_X3 _3022_ (.A(_1158_),
    .Z(_1159_));
 NOR2_X2 _3023_ (.A1(_1134_),
    .A2(_1158_),
    .ZN(_1160_));
 CLKBUF_X3 _3024_ (.A(_1160_),
    .Z(_1161_));
 AOI22_X1 _3025_ (.A1(_0241_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0211_),
    .ZN(_1162_));
 NOR2_X2 _3026_ (.A1(_1132_),
    .A2(_1158_),
    .ZN(_1163_));
 CLKBUF_X3 _3027_ (.A(_1163_),
    .Z(_1164_));
 INV_X1 _3028_ (.A(_0303_),
    .ZN(_1165_));
 NOR3_X2 _3029_ (.A1(_1381_),
    .A2(_1165_),
    .A3(_1323_),
    .ZN(_1166_));
 NAND2_X2 _3030_ (.A1(_0352_),
    .A2(_1166_),
    .ZN(_1167_));
 CLKBUF_X3 _3031_ (.A(_1167_),
    .Z(_1168_));
 OAI21_X1 _3032_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1387_),
    .ZN(_1169_));
 NOR2_X4 _3033_ (.A1(_1165_),
    .A2(_0377_),
    .ZN(_1170_));
 BUF_X4 _3034_ (.A(_1170_),
    .Z(_1171_));
 AND2_X1 _3035_ (.A1(_0287_),
    .A2(_1342_),
    .ZN(_1172_));
 BUF_X4 _3036_ (.A(_1172_),
    .Z(_1173_));
 BUF_X4 _3037_ (.A(_1173_),
    .Z(_1174_));
 NOR2_X2 _3038_ (.A1(_1145_),
    .A2(_1147_),
    .ZN(_1175_));
 BUF_X4 _3039_ (.A(_1175_),
    .Z(_1176_));
 AOI221_X2 _3040_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0399_),
    .C1(_1176_),
    .C2(_0398_),
    .ZN(_1177_));
 OAI21_X1 _3041_ (.A(_1162_),
    .B1(_1169_),
    .B2(_1177_),
    .ZN(net309));
 AOI22_X1 _3042_ (.A1(_0242_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0212_),
    .ZN(_1178_));
 OAI21_X1 _3043_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1388_),
    .ZN(_1179_));
 AOI221_X2 _3044_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0405_),
    .C1(_1176_),
    .C2(_0404_),
    .ZN(_1180_));
 OAI21_X1 _3045_ (.A(_1178_),
    .B1(_1179_),
    .B2(_1180_),
    .ZN(net310));
 AOI22_X1 _3046_ (.A1(_0243_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0213_),
    .ZN(_1181_));
 OAI21_X1 _3047_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1389_),
    .ZN(_1182_));
 AOI221_X2 _3048_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0410_),
    .C1(_1176_),
    .C2(_0409_),
    .ZN(_1183_));
 OAI21_X1 _3049_ (.A(_1181_),
    .B1(_1182_),
    .B2(_1183_),
    .ZN(net311));
 AOI22_X1 _3050_ (.A1(_0244_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0214_),
    .ZN(_1184_));
 OAI21_X1 _3051_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1390_),
    .ZN(_1185_));
 AOI221_X2 _3052_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0415_),
    .C1(_1176_),
    .C2(_0414_),
    .ZN(_1186_));
 OAI21_X1 _3053_ (.A(_1184_),
    .B1(_1185_),
    .B2(_1186_),
    .ZN(net312));
 AOI22_X1 _3054_ (.A1(_0245_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0215_),
    .ZN(_1187_));
 OAI21_X1 _3055_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1391_),
    .ZN(_1188_));
 AOI221_X2 _3056_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0421_),
    .C1(_1176_),
    .C2(_0420_),
    .ZN(_1189_));
 OAI21_X1 _3057_ (.A(_1187_),
    .B1(_1188_),
    .B2(_1189_),
    .ZN(net313));
 AOI22_X1 _3058_ (.A1(_0246_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0216_),
    .ZN(_1190_));
 OAI21_X1 _3059_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1392_),
    .ZN(_1191_));
 AOI221_X1 _3060_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0427_),
    .C1(_1176_),
    .C2(_0425_),
    .ZN(_1192_));
 OAI21_X1 _3061_ (.A(_1190_),
    .B1(_1191_),
    .B2(_1192_),
    .ZN(net314));
 AOI22_X1 _3062_ (.A1(_0247_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0217_),
    .ZN(_1193_));
 OAI21_X1 _3063_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1393_),
    .ZN(_1194_));
 AOI221_X1 _3064_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0433_),
    .C1(_1176_),
    .C2(_0432_),
    .ZN(_1195_));
 OAI21_X1 _3065_ (.A(_1193_),
    .B1(_1194_),
    .B2(_1195_),
    .ZN(net315));
 AOI22_X1 _3066_ (.A1(_0248_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0218_),
    .ZN(_1196_));
 OAI21_X1 _3067_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1394_),
    .ZN(_1197_));
 AOI221_X1 _3068_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0441_),
    .C1(_1176_),
    .C2(_0440_),
    .ZN(_1198_));
 OAI21_X1 _3069_ (.A(_1196_),
    .B1(_1197_),
    .B2(_1198_),
    .ZN(net316));
 AOI22_X1 _3070_ (.A1(_0250_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0220_),
    .ZN(_1199_));
 OAI21_X1 _3071_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1396_),
    .ZN(_1200_));
 AOI221_X1 _3072_ (.A(_1171_),
    .B1(_1174_),
    .B2(_0448_),
    .C1(_1176_),
    .C2(_0447_),
    .ZN(_1201_));
 OAI21_X1 _3073_ (.A(_1199_),
    .B1(_1200_),
    .B2(_1201_),
    .ZN(net317));
 NOR2_X1 _3074_ (.A1(_0251_),
    .A2(_1127_),
    .ZN(_1202_));
 AOI21_X1 _3075_ (.A(_1130_),
    .B1(_1132_),
    .B2(_0221_),
    .ZN(_1203_));
 NOR4_X1 _3076_ (.A1(_1145_),
    .A2(_0380_),
    .A3(_0453_),
    .A4(_1147_),
    .ZN(_1204_));
 NAND2_X1 _3077_ (.A1(_0284_),
    .A2(\input_buffer[1][20] ),
    .ZN(_1205_));
 OAI21_X1 _3078_ (.A(_1135_),
    .B1(_1137_),
    .B2(_1205_),
    .ZN(_1206_));
 OAI221_X1 _3079_ (.A(_1134_),
    .B1(_1204_),
    .B2(_1206_),
    .C1(_1136_),
    .C2(_1397_),
    .ZN(_1207_));
 AOI21_X1 _3080_ (.A(_1202_),
    .B1(_1203_),
    .B2(_1207_),
    .ZN(net318));
 AOI22_X1 _3081_ (.A1(_0252_),
    .A2(_1159_),
    .B1(_1161_),
    .B2(_0222_),
    .ZN(_1208_));
 OAI21_X1 _3082_ (.A(_1164_),
    .B1(_1168_),
    .B2(_1398_),
    .ZN(_1209_));
 AOI221_X1 _3083_ (.A(_1170_),
    .B1(_1174_),
    .B2(_0461_),
    .C1(_1176_),
    .C2(_0460_),
    .ZN(_1210_));
 OAI21_X1 _3084_ (.A(_1208_),
    .B1(_1209_),
    .B2(_1210_),
    .ZN(net319));
 CLKBUF_X3 _3085_ (.A(_1158_),
    .Z(_1211_));
 CLKBUF_X3 _3086_ (.A(_1160_),
    .Z(_1212_));
 AOI22_X1 _3087_ (.A1(_0253_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0223_),
    .ZN(_1213_));
 CLKBUF_X3 _3088_ (.A(_1163_),
    .Z(_1214_));
 CLKBUF_X3 _3089_ (.A(_1167_),
    .Z(_1215_));
 OAI21_X1 _3090_ (.A(_1214_),
    .B1(_1215_),
    .B2(_1399_),
    .ZN(_1216_));
 BUF_X4 _3091_ (.A(_1175_),
    .Z(_1217_));
 AOI221_X1 _3092_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0466_),
    .C1(_1217_),
    .C2(_0465_),
    .ZN(_1218_));
 OAI21_X1 _3093_ (.A(_1213_),
    .B1(_1216_),
    .B2(_1218_),
    .ZN(net320));
 AOI22_X1 _3094_ (.A1(_0254_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0224_),
    .ZN(_1219_));
 OAI21_X1 _3095_ (.A(_1214_),
    .B1(_1215_),
    .B2(_1400_),
    .ZN(_1220_));
 AOI221_X1 _3096_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0471_),
    .C1(_1217_),
    .C2(_0470_),
    .ZN(_1221_));
 OAI21_X1 _3097_ (.A(_1219_),
    .B1(_1220_),
    .B2(_1221_),
    .ZN(net321));
 NOR4_X2 _3098_ (.A1(_1145_),
    .A2(_0380_),
    .A3(_0477_),
    .A4(_1147_),
    .ZN(_1222_));
 OAI21_X1 _3099_ (.A(_1135_),
    .B1(_1140_),
    .B2(_1334_),
    .ZN(_1223_));
 OAI221_X2 _3100_ (.A(_1134_),
    .B1(_1222_),
    .B2(_1223_),
    .C1(_1136_),
    .C2(_1314_),
    .ZN(_1224_));
 AOI21_X1 _3101_ (.A(_1130_),
    .B1(_1132_),
    .B2(_1300_),
    .ZN(_1225_));
 AOI22_X2 _3102_ (.A1(_1278_),
    .A2(_1130_),
    .B1(_1224_),
    .B2(_1225_),
    .ZN(net322));
 AOI22_X1 _3103_ (.A1(_1279_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_1305_),
    .ZN(_1226_));
 OAI21_X1 _3104_ (.A(_1214_),
    .B1(_1215_),
    .B2(_1316_),
    .ZN(_1227_));
 AOI221_X1 _3105_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0483_),
    .C1(_1217_),
    .C2(_0482_),
    .ZN(_1228_));
 OAI21_X1 _3106_ (.A(_1226_),
    .B1(_1227_),
    .B2(_1228_),
    .ZN(net323));
 AOI22_X1 _3107_ (.A1(_1280_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_1295_),
    .ZN(_1229_));
 OAI21_X1 _3108_ (.A(_1214_),
    .B1(_1215_),
    .B2(_1315_),
    .ZN(_1230_));
 NOR2_X1 _3109_ (.A1(_1339_),
    .A2(_1140_),
    .ZN(_1231_));
 NOR4_X1 _3110_ (.A1(_1145_),
    .A2(_0380_),
    .A3(_0488_),
    .A4(_1147_),
    .ZN(_1232_));
 NOR3_X1 _3111_ (.A1(_1171_),
    .A2(_1231_),
    .A3(_1232_),
    .ZN(_1233_));
 OAI21_X1 _3112_ (.A(_1229_),
    .B1(_1230_),
    .B2(_1233_),
    .ZN(net324));
 NOR3_X1 _3113_ (.A1(_1145_),
    .A2(_0494_),
    .A3(_1147_),
    .ZN(_1234_));
 NAND2_X1 _3114_ (.A1(_0287_),
    .A2(_0675_),
    .ZN(_1235_));
 OAI21_X1 _3115_ (.A(_1135_),
    .B1(_1235_),
    .B2(_0496_),
    .ZN(_1236_));
 OAI221_X2 _3116_ (.A(_1134_),
    .B1(_1234_),
    .B2(_1236_),
    .C1(_1136_),
    .C2(_1319_),
    .ZN(_1237_));
 AOI21_X1 _3117_ (.A(_1130_),
    .B1(_1132_),
    .B2(_1302_),
    .ZN(_1238_));
 AOI22_X2 _3118_ (.A1(_1287_),
    .A2(_1130_),
    .B1(_1237_),
    .B2(_1238_),
    .ZN(net325));
 NOR3_X2 _3119_ (.A1(_1145_),
    .A2(_0380_),
    .A3(_1132_),
    .ZN(_1239_));
 NAND4_X4 _3120_ (.A1(_1140_),
    .A2(_1136_),
    .A3(_1127_),
    .A4(_1239_),
    .ZN(_1240_));
 NOR2_X1 _3121_ (.A1(_0501_),
    .A2(_1240_),
    .ZN(net326));
 NOR2_X1 _3122_ (.A1(_0504_),
    .A2(_1240_),
    .ZN(net327));
 AOI22_X1 _3123_ (.A1(_0256_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0226_),
    .ZN(_1241_));
 OAI21_X1 _3124_ (.A(_1214_),
    .B1(_1215_),
    .B2(_1402_),
    .ZN(_1242_));
 AOI221_X1 _3125_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0508_),
    .C1(_1217_),
    .C2(_0507_),
    .ZN(_1243_));
 OAI21_X1 _3126_ (.A(_1241_),
    .B1(_1242_),
    .B2(_1243_),
    .ZN(net328));
 NOR2_X1 _3127_ (.A1(_0510_),
    .A2(_1240_),
    .ZN(net329));
 NOR2_X1 _3128_ (.A1(_0511_),
    .A2(_1240_),
    .ZN(net330));
 AOI22_X1 _3129_ (.A1(_0257_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0227_),
    .ZN(_1244_));
 OAI21_X1 _3130_ (.A(_1214_),
    .B1(_1215_),
    .B2(_0197_),
    .ZN(_1245_));
 AOI221_X1 _3131_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0515_),
    .C1(_1217_),
    .C2(_0514_),
    .ZN(_1246_));
 OAI21_X1 _3132_ (.A(_1244_),
    .B1(_1245_),
    .B2(_1246_),
    .ZN(net331));
 AOI22_X1 _3133_ (.A1(_0258_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0228_),
    .ZN(_1247_));
 OAI21_X1 _3134_ (.A(_1214_),
    .B1(_1215_),
    .B2(_0198_),
    .ZN(_1248_));
 AOI221_X1 _3135_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0520_),
    .C1(_1217_),
    .C2(_0519_),
    .ZN(_1249_));
 OAI21_X1 _3136_ (.A(_1247_),
    .B1(_1248_),
    .B2(_1249_),
    .ZN(net332));
 AOI22_X1 _3137_ (.A1(_0259_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0229_),
    .ZN(_1250_));
 OAI21_X1 _3138_ (.A(_1214_),
    .B1(_1215_),
    .B2(_0199_),
    .ZN(_1251_));
 AND2_X1 _3139_ (.A1(_0352_),
    .A2(_1166_),
    .ZN(_1252_));
 AND2_X1 _3140_ (.A1(_0287_),
    .A2(_0525_),
    .ZN(_1253_));
 AOI221_X2 _3141_ (.A(_1252_),
    .B1(_1253_),
    .B2(_1342_),
    .C1(_0524_),
    .C2(_1217_),
    .ZN(_1254_));
 OAI21_X1 _3142_ (.A(_1250_),
    .B1(_1251_),
    .B2(_1254_),
    .ZN(net333));
 AOI22_X1 _3143_ (.A1(_0260_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0230_),
    .ZN(_1255_));
 OAI21_X1 _3144_ (.A(_1214_),
    .B1(_1215_),
    .B2(_0200_),
    .ZN(_1256_));
 AOI221_X2 _3145_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0530_),
    .C1(_1217_),
    .C2(_0529_),
    .ZN(_1257_));
 OAI21_X1 _3146_ (.A(_1255_),
    .B1(_1256_),
    .B2(_1257_),
    .ZN(net334));
 AOI22_X1 _3147_ (.A1(_0261_),
    .A2(_1211_),
    .B1(_1212_),
    .B2(_0231_),
    .ZN(_1258_));
 OAI21_X1 _3148_ (.A(_1214_),
    .B1(_1215_),
    .B2(_0201_),
    .ZN(_1259_));
 AND2_X1 _3149_ (.A1(_0287_),
    .A2(_0535_),
    .ZN(_1260_));
 AOI221_X2 _3150_ (.A(_1252_),
    .B1(_1260_),
    .B2(_1342_),
    .C1(_0534_),
    .C2(_1217_),
    .ZN(_1261_));
 OAI21_X1 _3151_ (.A(_1258_),
    .B1(_1259_),
    .B2(_1261_),
    .ZN(net335));
 AOI22_X1 _3152_ (.A1(_0262_),
    .A2(_1158_),
    .B1(_1160_),
    .B2(_0232_),
    .ZN(_1262_));
 OAI21_X1 _3153_ (.A(_1163_),
    .B1(_1167_),
    .B2(_0202_),
    .ZN(_1263_));
 AND2_X1 _3154_ (.A1(_0287_),
    .A2(_0540_),
    .ZN(_1264_));
 AOI221_X1 _3155_ (.A(_1252_),
    .B1(_1264_),
    .B2(_1342_),
    .C1(_0539_),
    .C2(_1175_),
    .ZN(_1265_));
 OAI21_X1 _3156_ (.A(_1262_),
    .B1(_1263_),
    .B2(_1265_),
    .ZN(net336));
 AOI22_X1 _3157_ (.A1(_0263_),
    .A2(_1158_),
    .B1(_1160_),
    .B2(_0233_),
    .ZN(_1266_));
 OAI21_X1 _3158_ (.A(_1163_),
    .B1(_1167_),
    .B2(_0203_),
    .ZN(_1267_));
 AOI221_X1 _3159_ (.A(_1170_),
    .B1(_1173_),
    .B2(_0546_),
    .C1(_1217_),
    .C2(_0545_),
    .ZN(_1268_));
 OAI21_X1 _3160_ (.A(_1266_),
    .B1(_1267_),
    .B2(_1268_),
    .ZN(net337));
 NAND3_X1 _3161_ (.A1(_0576_),
    .A2(_1545_),
    .A3(_0268_),
    .ZN(_1269_));
 NAND2_X1 _3162_ (.A1(net344),
    .A2(_0548_),
    .ZN(_1270_));
 NAND3_X1 _3163_ (.A1(_0314_),
    .A2(_1590_),
    .A3(_0327_),
    .ZN(_1271_));
 AND3_X1 _3164_ (.A1(_0284_),
    .A2(_1560_),
    .A3(_0287_),
    .ZN(_1272_));
 AOI21_X1 _3165_ (.A(_1272_),
    .B1(_0549_),
    .B2(_0303_),
    .ZN(_1273_));
 NAND4_X1 _3166_ (.A1(_1269_),
    .A2(_1270_),
    .A3(_1271_),
    .A4(_1273_),
    .ZN(net338));
 HA_X1 _3167_ (.A(_1531_),
    .B(_1532_),
    .CO(_1533_),
    .S(_1534_));
 HA_X1 _3168_ (.A(_1531_),
    .B(_1535_),
    .CO(_1536_),
    .S(_1537_));
 HA_X1 _3169_ (.A(_1538_),
    .B(_1532_),
    .CO(_1539_),
    .S(_1540_));
 HA_X1 _3170_ (.A(_1538_),
    .B(_1535_),
    .CO(_1541_),
    .S(_1542_));
 HA_X1 _3171_ (.A(_1539_),
    .B(_1543_),
    .CO(_1544_),
    .S(_1545_));
 HA_X1 _3172_ (.A(_1546_),
    .B(_1547_),
    .CO(_1548_),
    .S(_1549_));
 HA_X1 _3173_ (.A(_1546_),
    .B(_1550_),
    .CO(_1551_),
    .S(_1552_));
 HA_X1 _3174_ (.A(_1553_),
    .B(_1547_),
    .CO(_1554_),
    .S(_1555_));
 HA_X1 _3175_ (.A(_1553_),
    .B(_1550_),
    .CO(_1556_),
    .S(_1557_));
 HA_X1 _3176_ (.A(_1551_),
    .B(_1558_),
    .CO(_1559_),
    .S(_1560_));
 HA_X1 _3177_ (.A(_1561_),
    .B(_1562_),
    .CO(_1563_),
    .S(_1564_));
 HA_X1 _3178_ (.A(_1561_),
    .B(_1565_),
    .CO(_1566_),
    .S(_1567_));
 HA_X1 _3179_ (.A(_1568_),
    .B(_1562_),
    .CO(_1569_),
    .S(_1570_));
 HA_X1 _3180_ (.A(_1568_),
    .B(_1565_),
    .CO(_1571_),
    .S(_1572_));
 HA_X1 _3181_ (.A(_1566_),
    .B(_1573_),
    .CO(_1574_),
    .S(_1575_));
 HA_X1 _3182_ (.A(_1576_),
    .B(_1577_),
    .CO(_1578_),
    .S(_1579_));
 HA_X1 _3183_ (.A(_1576_),
    .B(_1580_),
    .CO(_1581_),
    .S(_1582_));
 HA_X1 _3184_ (.A(_1583_),
    .B(_1577_),
    .CO(_1584_),
    .S(_1585_));
 HA_X1 _3185_ (.A(_1583_),
    .B(_1580_),
    .CO(_1586_),
    .S(_1587_));
 HA_X1 _3186_ (.A(_1581_),
    .B(_1588_),
    .CO(_1589_),
    .S(_1590_));
 HA_X1 _3187_ (.A(_1591_),
    .B(_1592_),
    .CO(_1593_),
    .S(_1594_));
 HA_X1 _3188_ (.A(_1591_),
    .B(_1595_),
    .CO(_1596_),
    .S(_1597_));
 HA_X1 _3189_ (.A(_1598_),
    .B(_1592_),
    .CO(_1599_),
    .S(_1600_));
 HA_X1 _3190_ (.A(_1598_),
    .B(_1595_),
    .CO(_1601_),
    .S(_1602_));
 HA_X1 _3191_ (.A(_1596_),
    .B(_1603_),
    .CO(_1604_),
    .S(_1605_));
 DFF_X1 \input_buffer[0][0]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][0] ),
    .QN(_0005_));
 DFF_X1 \input_buffer[0][10]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][10] ),
    .QN(_0015_));
 DFF_X1 \input_buffer[0][11]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][11] ),
    .QN(_0016_));
 DFF_X2 \input_buffer[0][12]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][12] ),
    .QN(_0017_));
 DFF_X2 \input_buffer[0][13]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][13] ),
    .QN(_0018_));
 DFF_X2 \input_buffer[0][14]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][14] ),
    .QN(_0019_));
 DFF_X2 \input_buffer[0][15]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][15] ),
    .QN(_0020_));
 DFF_X2 \input_buffer[0][16]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][16] ),
    .QN(_0021_));
 DFF_X2 \input_buffer[0][17]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][17] ),
    .QN(_0022_));
 DFF_X2 \input_buffer[0][18]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][18] ),
    .QN(_0023_));
 DFF_X2 \input_buffer[0][19]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][19] ),
    .QN(_0024_));
 DFF_X2 \input_buffer[0][1]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[0][1] ),
    .QN(_0006_));
 DFF_X1 \input_buffer[0][20]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][20] ),
    .QN(_0025_));
 DFF_X2 \input_buffer[0][21]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][21] ),
    .QN(_0026_));
 DFF_X2 \input_buffer[0][22]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[0][22] ),
    .QN(_0027_));
 DFF_X2 \input_buffer[0][23]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_4_4_0_clk),
    .Q(\input_buffer[0][23] ),
    .QN(_0028_));
 DFF_X2 \input_buffer[0][24]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_4_4_0_clk),
    .Q(\dest_id[0][0] ),
    .QN(_0029_));
 DFF_X2 \input_buffer[0][25]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_4_1_0_clk),
    .Q(\dest_id[0][1] ),
    .QN(_0030_));
 DFF_X2 \input_buffer[0][26]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_4_1_0_clk),
    .Q(\dest_id[0][2] ),
    .QN(_0031_));
 DFF_X1 \input_buffer[0][27]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_4_1_0_clk),
    .Q(\dest_id[0][3] ),
    .QN(_0000_));
 DFF_X2 \input_buffer[0][28]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[0][4] ),
    .QN(_0001_));
 DFF_X2 \input_buffer[0][29]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[0][5] ),
    .QN(_0002_));
 DFF_X2 \input_buffer[0][2]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer[0][2] ),
    .QN(_0007_));
 DFF_X1 \input_buffer[0][30]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[0][6] ),
    .QN(_0003_));
 DFF_X2 \input_buffer[0][31]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[0][7] ),
    .QN(_0004_));
 DFF_X2 \input_buffer[0][3]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[0][3] ),
    .QN(_0008_));
 DFF_X2 \input_buffer[0][4]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer[0][4] ),
    .QN(_0009_));
 DFF_X2 \input_buffer[0][5]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[0][5] ),
    .QN(_0010_));
 DFF_X2 \input_buffer[0][6]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[0][6] ),
    .QN(_0011_));
 DFF_X2 \input_buffer[0][7]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[0][7] ),
    .QN(_0012_));
 DFF_X2 \input_buffer[0][8]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer[0][8] ),
    .QN(_0013_));
 DFF_X1 \input_buffer[0][9]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_4_3_0_clk),
    .Q(\input_buffer[0][9] ),
    .QN(_0014_));
 DFF_X1 \input_buffer[1][0]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][0] ),
    .QN(_1530_));
 DFF_X1 \input_buffer[1][10]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][10] ),
    .QN(_1529_));
 DFF_X1 \input_buffer[1][11]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][11] ),
    .QN(_1528_));
 DFF_X1 \input_buffer[1][12]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][12] ),
    .QN(_1527_));
 DFF_X1 \input_buffer[1][13]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[1][13] ),
    .QN(_1526_));
 DFF_X1 \input_buffer[1][14]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[1][14] ),
    .QN(_1525_));
 DFF_X1 \input_buffer[1][15]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[1][15] ),
    .QN(_1524_));
 DFF_X1 \input_buffer[1][16]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[1][16] ),
    .QN(_1523_));
 DFF_X1 \input_buffer[1][17]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][17] ),
    .QN(_1522_));
 DFF_X1 \input_buffer[1][18]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_4_6_0_clk),
    .Q(\input_buffer[1][18] ),
    .QN(_1521_));
 DFF_X1 \input_buffer[1][19]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[1][19] ),
    .QN(_1520_));
 DFF_X1 \input_buffer[1][1]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[1][1] ),
    .QN(_1519_));
 DFF_X1 \input_buffer[1][20]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_4_4_0_clk),
    .Q(\input_buffer[1][20] ),
    .QN(_1518_));
 DFF_X2 \input_buffer[1][21]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_4_5_0_clk),
    .Q(\input_buffer[1][21] ),
    .QN(_1517_));
 DFF_X2 \input_buffer[1][22]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_4_4_0_clk),
    .Q(\input_buffer[1][22] ),
    .QN(_1516_));
 DFF_X2 \input_buffer[1][23]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_4_4_0_clk),
    .Q(\input_buffer[1][23] ),
    .QN(_1515_));
 DFF_X1 \input_buffer[1][24]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_4_4_0_clk),
    .Q(\dest_id[1][0] ),
    .QN(_1514_));
 DFF_X1 \input_buffer[1][25]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_4_4_0_clk),
    .Q(\dest_id[1][1] ),
    .QN(_1513_));
 DFF_X1 \input_buffer[1][26]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_4_4_0_clk),
    .Q(\dest_id[1][2] ),
    .QN(_1512_));
 DFF_X1 \input_buffer[1][27]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_4_4_0_clk),
    .Q(\dest_id[1][3] ),
    .QN(_1511_));
 DFF_X1 \input_buffer[1][28]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[1][4] ),
    .QN(_1510_));
 DFF_X1 \input_buffer[1][29]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_4_0_0_clk),
    .Q(\dest_id[1][5] ),
    .QN(_1509_));
 DFF_X2 \input_buffer[1][2]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[1][2] ),
    .QN(_1508_));
 DFF_X1 \input_buffer[1][30]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_4_3_0_clk),
    .Q(\dest_id[1][6] ),
    .QN(_1507_));
 DFF_X1 \input_buffer[1][31]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_4_3_0_clk),
    .Q(\dest_id[1][7] ),
    .QN(_1506_));
 DFF_X1 \input_buffer[1][3]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_4_3_0_clk),
    .Q(\input_buffer[1][3] ),
    .QN(_1505_));
 DFF_X1 \input_buffer[1][4]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[1][4] ),
    .QN(_1504_));
 DFF_X1 \input_buffer[1][5]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_4_3_0_clk),
    .Q(\input_buffer[1][5] ),
    .QN(_1503_));
 DFF_X1 \input_buffer[1][6]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[1][6] ),
    .QN(_1502_));
 DFF_X1 \input_buffer[1][7]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_4_0_0_clk),
    .Q(\input_buffer[1][7] ),
    .QN(_1501_));
 DFF_X1 \input_buffer[1][8]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer[1][8] ),
    .QN(_1500_));
 DFF_X1 \input_buffer[1][9]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer[1][9] ),
    .QN(_1499_));
 DFF_X1 \input_buffer[2][0]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][0] ),
    .QN(_1498_));
 DFF_X1 \input_buffer[2][10]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][10] ),
    .QN(_1497_));
 DFF_X1 \input_buffer[2][11]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][11] ),
    .QN(_1496_));
 DFF_X1 \input_buffer[2][12]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][12] ),
    .QN(_1495_));
 DFF_X1 \input_buffer[2][13]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][13] ),
    .QN(_1494_));
 DFF_X1 \input_buffer[2][14]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[2][14] ),
    .QN(_1493_));
 DFF_X1 \input_buffer[2][15]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[2][15] ),
    .QN(_1492_));
 DFF_X1 \input_buffer[2][16]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[2][16] ),
    .QN(_1491_));
 DFF_X1 \input_buffer[2][17]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[2][17] ),
    .QN(_1490_));
 DFF_X1 \input_buffer[2][18]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[2][18] ),
    .QN(_1489_));
 DFF_X1 \input_buffer[2][19]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[2][19] ),
    .QN(_1488_));
 DFF_X1 \input_buffer[2][1]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[2][1] ),
    .QN(_1487_));
 DFF_X1 \input_buffer[2][20]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[2][20] ),
    .QN(_1486_));
 DFF_X1 \input_buffer[2][21]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[2][21] ),
    .QN(_1485_));
 DFF_X1 \input_buffer[2][22]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[2][22] ),
    .QN(_1484_));
 DFF_X1 \input_buffer[2][23]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[2][23] ),
    .QN(_1483_));
 DFF_X1 \input_buffer[2][24]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[2][0] ),
    .QN(_1482_));
 DFF_X1 \input_buffer[2][25]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[2][1] ),
    .QN(_1481_));
 DFF_X1 \input_buffer[2][26]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[2][2] ),
    .QN(_1480_));
 DFF_X1 \input_buffer[2][27]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[2][3] ),
    .QN(_1479_));
 DFF_X1 \input_buffer[2][28]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_2_0_clk),
    .Q(\dest_id[2][4] ),
    .QN(_1478_));
 DFF_X1 \input_buffer[2][29]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_2_0_clk),
    .Q(\dest_id[2][5] ),
    .QN(_1477_));
 DFF_X1 \input_buffer[2][2]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[2][2] ),
    .QN(_1476_));
 DFF_X1 \input_buffer[2][30]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_2_0_clk),
    .Q(\dest_id[2][6] ),
    .QN(_1475_));
 DFF_X1 \input_buffer[2][31]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_2_0_clk),
    .Q(\dest_id[2][7] ),
    .QN(_1474_));
 DFF_X1 \input_buffer[2][3]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[2][3] ),
    .QN(_1473_));
 DFF_X1 \input_buffer[2][4]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_8_0_clk),
    .Q(\input_buffer[2][4] ),
    .QN(_1472_));
 DFF_X1 \input_buffer[2][5]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_8_0_clk),
    .Q(\input_buffer[2][5] ),
    .QN(_1471_));
 DFF_X1 \input_buffer[2][6]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_8_0_clk),
    .Q(\input_buffer[2][6] ),
    .QN(_1470_));
 DFF_X1 \input_buffer[2][7]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[2][7] ),
    .QN(_1469_));
 DFF_X1 \input_buffer[2][8]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_4_11_0_clk),
    .Q(\input_buffer[2][8] ),
    .QN(_1468_));
 DFF_X1 \input_buffer[2][9]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[2][9] ),
    .QN(_1467_));
 DFF_X1 \input_buffer[3][0]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[3][0] ),
    .QN(_1466_));
 DFF_X1 \input_buffer[3][10]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[3][10] ),
    .QN(_1465_));
 DFF_X1 \input_buffer[3][11]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[3][11] ),
    .QN(_1464_));
 DFF_X1 \input_buffer[3][12]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[3][12] ),
    .QN(_1463_));
 DFF_X1 \input_buffer[3][13]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_4_7_0_clk),
    .Q(\input_buffer[3][13] ),
    .QN(_1462_));
 DFF_X1 \input_buffer[3][14]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[3][14] ),
    .QN(_1461_));
 DFF_X1 \input_buffer[3][15]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[3][15] ),
    .QN(_1460_));
 DFF_X1 \input_buffer[3][16]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[3][16] ),
    .QN(_1459_));
 DFF_X1 \input_buffer[3][17]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[3][17] ),
    .QN(_1458_));
 DFF_X1 \input_buffer[3][18]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[3][18] ),
    .QN(_1457_));
 DFF_X1 \input_buffer[3][19]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[3][19] ),
    .QN(_1456_));
 DFF_X1 \input_buffer[3][1]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[3][1] ),
    .QN(_1455_));
 DFF_X1 \input_buffer[3][20]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[3][20] ),
    .QN(_1454_));
 DFF_X1 \input_buffer[3][21]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[3][21] ),
    .QN(_1453_));
 DFF_X1 \input_buffer[3][22]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[3][22] ),
    .QN(_1452_));
 DFF_X1 \input_buffer[3][23]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[3][23] ),
    .QN(_1451_));
 DFF_X2 \input_buffer[3][24]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[3][0] ),
    .QN(_1450_));
 DFF_X2 \input_buffer[3][25]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[3][1] ),
    .QN(_1449_));
 DFF_X1 \input_buffer[3][26]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_4_14_0_clk),
    .Q(\dest_id[3][2] ),
    .QN(_1448_));
 DFF_X2 \input_buffer[3][27]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[3][3] ),
    .QN(_1447_));
 DFF_X1 \input_buffer[3][28]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[3][4] ),
    .QN(_1446_));
 DFF_X1 \input_buffer[3][29]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_4_2_0_clk),
    .Q(\dest_id[3][5] ),
    .QN(_1445_));
 DFF_X1 \input_buffer[3][2]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[3][2] ),
    .QN(_1444_));
 DFF_X1 \input_buffer[3][30]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[3][6] ),
    .QN(_1443_));
 DFF_X1 \input_buffer[3][31]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[3][7] ),
    .QN(_1442_));
 DFF_X1 \input_buffer[3][3]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[3][3] ),
    .QN(_1441_));
 DFF_X1 \input_buffer[3][4]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[3][4] ),
    .QN(_1440_));
 DFF_X1 \input_buffer[3][5]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[3][5] ),
    .QN(_1439_));
 DFF_X1 \input_buffer[3][6]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[3][6] ),
    .QN(_1438_));
 DFF_X1 \input_buffer[3][7]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[3][7] ),
    .QN(_1437_));
 DFF_X1 \input_buffer[3][8]$_DFFE_PP_  (.D(_0158_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[3][8] ),
    .QN(_1436_));
 DFF_X1 \input_buffer[3][9]$_DFFE_PP_  (.D(_0159_),
    .CK(clknet_4_9_0_clk),
    .Q(\input_buffer[3][9] ),
    .QN(_1435_));
 DFF_X1 \input_buffer[4][0]$_DFFE_PP_  (.D(_0160_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[4][0] ),
    .QN(_1434_));
 DFF_X1 \input_buffer[4][10]$_DFFE_PP_  (.D(_0161_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[4][10] ),
    .QN(_1433_));
 DFF_X1 \input_buffer[4][11]$_DFFE_PP_  (.D(_0162_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][11] ),
    .QN(_1432_));
 DFF_X1 \input_buffer[4][12]$_DFFE_PP_  (.D(_0163_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][12] ),
    .QN(_1431_));
 DFF_X1 \input_buffer[4][13]$_DFFE_PP_  (.D(_0164_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[4][13] ),
    .QN(_1430_));
 DFF_X1 \input_buffer[4][14]$_DFFE_PP_  (.D(_0165_),
    .CK(clknet_4_13_0_clk),
    .Q(\input_buffer[4][14] ),
    .QN(_1429_));
 DFF_X1 \input_buffer[4][15]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_4_12_0_clk),
    .Q(\input_buffer[4][15] ),
    .QN(_1428_));
 DFF_X1 \input_buffer[4][16]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][16] ),
    .QN(_1427_));
 DFF_X1 \input_buffer[4][17]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][17] ),
    .QN(_1426_));
 DFF_X1 \input_buffer[4][18]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][18] ),
    .QN(_1425_));
 DFF_X1 \input_buffer[4][19]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][19] ),
    .QN(_1424_));
 DFF_X1 \input_buffer[4][1]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][1] ),
    .QN(_1423_));
 DFF_X1 \input_buffer[4][20]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_4_15_0_clk),
    .Q(\input_buffer[4][20] ),
    .QN(_1422_));
 DFF_X1 \input_buffer[4][21]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[4][21] ),
    .QN(_1421_));
 DFF_X1 \input_buffer[4][22]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[4][22] ),
    .QN(_1420_));
 DFF_X1 \input_buffer[4][23]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_4_14_0_clk),
    .Q(\input_buffer[4][23] ),
    .QN(_1419_));
 DFF_X1 \input_buffer[4][24]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[4][0] ),
    .QN(_1418_));
 DFF_X1 \input_buffer[4][25]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[4][1] ),
    .QN(_1417_));
 DFF_X1 \input_buffer[4][26]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[4][2] ),
    .QN(_1416_));
 DFF_X1 \input_buffer[4][27]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_4_11_0_clk),
    .Q(\dest_id[4][3] ),
    .QN(_1415_));
 DFF_X1 \input_buffer[4][28]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[4][4] ),
    .QN(_1414_));
 DFF_X1 \input_buffer[4][29]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[4][5] ),
    .QN(_1413_));
 DFF_X1 \input_buffer[4][2]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][2] ),
    .QN(_1412_));
 DFF_X1 \input_buffer[4][30]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[4][6] ),
    .QN(_1411_));
 DFF_X1 \input_buffer[4][31]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_4_8_0_clk),
    .Q(\dest_id[4][7] ),
    .QN(_1410_));
 DFF_X1 \input_buffer[4][3]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][3] ),
    .QN(_1409_));
 DFF_X1 \input_buffer[4][4]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][4] ),
    .QN(_1408_));
 DFF_X1 \input_buffer[4][5]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][5] ),
    .QN(_1407_));
 DFF_X1 \input_buffer[4][6]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][6] ),
    .QN(_1406_));
 DFF_X1 \input_buffer[4][7]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][7] ),
    .QN(_1405_));
 DFF_X1 \input_buffer[4][8]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_4_11_0_clk),
    .Q(\input_buffer[4][8] ),
    .QN(_1404_));
 DFF_X1 \input_buffer[4][9]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_4_10_0_clk),
    .Q(\input_buffer[4][9] ),
    .QN(_1403_));
 DFF_X1 \input_buffer_valid[0]$_SDFF_PN0_  (.D(_0192_),
    .CK(clknet_4_1_0_clk),
    .Q(\input_buffer_valid[0] ),
    .QN(net237));
 DFF_X1 \input_buffer_valid[1]$_SDFF_PN0_  (.D(_0193_),
    .CK(clknet_4_3_0_clk),
    .Q(\input_buffer_valid[1] ),
    .QN(net169));
 DFF_X1 \input_buffer_valid[2]$_SDFF_PN0_  (.D(_0194_),
    .CK(clknet_4_2_0_clk),
    .Q(\input_buffer_valid[2] ),
    .QN(net271));
 DFF_X1 \input_buffer_valid[3]$_SDFF_PN0_  (.D(_0195_),
    .CK(clknet_4_2_0_clk),
    .Q(\input_buffer_valid[3] ),
    .QN(net305));
 DFF_X1 \input_buffer_valid[4]$_SDFF_PN0_  (.D(_0196_),
    .CK(clknet_4_2_0_clk),
    .Q(\input_buffer_valid[4] ),
    .QN(net203));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_103 ();
 BUF_X1 input1 (.A(east_in_data[0]),
    .Z(net1));
 BUF_X1 input2 (.A(east_in_data[10]),
    .Z(net2));
 BUF_X1 input3 (.A(east_in_data[11]),
    .Z(net3));
 BUF_X1 input4 (.A(east_in_data[12]),
    .Z(net4));
 BUF_X1 input5 (.A(east_in_data[13]),
    .Z(net5));
 BUF_X1 input6 (.A(east_in_data[14]),
    .Z(net6));
 BUF_X1 input7 (.A(east_in_data[15]),
    .Z(net7));
 BUF_X1 input8 (.A(east_in_data[16]),
    .Z(net8));
 BUF_X1 input9 (.A(east_in_data[17]),
    .Z(net9));
 BUF_X1 input10 (.A(east_in_data[18]),
    .Z(net10));
 BUF_X1 input11 (.A(east_in_data[19]),
    .Z(net11));
 BUF_X1 input12 (.A(east_in_data[1]),
    .Z(net12));
 BUF_X1 input13 (.A(east_in_data[20]),
    .Z(net13));
 BUF_X1 input14 (.A(east_in_data[21]),
    .Z(net14));
 BUF_X1 input15 (.A(east_in_data[22]),
    .Z(net15));
 BUF_X1 input16 (.A(east_in_data[23]),
    .Z(net16));
 BUF_X1 input17 (.A(east_in_data[24]),
    .Z(net17));
 BUF_X1 input18 (.A(east_in_data[25]),
    .Z(net18));
 BUF_X1 input19 (.A(east_in_data[26]),
    .Z(net19));
 BUF_X1 input20 (.A(east_in_data[27]),
    .Z(net20));
 BUF_X1 input21 (.A(east_in_data[28]),
    .Z(net21));
 BUF_X1 input22 (.A(east_in_data[29]),
    .Z(net22));
 BUF_X1 input23 (.A(east_in_data[2]),
    .Z(net23));
 BUF_X1 input24 (.A(east_in_data[30]),
    .Z(net24));
 BUF_X1 input25 (.A(east_in_data[31]),
    .Z(net25));
 BUF_X1 input26 (.A(east_in_data[3]),
    .Z(net26));
 BUF_X1 input27 (.A(east_in_data[4]),
    .Z(net27));
 BUF_X1 input28 (.A(east_in_data[5]),
    .Z(net28));
 BUF_X1 input29 (.A(east_in_data[6]),
    .Z(net29));
 BUF_X1 input30 (.A(east_in_data[7]),
    .Z(net30));
 BUF_X1 input31 (.A(east_in_data[8]),
    .Z(net31));
 BUF_X1 input32 (.A(east_in_data[9]),
    .Z(net32));
 BUF_X1 input33 (.A(east_in_valid),
    .Z(net33));
 BUF_X1 input34 (.A(east_out_ready),
    .Z(net34));
 BUF_X1 input35 (.A(local_in_data[0]),
    .Z(net35));
 BUF_X1 input36 (.A(local_in_data[10]),
    .Z(net36));
 BUF_X1 input37 (.A(local_in_data[11]),
    .Z(net37));
 BUF_X1 input38 (.A(local_in_data[12]),
    .Z(net38));
 BUF_X1 input39 (.A(local_in_data[13]),
    .Z(net39));
 BUF_X1 input40 (.A(local_in_data[14]),
    .Z(net40));
 BUF_X1 input41 (.A(local_in_data[15]),
    .Z(net41));
 BUF_X1 input42 (.A(local_in_data[16]),
    .Z(net42));
 BUF_X1 input43 (.A(local_in_data[17]),
    .Z(net43));
 BUF_X1 input44 (.A(local_in_data[18]),
    .Z(net44));
 BUF_X1 input45 (.A(local_in_data[19]),
    .Z(net45));
 BUF_X1 input46 (.A(local_in_data[1]),
    .Z(net46));
 BUF_X1 input47 (.A(local_in_data[20]),
    .Z(net47));
 BUF_X1 input48 (.A(local_in_data[21]),
    .Z(net48));
 BUF_X1 input49 (.A(local_in_data[22]),
    .Z(net49));
 BUF_X1 input50 (.A(local_in_data[23]),
    .Z(net50));
 BUF_X1 input51 (.A(local_in_data[24]),
    .Z(net51));
 BUF_X1 input52 (.A(local_in_data[25]),
    .Z(net52));
 BUF_X1 input53 (.A(local_in_data[26]),
    .Z(net53));
 BUF_X1 input54 (.A(local_in_data[27]),
    .Z(net54));
 BUF_X1 input55 (.A(local_in_data[28]),
    .Z(net55));
 BUF_X1 input56 (.A(local_in_data[29]),
    .Z(net56));
 BUF_X1 input57 (.A(local_in_data[2]),
    .Z(net57));
 BUF_X1 input58 (.A(local_in_data[30]),
    .Z(net58));
 BUF_X1 input59 (.A(local_in_data[31]),
    .Z(net59));
 BUF_X1 input60 (.A(local_in_data[3]),
    .Z(net60));
 BUF_X1 input61 (.A(local_in_data[4]),
    .Z(net61));
 BUF_X1 input62 (.A(local_in_data[5]),
    .Z(net62));
 BUF_X1 input63 (.A(local_in_data[6]),
    .Z(net63));
 BUF_X1 input64 (.A(local_in_data[7]),
    .Z(net64));
 BUF_X1 input65 (.A(local_in_data[8]),
    .Z(net65));
 BUF_X1 input66 (.A(local_in_data[9]),
    .Z(net66));
 BUF_X1 input67 (.A(local_in_valid),
    .Z(net67));
 BUF_X1 input68 (.A(north_in_data[0]),
    .Z(net68));
 BUF_X1 input69 (.A(north_in_data[10]),
    .Z(net69));
 BUF_X1 input70 (.A(north_in_data[11]),
    .Z(net70));
 BUF_X1 input71 (.A(north_in_data[12]),
    .Z(net71));
 BUF_X1 input72 (.A(north_in_data[13]),
    .Z(net72));
 BUF_X1 input73 (.A(north_in_data[14]),
    .Z(net73));
 BUF_X1 input74 (.A(north_in_data[15]),
    .Z(net74));
 BUF_X1 input75 (.A(north_in_data[16]),
    .Z(net75));
 BUF_X1 input76 (.A(north_in_data[17]),
    .Z(net76));
 BUF_X1 input77 (.A(north_in_data[18]),
    .Z(net77));
 BUF_X1 input78 (.A(north_in_data[19]),
    .Z(net78));
 BUF_X1 input79 (.A(north_in_data[1]),
    .Z(net79));
 BUF_X1 input80 (.A(north_in_data[20]),
    .Z(net80));
 BUF_X1 input81 (.A(north_in_data[21]),
    .Z(net81));
 BUF_X1 input82 (.A(north_in_data[22]),
    .Z(net82));
 BUF_X1 input83 (.A(north_in_data[23]),
    .Z(net83));
 BUF_X1 input84 (.A(north_in_data[24]),
    .Z(net84));
 BUF_X1 input85 (.A(north_in_data[25]),
    .Z(net85));
 BUF_X1 input86 (.A(north_in_data[26]),
    .Z(net86));
 BUF_X1 input87 (.A(north_in_data[27]),
    .Z(net87));
 BUF_X1 input88 (.A(north_in_data[28]),
    .Z(net88));
 BUF_X1 input89 (.A(north_in_data[29]),
    .Z(net89));
 BUF_X1 input90 (.A(north_in_data[2]),
    .Z(net90));
 BUF_X1 input91 (.A(north_in_data[30]),
    .Z(net91));
 BUF_X1 input92 (.A(north_in_data[31]),
    .Z(net92));
 BUF_X1 input93 (.A(north_in_data[3]),
    .Z(net93));
 BUF_X1 input94 (.A(north_in_data[4]),
    .Z(net94));
 BUF_X1 input95 (.A(north_in_data[5]),
    .Z(net95));
 BUF_X1 input96 (.A(north_in_data[6]),
    .Z(net96));
 BUF_X1 input97 (.A(north_in_data[7]),
    .Z(net97));
 BUF_X1 input98 (.A(north_in_data[8]),
    .Z(net98));
 BUF_X1 input99 (.A(north_in_data[9]),
    .Z(net99));
 BUF_X1 input100 (.A(north_in_valid),
    .Z(net100));
 BUF_X1 input101 (.A(south_in_data[0]),
    .Z(net101));
 BUF_X1 input102 (.A(south_in_data[10]),
    .Z(net102));
 BUF_X1 input103 (.A(south_in_data[11]),
    .Z(net103));
 BUF_X1 input104 (.A(south_in_data[12]),
    .Z(net104));
 BUF_X1 input105 (.A(south_in_data[13]),
    .Z(net105));
 BUF_X1 input106 (.A(south_in_data[14]),
    .Z(net106));
 BUF_X1 input107 (.A(south_in_data[15]),
    .Z(net107));
 BUF_X1 input108 (.A(south_in_data[16]),
    .Z(net108));
 BUF_X1 input109 (.A(south_in_data[17]),
    .Z(net109));
 BUF_X1 input110 (.A(south_in_data[18]),
    .Z(net110));
 BUF_X1 input111 (.A(south_in_data[19]),
    .Z(net111));
 BUF_X1 input112 (.A(south_in_data[1]),
    .Z(net112));
 BUF_X1 input113 (.A(south_in_data[20]),
    .Z(net113));
 BUF_X1 input114 (.A(south_in_data[21]),
    .Z(net114));
 BUF_X1 input115 (.A(south_in_data[22]),
    .Z(net115));
 BUF_X1 input116 (.A(south_in_data[23]),
    .Z(net116));
 BUF_X1 input117 (.A(south_in_data[24]),
    .Z(net117));
 BUF_X1 input118 (.A(south_in_data[25]),
    .Z(net118));
 BUF_X1 input119 (.A(south_in_data[26]),
    .Z(net119));
 BUF_X1 input120 (.A(south_in_data[27]),
    .Z(net120));
 BUF_X1 input121 (.A(south_in_data[28]),
    .Z(net121));
 BUF_X1 input122 (.A(south_in_data[29]),
    .Z(net122));
 BUF_X1 input123 (.A(south_in_data[2]),
    .Z(net123));
 BUF_X1 input124 (.A(south_in_data[30]),
    .Z(net124));
 BUF_X1 input125 (.A(south_in_data[31]),
    .Z(net125));
 BUF_X1 input126 (.A(south_in_data[3]),
    .Z(net126));
 BUF_X1 input127 (.A(south_in_data[4]),
    .Z(net127));
 BUF_X1 input128 (.A(south_in_data[5]),
    .Z(net128));
 BUF_X1 input129 (.A(south_in_data[6]),
    .Z(net129));
 BUF_X1 input130 (.A(south_in_data[7]),
    .Z(net130));
 BUF_X1 input131 (.A(south_in_data[8]),
    .Z(net131));
 BUF_X1 input132 (.A(south_in_data[9]),
    .Z(net132));
 BUF_X1 input133 (.A(south_in_valid),
    .Z(net133));
 BUF_X1 input134 (.A(south_out_ready),
    .Z(net134));
 BUF_X1 input135 (.A(west_in_data[0]),
    .Z(net135));
 BUF_X1 input136 (.A(west_in_data[10]),
    .Z(net136));
 BUF_X1 input137 (.A(west_in_data[11]),
    .Z(net137));
 BUF_X1 input138 (.A(west_in_data[12]),
    .Z(net138));
 BUF_X1 input139 (.A(west_in_data[13]),
    .Z(net139));
 BUF_X1 input140 (.A(west_in_data[14]),
    .Z(net140));
 BUF_X1 input141 (.A(west_in_data[15]),
    .Z(net141));
 BUF_X1 input142 (.A(west_in_data[16]),
    .Z(net142));
 BUF_X1 input143 (.A(west_in_data[17]),
    .Z(net143));
 BUF_X1 input144 (.A(west_in_data[18]),
    .Z(net144));
 BUF_X1 input145 (.A(west_in_data[19]),
    .Z(net145));
 BUF_X1 input146 (.A(west_in_data[1]),
    .Z(net146));
 BUF_X1 input147 (.A(west_in_data[20]),
    .Z(net147));
 BUF_X1 input148 (.A(west_in_data[21]),
    .Z(net148));
 BUF_X1 input149 (.A(west_in_data[22]),
    .Z(net149));
 BUF_X1 input150 (.A(west_in_data[23]),
    .Z(net150));
 BUF_X1 input151 (.A(west_in_data[24]),
    .Z(net151));
 BUF_X1 input152 (.A(west_in_data[25]),
    .Z(net152));
 BUF_X1 input153 (.A(west_in_data[26]),
    .Z(net153));
 BUF_X1 input154 (.A(west_in_data[27]),
    .Z(net154));
 BUF_X1 input155 (.A(west_in_data[28]),
    .Z(net155));
 BUF_X1 input156 (.A(west_in_data[29]),
    .Z(net156));
 BUF_X1 input157 (.A(west_in_data[2]),
    .Z(net157));
 BUF_X1 input158 (.A(west_in_data[30]),
    .Z(net158));
 BUF_X1 input159 (.A(west_in_data[31]),
    .Z(net159));
 BUF_X1 input160 (.A(west_in_data[3]),
    .Z(net160));
 BUF_X1 input161 (.A(west_in_data[4]),
    .Z(net161));
 BUF_X1 input162 (.A(west_in_data[5]),
    .Z(net162));
 BUF_X1 input163 (.A(west_in_data[6]),
    .Z(net163));
 BUF_X1 input164 (.A(west_in_data[7]),
    .Z(net164));
 BUF_X1 input165 (.A(west_in_data[8]),
    .Z(net165));
 BUF_X1 input166 (.A(west_in_data[9]),
    .Z(net166));
 CLKBUF_X2 input167 (.A(west_in_valid),
    .Z(net167));
 BUF_X1 input168 (.A(west_out_ready),
    .Z(net168));
 BUF_X1 output169 (.A(net169),
    .Z(east_in_ready));
 BUF_X1 output170 (.A(net170),
    .Z(east_out_data[0]));
 BUF_X1 output171 (.A(net171),
    .Z(east_out_data[10]));
 BUF_X1 output172 (.A(net172),
    .Z(east_out_data[11]));
 BUF_X1 output173 (.A(net173),
    .Z(east_out_data[12]));
 BUF_X1 output174 (.A(net174),
    .Z(east_out_data[13]));
 BUF_X1 output175 (.A(net175),
    .Z(east_out_data[14]));
 BUF_X1 output176 (.A(net176),
    .Z(east_out_data[15]));
 BUF_X1 output177 (.A(net177),
    .Z(east_out_data[16]));
 BUF_X1 output178 (.A(net178),
    .Z(east_out_data[17]));
 BUF_X1 output179 (.A(net179),
    .Z(east_out_data[18]));
 BUF_X1 output180 (.A(net180),
    .Z(east_out_data[19]));
 BUF_X1 output181 (.A(net181),
    .Z(east_out_data[1]));
 BUF_X1 output182 (.A(net182),
    .Z(east_out_data[20]));
 BUF_X1 output183 (.A(net183),
    .Z(east_out_data[21]));
 BUF_X1 output184 (.A(net184),
    .Z(east_out_data[22]));
 BUF_X1 output185 (.A(net185),
    .Z(east_out_data[23]));
 BUF_X1 output186 (.A(net186),
    .Z(east_out_data[24]));
 BUF_X1 output187 (.A(net187),
    .Z(east_out_data[25]));
 BUF_X1 output188 (.A(net188),
    .Z(east_out_data[26]));
 BUF_X1 output189 (.A(net189),
    .Z(east_out_data[27]));
 BUF_X1 output190 (.A(net190),
    .Z(east_out_data[28]));
 BUF_X1 output191 (.A(net191),
    .Z(east_out_data[29]));
 BUF_X1 output192 (.A(net192),
    .Z(east_out_data[2]));
 BUF_X1 output193 (.A(net193),
    .Z(east_out_data[30]));
 BUF_X1 output194 (.A(net194),
    .Z(east_out_data[31]));
 BUF_X1 output195 (.A(net195),
    .Z(east_out_data[3]));
 BUF_X1 output196 (.A(net196),
    .Z(east_out_data[4]));
 BUF_X1 output197 (.A(net197),
    .Z(east_out_data[5]));
 BUF_X1 output198 (.A(net198),
    .Z(east_out_data[6]));
 BUF_X1 output199 (.A(net199),
    .Z(east_out_data[7]));
 BUF_X1 output200 (.A(net200),
    .Z(east_out_data[8]));
 BUF_X1 output201 (.A(net201),
    .Z(east_out_data[9]));
 BUF_X1 output202 (.A(net202),
    .Z(east_out_valid));
 BUF_X1 output203 (.A(net203),
    .Z(local_in_ready));
 BUF_X1 output204 (.A(net204),
    .Z(local_out_data[0]));
 BUF_X1 output205 (.A(net205),
    .Z(local_out_data[10]));
 BUF_X1 output206 (.A(net206),
    .Z(local_out_data[11]));
 BUF_X1 output207 (.A(net207),
    .Z(local_out_data[12]));
 BUF_X1 output208 (.A(net208),
    .Z(local_out_data[13]));
 BUF_X1 output209 (.A(net209),
    .Z(local_out_data[14]));
 BUF_X1 output210 (.A(net210),
    .Z(local_out_data[15]));
 BUF_X1 output211 (.A(net211),
    .Z(local_out_data[16]));
 BUF_X1 output212 (.A(net212),
    .Z(local_out_data[17]));
 BUF_X1 output213 (.A(net213),
    .Z(local_out_data[18]));
 BUF_X1 output214 (.A(net214),
    .Z(local_out_data[19]));
 BUF_X1 output215 (.A(net215),
    .Z(local_out_data[1]));
 BUF_X1 output216 (.A(net216),
    .Z(local_out_data[20]));
 BUF_X1 output217 (.A(net217),
    .Z(local_out_data[21]));
 BUF_X1 output218 (.A(net218),
    .Z(local_out_data[22]));
 BUF_X1 output219 (.A(net219),
    .Z(local_out_data[23]));
 BUF_X1 output220 (.A(net220),
    .Z(local_out_data[24]));
 BUF_X1 output221 (.A(net221),
    .Z(local_out_data[25]));
 BUF_X1 output222 (.A(net222),
    .Z(local_out_data[26]));
 BUF_X1 output223 (.A(net223),
    .Z(local_out_data[27]));
 BUF_X1 output224 (.A(net224),
    .Z(local_out_data[28]));
 BUF_X1 output225 (.A(net225),
    .Z(local_out_data[29]));
 BUF_X1 output226 (.A(net226),
    .Z(local_out_data[2]));
 BUF_X1 output227 (.A(net227),
    .Z(local_out_data[30]));
 BUF_X1 output228 (.A(net228),
    .Z(local_out_data[31]));
 BUF_X1 output229 (.A(net229),
    .Z(local_out_data[3]));
 BUF_X1 output230 (.A(net230),
    .Z(local_out_data[4]));
 BUF_X1 output231 (.A(net231),
    .Z(local_out_data[5]));
 BUF_X1 output232 (.A(net232),
    .Z(local_out_data[6]));
 BUF_X1 output233 (.A(net233),
    .Z(local_out_data[7]));
 BUF_X1 output234 (.A(net234),
    .Z(local_out_data[8]));
 BUF_X1 output235 (.A(net235),
    .Z(local_out_data[9]));
 BUF_X1 output236 (.A(net236),
    .Z(local_out_valid));
 BUF_X1 output237 (.A(net237),
    .Z(north_in_ready));
 BUF_X1 output238 (.A(net238),
    .Z(north_out_data[0]));
 BUF_X1 output239 (.A(net239),
    .Z(north_out_data[10]));
 BUF_X1 output240 (.A(net240),
    .Z(north_out_data[11]));
 BUF_X1 output241 (.A(net241),
    .Z(north_out_data[12]));
 BUF_X1 output242 (.A(net242),
    .Z(north_out_data[13]));
 BUF_X1 output243 (.A(net243),
    .Z(north_out_data[14]));
 BUF_X1 output244 (.A(net244),
    .Z(north_out_data[15]));
 BUF_X1 output245 (.A(net245),
    .Z(north_out_data[16]));
 BUF_X1 output246 (.A(net246),
    .Z(north_out_data[17]));
 BUF_X1 output247 (.A(net247),
    .Z(north_out_data[18]));
 BUF_X1 output248 (.A(net248),
    .Z(north_out_data[19]));
 BUF_X1 output249 (.A(net249),
    .Z(north_out_data[1]));
 BUF_X1 output250 (.A(net250),
    .Z(north_out_data[20]));
 BUF_X1 output251 (.A(net251),
    .Z(north_out_data[21]));
 BUF_X1 output252 (.A(net252),
    .Z(north_out_data[22]));
 BUF_X1 output253 (.A(net253),
    .Z(north_out_data[23]));
 BUF_X1 output254 (.A(net254),
    .Z(north_out_data[24]));
 BUF_X1 output255 (.A(net255),
    .Z(north_out_data[25]));
 BUF_X1 output256 (.A(net256),
    .Z(north_out_data[26]));
 BUF_X1 output257 (.A(net257),
    .Z(north_out_data[27]));
 BUF_X1 output258 (.A(net258),
    .Z(north_out_data[28]));
 BUF_X1 output259 (.A(net259),
    .Z(north_out_data[29]));
 BUF_X1 output260 (.A(net260),
    .Z(north_out_data[2]));
 BUF_X1 output261 (.A(net261),
    .Z(north_out_data[30]));
 BUF_X1 output262 (.A(net262),
    .Z(north_out_data[31]));
 BUF_X1 output263 (.A(net263),
    .Z(north_out_data[3]));
 BUF_X1 output264 (.A(net264),
    .Z(north_out_data[4]));
 BUF_X1 output265 (.A(net265),
    .Z(north_out_data[5]));
 BUF_X1 output266 (.A(net266),
    .Z(north_out_data[6]));
 BUF_X1 output267 (.A(net267),
    .Z(north_out_data[7]));
 BUF_X1 output268 (.A(net268),
    .Z(north_out_data[8]));
 BUF_X1 output269 (.A(net269),
    .Z(north_out_data[9]));
 BUF_X1 output270 (.A(net270),
    .Z(north_out_valid));
 BUF_X1 output271 (.A(net271),
    .Z(south_in_ready));
 BUF_X1 output272 (.A(net272),
    .Z(south_out_data[0]));
 BUF_X1 output273 (.A(net273),
    .Z(south_out_data[10]));
 BUF_X1 output274 (.A(net274),
    .Z(south_out_data[11]));
 BUF_X1 output275 (.A(net275),
    .Z(south_out_data[12]));
 BUF_X1 output276 (.A(net276),
    .Z(south_out_data[13]));
 BUF_X1 output277 (.A(net277),
    .Z(south_out_data[14]));
 BUF_X1 output278 (.A(net278),
    .Z(south_out_data[15]));
 BUF_X1 output279 (.A(net279),
    .Z(south_out_data[16]));
 BUF_X1 output280 (.A(net280),
    .Z(south_out_data[17]));
 BUF_X1 output281 (.A(net281),
    .Z(south_out_data[18]));
 BUF_X1 output282 (.A(net282),
    .Z(south_out_data[19]));
 BUF_X1 output283 (.A(net283),
    .Z(south_out_data[1]));
 BUF_X1 output284 (.A(net284),
    .Z(south_out_data[20]));
 BUF_X1 output285 (.A(net285),
    .Z(south_out_data[21]));
 BUF_X1 output286 (.A(net286),
    .Z(south_out_data[22]));
 BUF_X1 output287 (.A(net287),
    .Z(south_out_data[23]));
 BUF_X1 output288 (.A(net288),
    .Z(south_out_data[24]));
 BUF_X1 output289 (.A(net289),
    .Z(south_out_data[25]));
 BUF_X1 output290 (.A(net290),
    .Z(south_out_data[26]));
 BUF_X1 output291 (.A(net291),
    .Z(south_out_data[27]));
 BUF_X1 output292 (.A(net292),
    .Z(south_out_data[28]));
 BUF_X1 output293 (.A(net293),
    .Z(south_out_data[29]));
 BUF_X1 output294 (.A(net294),
    .Z(south_out_data[2]));
 BUF_X1 output295 (.A(net295),
    .Z(south_out_data[30]));
 BUF_X1 output296 (.A(net296),
    .Z(south_out_data[31]));
 BUF_X1 output297 (.A(net297),
    .Z(south_out_data[3]));
 BUF_X1 output298 (.A(net298),
    .Z(south_out_data[4]));
 BUF_X1 output299 (.A(net299),
    .Z(south_out_data[5]));
 BUF_X1 output300 (.A(net300),
    .Z(south_out_data[6]));
 BUF_X1 output301 (.A(net301),
    .Z(south_out_data[7]));
 BUF_X1 output302 (.A(net302),
    .Z(south_out_data[8]));
 BUF_X1 output303 (.A(net303),
    .Z(south_out_data[9]));
 BUF_X1 output304 (.A(net304),
    .Z(south_out_valid));
 BUF_X1 output305 (.A(net305),
    .Z(west_in_ready));
 BUF_X1 output306 (.A(net306),
    .Z(west_out_data[0]));
 BUF_X1 output307 (.A(net307),
    .Z(west_out_data[10]));
 BUF_X1 output308 (.A(net308),
    .Z(west_out_data[11]));
 BUF_X1 output309 (.A(net309),
    .Z(west_out_data[12]));
 BUF_X1 output310 (.A(net310),
    .Z(west_out_data[13]));
 BUF_X1 output311 (.A(net311),
    .Z(west_out_data[14]));
 BUF_X1 output312 (.A(net312),
    .Z(west_out_data[15]));
 BUF_X1 output313 (.A(net313),
    .Z(west_out_data[16]));
 BUF_X1 output314 (.A(net314),
    .Z(west_out_data[17]));
 BUF_X1 output315 (.A(net315),
    .Z(west_out_data[18]));
 BUF_X1 output316 (.A(net316),
    .Z(west_out_data[19]));
 BUF_X1 output317 (.A(net317),
    .Z(west_out_data[1]));
 BUF_X1 output318 (.A(net318),
    .Z(west_out_data[20]));
 BUF_X1 output319 (.A(net319),
    .Z(west_out_data[21]));
 BUF_X1 output320 (.A(net320),
    .Z(west_out_data[22]));
 BUF_X1 output321 (.A(net321),
    .Z(west_out_data[23]));
 BUF_X1 output322 (.A(net322),
    .Z(west_out_data[24]));
 BUF_X1 output323 (.A(net323),
    .Z(west_out_data[25]));
 BUF_X1 output324 (.A(net324),
    .Z(west_out_data[26]));
 BUF_X1 output325 (.A(net325),
    .Z(west_out_data[27]));
 BUF_X1 output326 (.A(net326),
    .Z(west_out_data[28]));
 BUF_X1 output327 (.A(net327),
    .Z(west_out_data[29]));
 BUF_X1 output328 (.A(net328),
    .Z(west_out_data[2]));
 BUF_X1 output329 (.A(net329),
    .Z(west_out_data[30]));
 BUF_X1 output330 (.A(net330),
    .Z(west_out_data[31]));
 BUF_X1 output331 (.A(net331),
    .Z(west_out_data[3]));
 BUF_X1 output332 (.A(net332),
    .Z(west_out_data[4]));
 BUF_X1 output333 (.A(net333),
    .Z(west_out_data[5]));
 BUF_X1 output334 (.A(net334),
    .Z(west_out_data[6]));
 BUF_X1 output335 (.A(net335),
    .Z(west_out_data[7]));
 BUF_X1 output336 (.A(net336),
    .Z(west_out_data[8]));
 BUF_X1 output337 (.A(net337),
    .Z(west_out_data[9]));
 BUF_X1 output338 (.A(net338),
    .Z(west_out_valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X2 clkload0 (.A(clknet_4_0_0_clk));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk));
 INV_X4 clkload2 (.A(clknet_4_2_0_clk));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk));
 INV_X4 clkload4 (.A(clknet_4_4_0_clk));
 INV_X2 clkload5 (.A(clknet_4_5_0_clk));
 INV_X2 clkload6 (.A(clknet_4_6_0_clk));
 INV_X2 clkload7 (.A(clknet_4_8_0_clk));
 INV_X4 clkload8 (.A(clknet_4_9_0_clk));
 INV_X2 clkload9 (.A(clknet_4_10_0_clk));
 INV_X1 clkload10 (.A(clknet_4_11_0_clk));
 INV_X4 clkload11 (.A(clknet_4_12_0_clk));
 INV_X4 clkload12 (.A(clknet_4_13_0_clk));
 INV_X2 clkload13 (.A(clknet_4_14_0_clk));
 INV_X2 clkload14 (.A(clknet_4_15_0_clk));
 BUF_X1 rebuffer1 (.A(_1332_),
    .Z(net339));
 BUF_X1 rebuffer2 (.A(_1332_),
    .Z(net340));
 BUF_X1 rebuffer3 (.A(net340),
    .Z(net341));
 BUF_X1 rebuffer4 (.A(_1332_),
    .Z(net342));
 BUF_X1 rebuffer6 (.A(net343),
    .Z(net344));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_33 ();
 FILLCELL_X2 FILLER_0_37 ();
 FILLCELL_X16 FILLER_0_42 ();
 FILLCELL_X4 FILLER_0_58 ();
 FILLCELL_X2 FILLER_0_68 ();
 FILLCELL_X1 FILLER_0_70 ();
 FILLCELL_X8 FILLER_0_74 ();
 FILLCELL_X4 FILLER_0_88 ();
 FILLCELL_X2 FILLER_0_92 ();
 FILLCELL_X1 FILLER_0_124 ();
 FILLCELL_X1 FILLER_0_134 ();
 FILLCELL_X1 FILLER_0_148 ();
 FILLCELL_X1 FILLER_0_221 ();
 FILLCELL_X4 FILLER_0_245 ();
 FILLCELL_X1 FILLER_0_249 ();
 FILLCELL_X4 FILLER_0_253 ();
 FILLCELL_X4 FILLER_0_263 ();
 FILLCELL_X2 FILLER_0_267 ();
 FILLCELL_X1 FILLER_0_276 ();
 FILLCELL_X1 FILLER_0_283 ();
 FILLCELL_X2 FILLER_0_294 ();
 FILLCELL_X1 FILLER_0_303 ();
 FILLCELL_X1 FILLER_0_317 ();
 FILLCELL_X1 FILLER_0_345 ();
 FILLCELL_X32 FILLER_0_349 ();
 FILLCELL_X4 FILLER_0_381 ();
 FILLCELL_X1 FILLER_0_385 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X16 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_81 ();
 FILLCELL_X4 FILLER_1_88 ();
 FILLCELL_X1 FILLER_1_217 ();
 FILLCELL_X2 FILLER_1_245 ();
 FILLCELL_X32 FILLER_1_350 ();
 FILLCELL_X4 FILLER_1_382 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_97 ();
 FILLCELL_X1 FILLER_2_101 ();
 FILLCELL_X16 FILLER_2_105 ();
 FILLCELL_X4 FILLER_2_121 ();
 FILLCELL_X2 FILLER_2_125 ();
 FILLCELL_X4 FILLER_2_155 ();
 FILLCELL_X2 FILLER_2_159 ();
 FILLCELL_X1 FILLER_2_161 ();
 FILLCELL_X2 FILLER_2_184 ();
 FILLCELL_X4 FILLER_2_192 ();
 FILLCELL_X2 FILLER_2_196 ();
 FILLCELL_X4 FILLER_2_202 ();
 FILLCELL_X2 FILLER_2_206 ();
 FILLCELL_X1 FILLER_2_208 ();
 FILLCELL_X2 FILLER_2_213 ();
 FILLCELL_X1 FILLER_2_215 ();
 FILLCELL_X8 FILLER_2_219 ();
 FILLCELL_X2 FILLER_2_227 ();
 FILLCELL_X8 FILLER_2_258 ();
 FILLCELL_X1 FILLER_2_266 ();
 FILLCELL_X4 FILLER_2_273 ();
 FILLCELL_X2 FILLER_2_277 ();
 FILLCELL_X1 FILLER_2_279 ();
 FILLCELL_X1 FILLER_2_286 ();
 FILLCELL_X8 FILLER_2_291 ();
 FILLCELL_X1 FILLER_2_303 ();
 FILLCELL_X32 FILLER_2_327 ();
 FILLCELL_X16 FILLER_2_359 ();
 FILLCELL_X8 FILLER_2_375 ();
 FILLCELL_X2 FILLER_2_383 ();
 FILLCELL_X1 FILLER_2_385 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_65 ();
 FILLCELL_X8 FILLER_3_73 ();
 FILLCELL_X4 FILLER_3_81 ();
 FILLCELL_X1 FILLER_3_85 ();
 FILLCELL_X16 FILLER_3_93 ();
 FILLCELL_X1 FILLER_3_109 ();
 FILLCELL_X4 FILLER_3_131 ();
 FILLCELL_X1 FILLER_3_135 ();
 FILLCELL_X4 FILLER_3_143 ();
 FILLCELL_X1 FILLER_3_147 ();
 FILLCELL_X2 FILLER_3_151 ();
 FILLCELL_X8 FILLER_3_157 ();
 FILLCELL_X8 FILLER_3_178 ();
 FILLCELL_X1 FILLER_3_186 ();
 FILLCELL_X1 FILLER_3_198 ();
 FILLCELL_X2 FILLER_3_202 ();
 FILLCELL_X4 FILLER_3_207 ();
 FILLCELL_X4 FILLER_3_214 ();
 FILLCELL_X1 FILLER_3_218 ();
 FILLCELL_X4 FILLER_3_225 ();
 FILLCELL_X1 FILLER_3_229 ();
 FILLCELL_X4 FILLER_3_237 ();
 FILLCELL_X1 FILLER_3_241 ();
 FILLCELL_X8 FILLER_3_262 ();
 FILLCELL_X2 FILLER_3_270 ();
 FILLCELL_X4 FILLER_3_275 ();
 FILLCELL_X2 FILLER_3_282 ();
 FILLCELL_X1 FILLER_3_284 ();
 FILLCELL_X2 FILLER_3_301 ();
 FILLCELL_X1 FILLER_3_303 ();
 FILLCELL_X4 FILLER_3_314 ();
 FILLCELL_X2 FILLER_3_318 ();
 FILLCELL_X1 FILLER_3_320 ();
 FILLCELL_X32 FILLER_3_328 ();
 FILLCELL_X16 FILLER_3_360 ();
 FILLCELL_X8 FILLER_3_376 ();
 FILLCELL_X2 FILLER_3_384 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_49 ();
 FILLCELL_X4 FILLER_4_57 ();
 FILLCELL_X2 FILLER_4_61 ();
 FILLCELL_X1 FILLER_4_63 ();
 FILLCELL_X2 FILLER_4_85 ();
 FILLCELL_X1 FILLER_4_87 ();
 FILLCELL_X16 FILLER_4_109 ();
 FILLCELL_X8 FILLER_4_125 ();
 FILLCELL_X2 FILLER_4_133 ();
 FILLCELL_X1 FILLER_4_135 ();
 FILLCELL_X1 FILLER_4_172 ();
 FILLCELL_X1 FILLER_4_186 ();
 FILLCELL_X1 FILLER_4_195 ();
 FILLCELL_X2 FILLER_4_207 ();
 FILLCELL_X1 FILLER_4_209 ();
 FILLCELL_X8 FILLER_4_217 ();
 FILLCELL_X1 FILLER_4_225 ();
 FILLCELL_X4 FILLER_4_243 ();
 FILLCELL_X2 FILLER_4_247 ();
 FILLCELL_X1 FILLER_4_249 ();
 FILLCELL_X2 FILLER_4_254 ();
 FILLCELL_X2 FILLER_4_264 ();
 FILLCELL_X1 FILLER_4_266 ();
 FILLCELL_X4 FILLER_4_270 ();
 FILLCELL_X1 FILLER_4_274 ();
 FILLCELL_X4 FILLER_4_282 ();
 FILLCELL_X2 FILLER_4_320 ();
 FILLCELL_X32 FILLER_4_343 ();
 FILLCELL_X8 FILLER_4_375 ();
 FILLCELL_X2 FILLER_4_383 ();
 FILLCELL_X1 FILLER_4_385 ();
 FILLCELL_X4 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_5 ();
 FILLCELL_X1 FILLER_5_7 ();
 FILLCELL_X16 FILLER_5_11 ();
 FILLCELL_X8 FILLER_5_27 ();
 FILLCELL_X4 FILLER_5_35 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_73 ();
 FILLCELL_X4 FILLER_5_81 ();
 FILLCELL_X2 FILLER_5_85 ();
 FILLCELL_X1 FILLER_5_87 ();
 FILLCELL_X16 FILLER_5_95 ();
 FILLCELL_X8 FILLER_5_111 ();
 FILLCELL_X4 FILLER_5_119 ();
 FILLCELL_X2 FILLER_5_125 ();
 FILLCELL_X1 FILLER_5_153 ();
 FILLCELL_X4 FILLER_5_177 ();
 FILLCELL_X1 FILLER_5_198 ();
 FILLCELL_X8 FILLER_5_203 ();
 FILLCELL_X4 FILLER_5_211 ();
 FILLCELL_X1 FILLER_5_215 ();
 FILLCELL_X16 FILLER_5_229 ();
 FILLCELL_X2 FILLER_5_245 ();
 FILLCELL_X1 FILLER_5_247 ();
 FILLCELL_X1 FILLER_5_261 ();
 FILLCELL_X2 FILLER_5_269 ();
 FILLCELL_X8 FILLER_5_292 ();
 FILLCELL_X2 FILLER_5_300 ();
 FILLCELL_X1 FILLER_5_306 ();
 FILLCELL_X4 FILLER_5_335 ();
 FILLCELL_X2 FILLER_5_339 ();
 FILLCELL_X16 FILLER_5_358 ();
 FILLCELL_X8 FILLER_5_374 ();
 FILLCELL_X4 FILLER_5_382 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_17 ();
 FILLCELL_X1 FILLER_6_21 ();
 FILLCELL_X4 FILLER_6_65 ();
 FILLCELL_X1 FILLER_6_69 ();
 FILLCELL_X2 FILLER_6_87 ();
 FILLCELL_X2 FILLER_6_114 ();
 FILLCELL_X1 FILLER_6_155 ();
 FILLCELL_X8 FILLER_6_210 ();
 FILLCELL_X4 FILLER_6_218 ();
 FILLCELL_X2 FILLER_6_222 ();
 FILLCELL_X4 FILLER_6_229 ();
 FILLCELL_X1 FILLER_6_233 ();
 FILLCELL_X8 FILLER_6_238 ();
 FILLCELL_X4 FILLER_6_267 ();
 FILLCELL_X1 FILLER_6_271 ();
 FILLCELL_X8 FILLER_6_279 ();
 FILLCELL_X2 FILLER_6_287 ();
 FILLCELL_X1 FILLER_6_289 ();
 FILLCELL_X8 FILLER_6_301 ();
 FILLCELL_X4 FILLER_6_309 ();
 FILLCELL_X8 FILLER_6_324 ();
 FILLCELL_X4 FILLER_6_332 ();
 FILLCELL_X2 FILLER_6_336 ();
 FILLCELL_X1 FILLER_6_338 ();
 FILLCELL_X8 FILLER_6_346 ();
 FILLCELL_X2 FILLER_6_354 ();
 FILLCELL_X16 FILLER_6_363 ();
 FILLCELL_X4 FILLER_6_379 ();
 FILLCELL_X2 FILLER_6_383 ();
 FILLCELL_X1 FILLER_6_385 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_5 ();
 FILLCELL_X1 FILLER_7_7 ();
 FILLCELL_X2 FILLER_7_14 ();
 FILLCELL_X1 FILLER_7_16 ();
 FILLCELL_X1 FILLER_7_43 ();
 FILLCELL_X2 FILLER_7_69 ();
 FILLCELL_X1 FILLER_7_71 ();
 FILLCELL_X2 FILLER_7_79 ();
 FILLCELL_X2 FILLER_7_120 ();
 FILLCELL_X1 FILLER_7_122 ();
 FILLCELL_X2 FILLER_7_147 ();
 FILLCELL_X1 FILLER_7_149 ();
 FILLCELL_X4 FILLER_7_157 ();
 FILLCELL_X2 FILLER_7_161 ();
 FILLCELL_X1 FILLER_7_163 ();
 FILLCELL_X2 FILLER_7_199 ();
 FILLCELL_X1 FILLER_7_201 ();
 FILLCELL_X8 FILLER_7_206 ();
 FILLCELL_X4 FILLER_7_214 ();
 FILLCELL_X2 FILLER_7_218 ();
 FILLCELL_X1 FILLER_7_220 ();
 FILLCELL_X2 FILLER_7_230 ();
 FILLCELL_X8 FILLER_7_261 ();
 FILLCELL_X4 FILLER_7_269 ();
 FILLCELL_X1 FILLER_7_273 ();
 FILLCELL_X1 FILLER_7_291 ();
 FILLCELL_X1 FILLER_7_309 ();
 FILLCELL_X32 FILLER_7_352 ();
 FILLCELL_X2 FILLER_7_384 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X16 FILLER_8_33 ();
 FILLCELL_X2 FILLER_8_49 ();
 FILLCELL_X1 FILLER_8_51 ();
 FILLCELL_X8 FILLER_8_58 ();
 FILLCELL_X2 FILLER_8_66 ();
 FILLCELL_X1 FILLER_8_68 ();
 FILLCELL_X2 FILLER_8_86 ();
 FILLCELL_X16 FILLER_8_95 ();
 FILLCELL_X4 FILLER_8_111 ();
 FILLCELL_X2 FILLER_8_115 ();
 FILLCELL_X8 FILLER_8_121 ();
 FILLCELL_X4 FILLER_8_129 ();
 FILLCELL_X1 FILLER_8_133 ();
 FILLCELL_X4 FILLER_8_138 ();
 FILLCELL_X4 FILLER_8_163 ();
 FILLCELL_X2 FILLER_8_167 ();
 FILLCELL_X1 FILLER_8_169 ();
 FILLCELL_X8 FILLER_8_190 ();
 FILLCELL_X4 FILLER_8_198 ();
 FILLCELL_X2 FILLER_8_202 ();
 FILLCELL_X1 FILLER_8_204 ();
 FILLCELL_X2 FILLER_8_208 ();
 FILLCELL_X2 FILLER_8_217 ();
 FILLCELL_X2 FILLER_8_224 ();
 FILLCELL_X2 FILLER_8_231 ();
 FILLCELL_X8 FILLER_8_242 ();
 FILLCELL_X1 FILLER_8_256 ();
 FILLCELL_X1 FILLER_8_261 ();
 FILLCELL_X16 FILLER_8_268 ();
 FILLCELL_X8 FILLER_8_284 ();
 FILLCELL_X1 FILLER_8_292 ();
 FILLCELL_X16 FILLER_8_302 ();
 FILLCELL_X8 FILLER_8_318 ();
 FILLCELL_X4 FILLER_8_326 ();
 FILLCELL_X2 FILLER_8_330 ();
 FILLCELL_X8 FILLER_8_339 ();
 FILLCELL_X4 FILLER_8_347 ();
 FILLCELL_X8 FILLER_8_372 ();
 FILLCELL_X2 FILLER_8_380 ();
 FILLCELL_X1 FILLER_8_382 ();
 FILLCELL_X4 FILLER_9_30 ();
 FILLCELL_X16 FILLER_9_41 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X8 FILLER_9_76 ();
 FILLCELL_X4 FILLER_9_84 ();
 FILLCELL_X2 FILLER_9_88 ();
 FILLCELL_X4 FILLER_9_107 ();
 FILLCELL_X1 FILLER_9_111 ();
 FILLCELL_X1 FILLER_9_136 ();
 FILLCELL_X4 FILLER_9_140 ();
 FILLCELL_X2 FILLER_9_144 ();
 FILLCELL_X2 FILLER_9_148 ();
 FILLCELL_X1 FILLER_9_150 ();
 FILLCELL_X2 FILLER_9_160 ();
 FILLCELL_X1 FILLER_9_162 ();
 FILLCELL_X16 FILLER_9_167 ();
 FILLCELL_X8 FILLER_9_183 ();
 FILLCELL_X4 FILLER_9_191 ();
 FILLCELL_X2 FILLER_9_195 ();
 FILLCELL_X2 FILLER_9_210 ();
 FILLCELL_X1 FILLER_9_217 ();
 FILLCELL_X4 FILLER_9_230 ();
 FILLCELL_X1 FILLER_9_236 ();
 FILLCELL_X1 FILLER_9_241 ();
 FILLCELL_X2 FILLER_9_254 ();
 FILLCELL_X16 FILLER_9_267 ();
 FILLCELL_X4 FILLER_9_283 ();
 FILLCELL_X2 FILLER_9_287 ();
 FILLCELL_X1 FILLER_9_289 ();
 FILLCELL_X8 FILLER_9_294 ();
 FILLCELL_X1 FILLER_9_302 ();
 FILLCELL_X16 FILLER_9_324 ();
 FILLCELL_X4 FILLER_9_340 ();
 FILLCELL_X1 FILLER_9_344 ();
 FILLCELL_X4 FILLER_9_359 ();
 FILLCELL_X2 FILLER_9_363 ();
 FILLCELL_X2 FILLER_9_368 ();
 FILLCELL_X2 FILLER_9_373 ();
 FILLCELL_X4 FILLER_9_381 ();
 FILLCELL_X1 FILLER_9_385 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X2 FILLER_10_5 ();
 FILLCELL_X1 FILLER_10_7 ();
 FILLCELL_X2 FILLER_10_11 ();
 FILLCELL_X1 FILLER_10_13 ();
 FILLCELL_X8 FILLER_10_17 ();
 FILLCELL_X4 FILLER_10_25 ();
 FILLCELL_X1 FILLER_10_29 ();
 FILLCELL_X8 FILLER_10_63 ();
 FILLCELL_X4 FILLER_10_71 ();
 FILLCELL_X16 FILLER_10_92 ();
 FILLCELL_X8 FILLER_10_108 ();
 FILLCELL_X2 FILLER_10_116 ();
 FILLCELL_X1 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_146 ();
 FILLCELL_X2 FILLER_10_160 ();
 FILLCELL_X1 FILLER_10_162 ();
 FILLCELL_X4 FILLER_10_183 ();
 FILLCELL_X2 FILLER_10_196 ();
 FILLCELL_X1 FILLER_10_200 ();
 FILLCELL_X1 FILLER_10_205 ();
 FILLCELL_X1 FILLER_10_211 ();
 FILLCELL_X4 FILLER_10_221 ();
 FILLCELL_X2 FILLER_10_225 ();
 FILLCELL_X4 FILLER_10_245 ();
 FILLCELL_X1 FILLER_10_249 ();
 FILLCELL_X1 FILLER_10_261 ();
 FILLCELL_X1 FILLER_10_268 ();
 FILLCELL_X1 FILLER_10_273 ();
 FILLCELL_X1 FILLER_10_287 ();
 FILLCELL_X8 FILLER_10_317 ();
 FILLCELL_X4 FILLER_10_325 ();
 FILLCELL_X2 FILLER_10_329 ();
 FILLCELL_X1 FILLER_10_331 ();
 FILLCELL_X4 FILLER_10_337 ();
 FILLCELL_X1 FILLER_10_341 ();
 FILLCELL_X4 FILLER_10_363 ();
 FILLCELL_X2 FILLER_10_367 ();
 FILLCELL_X8 FILLER_10_378 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_9 ();
 FILLCELL_X16 FILLER_11_42 ();
 FILLCELL_X2 FILLER_11_58 ();
 FILLCELL_X1 FILLER_11_60 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_80 ();
 FILLCELL_X4 FILLER_11_96 ();
 FILLCELL_X2 FILLER_11_100 ();
 FILLCELL_X1 FILLER_11_112 ();
 FILLCELL_X2 FILLER_11_116 ();
 FILLCELL_X4 FILLER_11_135 ();
 FILLCELL_X1 FILLER_11_184 ();
 FILLCELL_X1 FILLER_11_207 ();
 FILLCELL_X2 FILLER_11_214 ();
 FILLCELL_X1 FILLER_11_216 ();
 FILLCELL_X1 FILLER_11_225 ();
 FILLCELL_X2 FILLER_11_231 ();
 FILLCELL_X1 FILLER_11_253 ();
 FILLCELL_X2 FILLER_11_276 ();
 FILLCELL_X1 FILLER_11_293 ();
 FILLCELL_X2 FILLER_11_307 ();
 FILLCELL_X8 FILLER_11_323 ();
 FILLCELL_X1 FILLER_11_331 ();
 FILLCELL_X4 FILLER_11_349 ();
 FILLCELL_X2 FILLER_11_353 ();
 FILLCELL_X1 FILLER_11_355 ();
 FILLCELL_X16 FILLER_11_359 ();
 FILLCELL_X2 FILLER_11_375 ();
 FILLCELL_X1 FILLER_11_377 ();
 FILLCELL_X2 FILLER_11_384 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X2 FILLER_12_5 ();
 FILLCELL_X1 FILLER_12_7 ();
 FILLCELL_X16 FILLER_12_11 ();
 FILLCELL_X4 FILLER_12_27 ();
 FILLCELL_X16 FILLER_12_57 ();
 FILLCELL_X8 FILLER_12_73 ();
 FILLCELL_X4 FILLER_12_81 ();
 FILLCELL_X2 FILLER_12_85 ();
 FILLCELL_X1 FILLER_12_87 ();
 FILLCELL_X1 FILLER_12_92 ();
 FILLCELL_X1 FILLER_12_121 ();
 FILLCELL_X1 FILLER_12_173 ();
 FILLCELL_X1 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_190 ();
 FILLCELL_X1 FILLER_12_192 ();
 FILLCELL_X8 FILLER_12_200 ();
 FILLCELL_X4 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_212 ();
 FILLCELL_X2 FILLER_12_217 ();
 FILLCELL_X2 FILLER_12_225 ();
 FILLCELL_X1 FILLER_12_227 ();
 FILLCELL_X4 FILLER_12_242 ();
 FILLCELL_X2 FILLER_12_246 ();
 FILLCELL_X1 FILLER_12_270 ();
 FILLCELL_X2 FILLER_12_275 ();
 FILLCELL_X1 FILLER_12_277 ();
 FILLCELL_X4 FILLER_12_289 ();
 FILLCELL_X2 FILLER_12_293 ();
 FILLCELL_X1 FILLER_12_295 ();
 FILLCELL_X4 FILLER_12_304 ();
 FILLCELL_X8 FILLER_12_312 ();
 FILLCELL_X2 FILLER_12_320 ();
 FILLCELL_X4 FILLER_12_329 ();
 FILLCELL_X1 FILLER_12_333 ();
 FILLCELL_X2 FILLER_12_341 ();
 FILLCELL_X1 FILLER_12_343 ();
 FILLCELL_X4 FILLER_12_348 ();
 FILLCELL_X2 FILLER_12_352 ();
 FILLCELL_X4 FILLER_12_377 ();
 FILLCELL_X2 FILLER_12_381 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_3 ();
 FILLCELL_X8 FILLER_13_14 ();
 FILLCELL_X2 FILLER_13_22 ();
 FILLCELL_X8 FILLER_13_27 ();
 FILLCELL_X16 FILLER_13_38 ();
 FILLCELL_X1 FILLER_13_54 ();
 FILLCELL_X8 FILLER_13_81 ();
 FILLCELL_X2 FILLER_13_107 ();
 FILLCELL_X1 FILLER_13_109 ();
 FILLCELL_X2 FILLER_13_120 ();
 FILLCELL_X1 FILLER_13_129 ();
 FILLCELL_X2 FILLER_13_174 ();
 FILLCELL_X1 FILLER_13_196 ();
 FILLCELL_X8 FILLER_13_220 ();
 FILLCELL_X4 FILLER_13_257 ();
 FILLCELL_X2 FILLER_13_261 ();
 FILLCELL_X1 FILLER_13_263 ();
 FILLCELL_X1 FILLER_13_278 ();
 FILLCELL_X2 FILLER_13_298 ();
 FILLCELL_X1 FILLER_13_300 ();
 FILLCELL_X4 FILLER_13_314 ();
 FILLCELL_X1 FILLER_13_318 ();
 FILLCELL_X8 FILLER_13_340 ();
 FILLCELL_X4 FILLER_13_348 ();
 FILLCELL_X8 FILLER_13_359 ();
 FILLCELL_X1 FILLER_13_367 ();
 FILLCELL_X2 FILLER_13_372 ();
 FILLCELL_X1 FILLER_13_374 ();
 FILLCELL_X2 FILLER_13_378 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_25 ();
 FILLCELL_X2 FILLER_14_29 ();
 FILLCELL_X1 FILLER_14_31 ();
 FILLCELL_X1 FILLER_14_56 ();
 FILLCELL_X4 FILLER_14_62 ();
 FILLCELL_X1 FILLER_14_66 ();
 FILLCELL_X16 FILLER_14_74 ();
 FILLCELL_X1 FILLER_14_90 ();
 FILLCELL_X2 FILLER_14_93 ();
 FILLCELL_X1 FILLER_14_95 ();
 FILLCELL_X1 FILLER_14_100 ();
 FILLCELL_X2 FILLER_14_105 ();
 FILLCELL_X2 FILLER_14_111 ();
 FILLCELL_X1 FILLER_14_113 ();
 FILLCELL_X1 FILLER_14_190 ();
 FILLCELL_X4 FILLER_14_198 ();
 FILLCELL_X1 FILLER_14_202 ();
 FILLCELL_X8 FILLER_14_210 ();
 FILLCELL_X4 FILLER_14_218 ();
 FILLCELL_X2 FILLER_14_231 ();
 FILLCELL_X1 FILLER_14_233 ();
 FILLCELL_X2 FILLER_14_256 ();
 FILLCELL_X4 FILLER_14_284 ();
 FILLCELL_X2 FILLER_14_288 ();
 FILLCELL_X1 FILLER_14_290 ();
 FILLCELL_X2 FILLER_14_317 ();
 FILLCELL_X16 FILLER_14_322 ();
 FILLCELL_X8 FILLER_14_338 ();
 FILLCELL_X2 FILLER_14_349 ();
 FILLCELL_X1 FILLER_14_351 ();
 FILLCELL_X2 FILLER_14_363 ();
 FILLCELL_X1 FILLER_14_378 ();
 FILLCELL_X1 FILLER_15_7 ();
 FILLCELL_X2 FILLER_15_42 ();
 FILLCELL_X1 FILLER_15_85 ();
 FILLCELL_X2 FILLER_15_106 ();
 FILLCELL_X1 FILLER_15_144 ();
 FILLCELL_X4 FILLER_15_190 ();
 FILLCELL_X8 FILLER_15_198 ();
 FILLCELL_X4 FILLER_15_206 ();
 FILLCELL_X2 FILLER_15_221 ();
 FILLCELL_X1 FILLER_15_223 ();
 FILLCELL_X8 FILLER_15_256 ();
 FILLCELL_X4 FILLER_15_264 ();
 FILLCELL_X1 FILLER_15_268 ();
 FILLCELL_X2 FILLER_15_278 ();
 FILLCELL_X1 FILLER_15_302 ();
 FILLCELL_X2 FILLER_15_315 ();
 FILLCELL_X1 FILLER_15_331 ();
 FILLCELL_X2 FILLER_15_349 ();
 FILLCELL_X1 FILLER_15_351 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X8 FILLER_16_17 ();
 FILLCELL_X4 FILLER_16_25 ();
 FILLCELL_X2 FILLER_16_29 ();
 FILLCELL_X1 FILLER_16_31 ();
 FILLCELL_X8 FILLER_16_36 ();
 FILLCELL_X2 FILLER_16_44 ();
 FILLCELL_X1 FILLER_16_46 ();
 FILLCELL_X2 FILLER_16_71 ();
 FILLCELL_X16 FILLER_16_77 ();
 FILLCELL_X2 FILLER_16_93 ();
 FILLCELL_X1 FILLER_16_95 ();
 FILLCELL_X2 FILLER_16_99 ();
 FILLCELL_X4 FILLER_16_110 ();
 FILLCELL_X2 FILLER_16_114 ();
 FILLCELL_X1 FILLER_16_137 ();
 FILLCELL_X2 FILLER_16_145 ();
 FILLCELL_X2 FILLER_16_184 ();
 FILLCELL_X1 FILLER_16_206 ();
 FILLCELL_X1 FILLER_16_213 ();
 FILLCELL_X1 FILLER_16_240 ();
 FILLCELL_X2 FILLER_16_246 ();
 FILLCELL_X8 FILLER_16_254 ();
 FILLCELL_X2 FILLER_16_262 ();
 FILLCELL_X1 FILLER_16_264 ();
 FILLCELL_X8 FILLER_16_268 ();
 FILLCELL_X4 FILLER_16_276 ();
 FILLCELL_X2 FILLER_16_280 ();
 FILLCELL_X8 FILLER_16_287 ();
 FILLCELL_X2 FILLER_16_295 ();
 FILLCELL_X1 FILLER_16_297 ();
 FILLCELL_X4 FILLER_16_307 ();
 FILLCELL_X8 FILLER_16_358 ();
 FILLCELL_X2 FILLER_16_369 ();
 FILLCELL_X1 FILLER_16_371 ();
 FILLCELL_X1 FILLER_16_375 ();
 FILLCELL_X2 FILLER_16_383 ();
 FILLCELL_X1 FILLER_16_385 ();
 FILLCELL_X2 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_6 ();
 FILLCELL_X1 FILLER_17_8 ();
 FILLCELL_X2 FILLER_17_12 ();
 FILLCELL_X1 FILLER_17_14 ();
 FILLCELL_X4 FILLER_17_21 ();
 FILLCELL_X8 FILLER_17_51 ();
 FILLCELL_X4 FILLER_17_59 ();
 FILLCELL_X1 FILLER_17_63 ();
 FILLCELL_X4 FILLER_17_91 ();
 FILLCELL_X4 FILLER_17_108 ();
 FILLCELL_X1 FILLER_17_112 ();
 FILLCELL_X4 FILLER_17_123 ();
 FILLCELL_X2 FILLER_17_139 ();
 FILLCELL_X2 FILLER_17_148 ();
 FILLCELL_X1 FILLER_17_150 ();
 FILLCELL_X4 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_181 ();
 FILLCELL_X2 FILLER_17_196 ();
 FILLCELL_X1 FILLER_17_198 ();
 FILLCELL_X4 FILLER_17_206 ();
 FILLCELL_X2 FILLER_17_210 ();
 FILLCELL_X1 FILLER_17_260 ();
 FILLCELL_X4 FILLER_17_278 ();
 FILLCELL_X2 FILLER_17_303 ();
 FILLCELL_X1 FILLER_17_305 ();
 FILLCELL_X2 FILLER_17_311 ();
 FILLCELL_X4 FILLER_17_322 ();
 FILLCELL_X2 FILLER_17_326 ();
 FILLCELL_X4 FILLER_17_333 ();
 FILLCELL_X2 FILLER_17_337 ();
 FILLCELL_X2 FILLER_17_380 ();
 FILLCELL_X1 FILLER_17_382 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_33 ();
 FILLCELL_X2 FILLER_18_37 ();
 FILLCELL_X1 FILLER_18_39 ();
 FILLCELL_X4 FILLER_18_43 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X1 FILLER_18_55 ();
 FILLCELL_X4 FILLER_18_60 ();
 FILLCELL_X2 FILLER_18_64 ();
 FILLCELL_X1 FILLER_18_66 ();
 FILLCELL_X4 FILLER_18_72 ();
 FILLCELL_X1 FILLER_18_76 ();
 FILLCELL_X8 FILLER_18_81 ();
 FILLCELL_X1 FILLER_18_89 ();
 FILLCELL_X4 FILLER_18_95 ();
 FILLCELL_X2 FILLER_18_99 ();
 FILLCELL_X1 FILLER_18_101 ();
 FILLCELL_X1 FILLER_18_108 ();
 FILLCELL_X1 FILLER_18_113 ();
 FILLCELL_X4 FILLER_18_127 ();
 FILLCELL_X2 FILLER_18_131 ();
 FILLCELL_X2 FILLER_18_150 ();
 FILLCELL_X2 FILLER_18_154 ();
 FILLCELL_X2 FILLER_18_199 ();
 FILLCELL_X1 FILLER_18_201 ();
 FILLCELL_X2 FILLER_18_217 ();
 FILLCELL_X1 FILLER_18_219 ();
 FILLCELL_X4 FILLER_18_235 ();
 FILLCELL_X8 FILLER_18_248 ();
 FILLCELL_X1 FILLER_18_256 ();
 FILLCELL_X4 FILLER_18_271 ();
 FILLCELL_X2 FILLER_18_275 ();
 FILLCELL_X1 FILLER_18_284 ();
 FILLCELL_X16 FILLER_18_320 ();
 FILLCELL_X4 FILLER_18_336 ();
 FILLCELL_X2 FILLER_18_340 ();
 FILLCELL_X4 FILLER_18_355 ();
 FILLCELL_X2 FILLER_18_359 ();
 FILLCELL_X1 FILLER_18_361 ();
 FILLCELL_X2 FILLER_18_365 ();
 FILLCELL_X2 FILLER_18_384 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X2 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_15 ();
 FILLCELL_X32 FILLER_19_19 ();
 FILLCELL_X1 FILLER_19_51 ();
 FILLCELL_X8 FILLER_19_59 ();
 FILLCELL_X4 FILLER_19_89 ();
 FILLCELL_X1 FILLER_19_93 ();
 FILLCELL_X4 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_111 ();
 FILLCELL_X8 FILLER_19_122 ();
 FILLCELL_X1 FILLER_19_139 ();
 FILLCELL_X1 FILLER_19_176 ();
 FILLCELL_X1 FILLER_19_238 ();
 FILLCELL_X16 FILLER_19_246 ();
 FILLCELL_X2 FILLER_19_281 ();
 FILLCELL_X2 FILLER_19_290 ();
 FILLCELL_X2 FILLER_19_305 ();
 FILLCELL_X1 FILLER_19_307 ();
 FILLCELL_X1 FILLER_19_312 ();
 FILLCELL_X1 FILLER_19_317 ();
 FILLCELL_X2 FILLER_19_326 ();
 FILLCELL_X2 FILLER_19_363 ();
 FILLCELL_X1 FILLER_19_365 ();
 FILLCELL_X1 FILLER_19_379 ();
 FILLCELL_X2 FILLER_19_383 ();
 FILLCELL_X1 FILLER_19_385 ();
 FILLCELL_X2 FILLER_20_4 ();
 FILLCELL_X1 FILLER_20_6 ();
 FILLCELL_X16 FILLER_20_10 ();
 FILLCELL_X8 FILLER_20_26 ();
 FILLCELL_X2 FILLER_20_34 ();
 FILLCELL_X1 FILLER_20_36 ();
 FILLCELL_X4 FILLER_20_43 ();
 FILLCELL_X1 FILLER_20_47 ();
 FILLCELL_X8 FILLER_20_76 ();
 FILLCELL_X2 FILLER_20_84 ();
 FILLCELL_X2 FILLER_20_105 ();
 FILLCELL_X8 FILLER_20_115 ();
 FILLCELL_X4 FILLER_20_123 ();
 FILLCELL_X2 FILLER_20_127 ();
 FILLCELL_X2 FILLER_20_164 ();
 FILLCELL_X2 FILLER_20_171 ();
 FILLCELL_X1 FILLER_20_173 ();
 FILLCELL_X4 FILLER_20_232 ();
 FILLCELL_X2 FILLER_20_236 ();
 FILLCELL_X1 FILLER_20_238 ();
 FILLCELL_X8 FILLER_20_246 ();
 FILLCELL_X4 FILLER_20_254 ();
 FILLCELL_X1 FILLER_20_277 ();
 FILLCELL_X16 FILLER_20_288 ();
 FILLCELL_X4 FILLER_20_304 ();
 FILLCELL_X1 FILLER_20_313 ();
 FILLCELL_X16 FILLER_20_319 ();
 FILLCELL_X2 FILLER_20_335 ();
 FILLCELL_X1 FILLER_20_337 ();
 FILLCELL_X2 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_3 ();
 FILLCELL_X8 FILLER_21_10 ();
 FILLCELL_X4 FILLER_21_18 ();
 FILLCELL_X2 FILLER_21_22 ();
 FILLCELL_X8 FILLER_21_55 ();
 FILLCELL_X2 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_71 ();
 FILLCELL_X4 FILLER_21_79 ();
 FILLCELL_X2 FILLER_21_83 ();
 FILLCELL_X16 FILLER_21_90 ();
 FILLCELL_X8 FILLER_21_106 ();
 FILLCELL_X8 FILLER_21_120 ();
 FILLCELL_X4 FILLER_21_128 ();
 FILLCELL_X4 FILLER_21_140 ();
 FILLCELL_X1 FILLER_21_144 ();
 FILLCELL_X1 FILLER_21_150 ();
 FILLCELL_X4 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_165 ();
 FILLCELL_X1 FILLER_21_167 ();
 FILLCELL_X4 FILLER_21_171 ();
 FILLCELL_X1 FILLER_21_175 ();
 FILLCELL_X4 FILLER_21_182 ();
 FILLCELL_X2 FILLER_21_186 ();
 FILLCELL_X1 FILLER_21_197 ();
 FILLCELL_X2 FILLER_21_234 ();
 FILLCELL_X1 FILLER_21_240 ();
 FILLCELL_X8 FILLER_21_251 ();
 FILLCELL_X4 FILLER_21_259 ();
 FILLCELL_X2 FILLER_21_263 ();
 FILLCELL_X1 FILLER_21_265 ();
 FILLCELL_X4 FILLER_21_279 ();
 FILLCELL_X2 FILLER_21_287 ();
 FILLCELL_X1 FILLER_21_289 ();
 FILLCELL_X16 FILLER_21_293 ();
 FILLCELL_X8 FILLER_21_309 ();
 FILLCELL_X1 FILLER_21_317 ();
 FILLCELL_X8 FILLER_21_337 ();
 FILLCELL_X4 FILLER_21_345 ();
 FILLCELL_X1 FILLER_21_349 ();
 FILLCELL_X4 FILLER_21_353 ();
 FILLCELL_X2 FILLER_21_384 ();
 FILLCELL_X8 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_9 ();
 FILLCELL_X1 FILLER_22_13 ();
 FILLCELL_X1 FILLER_22_40 ();
 FILLCELL_X8 FILLER_22_43 ();
 FILLCELL_X2 FILLER_22_51 ();
 FILLCELL_X1 FILLER_22_53 ();
 FILLCELL_X2 FILLER_22_87 ();
 FILLCELL_X1 FILLER_22_89 ();
 FILLCELL_X2 FILLER_22_94 ();
 FILLCELL_X1 FILLER_22_122 ();
 FILLCELL_X1 FILLER_22_128 ();
 FILLCELL_X2 FILLER_22_153 ();
 FILLCELL_X2 FILLER_22_177 ();
 FILLCELL_X4 FILLER_22_184 ();
 FILLCELL_X4 FILLER_22_195 ();
 FILLCELL_X1 FILLER_22_203 ();
 FILLCELL_X4 FILLER_22_207 ();
 FILLCELL_X2 FILLER_22_211 ();
 FILLCELL_X2 FILLER_22_245 ();
 FILLCELL_X1 FILLER_22_247 ();
 FILLCELL_X2 FILLER_22_287 ();
 FILLCELL_X2 FILLER_22_294 ();
 FILLCELL_X4 FILLER_22_306 ();
 FILLCELL_X2 FILLER_22_314 ();
 FILLCELL_X1 FILLER_22_316 ();
 FILLCELL_X8 FILLER_22_329 ();
 FILLCELL_X4 FILLER_22_337 ();
 FILLCELL_X4 FILLER_22_348 ();
 FILLCELL_X2 FILLER_22_352 ();
 FILLCELL_X8 FILLER_22_357 ();
 FILLCELL_X1 FILLER_22_365 ();
 FILLCELL_X4 FILLER_22_379 ();
 FILLCELL_X2 FILLER_22_383 ();
 FILLCELL_X1 FILLER_22_385 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_9 ();
 FILLCELL_X2 FILLER_23_13 ();
 FILLCELL_X16 FILLER_23_18 ();
 FILLCELL_X4 FILLER_23_34 ();
 FILLCELL_X1 FILLER_23_38 ();
 FILLCELL_X2 FILLER_23_87 ();
 FILLCELL_X1 FILLER_23_92 ();
 FILLCELL_X8 FILLER_23_95 ();
 FILLCELL_X1 FILLER_23_103 ();
 FILLCELL_X4 FILLER_23_118 ();
 FILLCELL_X2 FILLER_23_122 ();
 FILLCELL_X1 FILLER_23_124 ();
 FILLCELL_X1 FILLER_23_133 ();
 FILLCELL_X8 FILLER_23_155 ();
 FILLCELL_X8 FILLER_23_174 ();
 FILLCELL_X1 FILLER_23_214 ();
 FILLCELL_X2 FILLER_23_222 ();
 FILLCELL_X2 FILLER_23_227 ();
 FILLCELL_X2 FILLER_23_240 ();
 FILLCELL_X4 FILLER_23_246 ();
 FILLCELL_X1 FILLER_23_250 ();
 FILLCELL_X1 FILLER_23_284 ();
 FILLCELL_X4 FILLER_23_306 ();
 FILLCELL_X1 FILLER_23_310 ();
 FILLCELL_X2 FILLER_23_315 ();
 FILLCELL_X1 FILLER_23_317 ();
 FILLCELL_X2 FILLER_23_340 ();
 FILLCELL_X1 FILLER_23_367 ();
 FILLCELL_X2 FILLER_23_378 ();
 FILLCELL_X1 FILLER_23_380 ();
 FILLCELL_X2 FILLER_23_384 ();
 FILLCELL_X2 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_6 ();
 FILLCELL_X1 FILLER_24_22 ();
 FILLCELL_X8 FILLER_24_30 ();
 FILLCELL_X4 FILLER_24_38 ();
 FILLCELL_X2 FILLER_24_75 ();
 FILLCELL_X1 FILLER_24_95 ();
 FILLCELL_X1 FILLER_24_104 ();
 FILLCELL_X1 FILLER_24_133 ();
 FILLCELL_X1 FILLER_24_143 ();
 FILLCELL_X2 FILLER_24_154 ();
 FILLCELL_X1 FILLER_24_163 ();
 FILLCELL_X1 FILLER_24_173 ();
 FILLCELL_X4 FILLER_24_223 ();
 FILLCELL_X1 FILLER_24_227 ();
 FILLCELL_X2 FILLER_24_251 ();
 FILLCELL_X2 FILLER_24_264 ();
 FILLCELL_X1 FILLER_24_266 ();
 FILLCELL_X2 FILLER_24_271 ();
 FILLCELL_X1 FILLER_24_273 ();
 FILLCELL_X2 FILLER_24_285 ();
 FILLCELL_X1 FILLER_24_291 ();
 FILLCELL_X4 FILLER_24_295 ();
 FILLCELL_X2 FILLER_24_299 ();
 FILLCELL_X1 FILLER_24_301 ();
 FILLCELL_X4 FILLER_24_307 ();
 FILLCELL_X4 FILLER_24_321 ();
 FILLCELL_X2 FILLER_24_330 ();
 FILLCELL_X2 FILLER_24_351 ();
 FILLCELL_X2 FILLER_24_360 ();
 FILLCELL_X1 FILLER_24_362 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_12 ();
 FILLCELL_X4 FILLER_25_20 ();
 FILLCELL_X16 FILLER_25_43 ();
 FILLCELL_X1 FILLER_25_59 ();
 FILLCELL_X4 FILLER_25_79 ();
 FILLCELL_X2 FILLER_25_106 ();
 FILLCELL_X2 FILLER_25_139 ();
 FILLCELL_X2 FILLER_25_143 ();
 FILLCELL_X1 FILLER_25_148 ();
 FILLCELL_X8 FILLER_25_191 ();
 FILLCELL_X2 FILLER_25_199 ();
 FILLCELL_X2 FILLER_25_223 ();
 FILLCELL_X2 FILLER_25_246 ();
 FILLCELL_X1 FILLER_25_252 ();
 FILLCELL_X8 FILLER_25_256 ();
 FILLCELL_X32 FILLER_25_271 ();
 FILLCELL_X2 FILLER_25_303 ();
 FILLCELL_X1 FILLER_25_305 ();
 FILLCELL_X1 FILLER_25_310 ();
 FILLCELL_X2 FILLER_25_316 ();
 FILLCELL_X8 FILLER_25_327 ();
 FILLCELL_X2 FILLER_25_335 ();
 FILLCELL_X4 FILLER_25_366 ();
 FILLCELL_X2 FILLER_25_370 ();
 FILLCELL_X4 FILLER_25_380 ();
 FILLCELL_X2 FILLER_25_384 ();
 FILLCELL_X4 FILLER_26_29 ();
 FILLCELL_X1 FILLER_26_69 ();
 FILLCELL_X1 FILLER_26_76 ();
 FILLCELL_X2 FILLER_26_92 ();
 FILLCELL_X1 FILLER_26_102 ();
 FILLCELL_X1 FILLER_26_113 ();
 FILLCELL_X4 FILLER_26_128 ();
 FILLCELL_X1 FILLER_26_132 ();
 FILLCELL_X4 FILLER_26_136 ();
 FILLCELL_X1 FILLER_26_150 ();
 FILLCELL_X1 FILLER_26_162 ();
 FILLCELL_X1 FILLER_26_167 ();
 FILLCELL_X1 FILLER_26_179 ();
 FILLCELL_X2 FILLER_26_194 ();
 FILLCELL_X2 FILLER_26_227 ();
 FILLCELL_X8 FILLER_26_254 ();
 FILLCELL_X4 FILLER_26_262 ();
 FILLCELL_X4 FILLER_26_289 ();
 FILLCELL_X2 FILLER_26_293 ();
 FILLCELL_X1 FILLER_26_295 ();
 FILLCELL_X1 FILLER_26_305 ();
 FILLCELL_X1 FILLER_26_323 ();
 FILLCELL_X16 FILLER_26_328 ();
 FILLCELL_X4 FILLER_26_344 ();
 FILLCELL_X2 FILLER_26_352 ();
 FILLCELL_X8 FILLER_26_357 ();
 FILLCELL_X4 FILLER_27_1 ();
 FILLCELL_X1 FILLER_27_5 ();
 FILLCELL_X8 FILLER_27_9 ();
 FILLCELL_X4 FILLER_27_17 ();
 FILLCELL_X1 FILLER_27_21 ();
 FILLCELL_X1 FILLER_27_46 ();
 FILLCELL_X32 FILLER_27_54 ();
 FILLCELL_X1 FILLER_27_86 ();
 FILLCELL_X4 FILLER_27_94 ();
 FILLCELL_X2 FILLER_27_98 ();
 FILLCELL_X1 FILLER_27_100 ();
 FILLCELL_X2 FILLER_27_104 ();
 FILLCELL_X1 FILLER_27_106 ();
 FILLCELL_X2 FILLER_27_123 ();
 FILLCELL_X2 FILLER_27_132 ();
 FILLCELL_X4 FILLER_27_169 ();
 FILLCELL_X1 FILLER_27_173 ();
 FILLCELL_X1 FILLER_27_181 ();
 FILLCELL_X2 FILLER_27_206 ();
 FILLCELL_X1 FILLER_27_208 ();
 FILLCELL_X1 FILLER_27_214 ();
 FILLCELL_X2 FILLER_27_219 ();
 FILLCELL_X2 FILLER_27_226 ();
 FILLCELL_X1 FILLER_27_228 ();
 FILLCELL_X1 FILLER_27_238 ();
 FILLCELL_X4 FILLER_27_244 ();
 FILLCELL_X2 FILLER_27_248 ();
 FILLCELL_X1 FILLER_27_260 ();
 FILLCELL_X2 FILLER_27_276 ();
 FILLCELL_X1 FILLER_27_278 ();
 FILLCELL_X1 FILLER_27_282 ();
 FILLCELL_X2 FILLER_27_294 ();
 FILLCELL_X1 FILLER_27_302 ();
 FILLCELL_X2 FILLER_27_307 ();
 FILLCELL_X4 FILLER_27_331 ();
 FILLCELL_X2 FILLER_27_335 ();
 FILLCELL_X1 FILLER_27_337 ();
 FILLCELL_X1 FILLER_27_382 ();
 FILLCELL_X4 FILLER_28_25 ();
 FILLCELL_X16 FILLER_28_36 ();
 FILLCELL_X4 FILLER_28_52 ();
 FILLCELL_X2 FILLER_28_56 ();
 FILLCELL_X1 FILLER_28_58 ();
 FILLCELL_X2 FILLER_28_104 ();
 FILLCELL_X1 FILLER_28_118 ();
 FILLCELL_X2 FILLER_28_123 ();
 FILLCELL_X4 FILLER_28_143 ();
 FILLCELL_X2 FILLER_28_147 ();
 FILLCELL_X1 FILLER_28_149 ();
 FILLCELL_X1 FILLER_28_153 ();
 FILLCELL_X2 FILLER_28_168 ();
 FILLCELL_X1 FILLER_28_193 ();
 FILLCELL_X8 FILLER_28_197 ();
 FILLCELL_X4 FILLER_28_205 ();
 FILLCELL_X4 FILLER_28_225 ();
 FILLCELL_X8 FILLER_28_233 ();
 FILLCELL_X4 FILLER_28_248 ();
 FILLCELL_X1 FILLER_28_272 ();
 FILLCELL_X1 FILLER_28_277 ();
 FILLCELL_X1 FILLER_28_320 ();
 FILLCELL_X1 FILLER_28_330 ();
 FILLCELL_X4 FILLER_28_335 ();
 FILLCELL_X2 FILLER_28_339 ();
 FILLCELL_X1 FILLER_28_341 ();
 FILLCELL_X8 FILLER_28_349 ();
 FILLCELL_X4 FILLER_28_364 ();
 FILLCELL_X2 FILLER_28_368 ();
 FILLCELL_X2 FILLER_28_377 ();
 FILLCELL_X1 FILLER_28_379 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_27 ();
 FILLCELL_X2 FILLER_29_31 ();
 FILLCELL_X1 FILLER_29_33 ();
 FILLCELL_X4 FILLER_29_53 ();
 FILLCELL_X2 FILLER_29_57 ();
 FILLCELL_X1 FILLER_29_59 ();
 FILLCELL_X2 FILLER_29_72 ();
 FILLCELL_X1 FILLER_29_74 ();
 FILLCELL_X2 FILLER_29_85 ();
 FILLCELL_X1 FILLER_29_87 ();
 FILLCELL_X2 FILLER_29_93 ();
 FILLCELL_X2 FILLER_29_99 ();
 FILLCELL_X1 FILLER_29_118 ();
 FILLCELL_X2 FILLER_29_132 ();
 FILLCELL_X2 FILLER_29_150 ();
 FILLCELL_X4 FILLER_29_166 ();
 FILLCELL_X4 FILLER_29_173 ();
 FILLCELL_X2 FILLER_29_177 ();
 FILLCELL_X1 FILLER_29_179 ();
 FILLCELL_X4 FILLER_29_185 ();
 FILLCELL_X2 FILLER_29_189 ();
 FILLCELL_X4 FILLER_29_205 ();
 FILLCELL_X1 FILLER_29_209 ();
 FILLCELL_X8 FILLER_29_217 ();
 FILLCELL_X1 FILLER_29_225 ();
 FILLCELL_X1 FILLER_29_231 ();
 FILLCELL_X2 FILLER_29_239 ();
 FILLCELL_X1 FILLER_29_250 ();
 FILLCELL_X2 FILLER_29_258 ();
 FILLCELL_X2 FILLER_29_274 ();
 FILLCELL_X1 FILLER_29_276 ();
 FILLCELL_X4 FILLER_29_281 ();
 FILLCELL_X1 FILLER_29_285 ();
 FILLCELL_X1 FILLER_29_289 ();
 FILLCELL_X1 FILLER_29_300 ();
 FILLCELL_X8 FILLER_29_306 ();
 FILLCELL_X4 FILLER_29_318 ();
 FILLCELL_X2 FILLER_29_322 ();
 FILLCELL_X1 FILLER_29_324 ();
 FILLCELL_X8 FILLER_29_329 ();
 FILLCELL_X2 FILLER_29_337 ();
 FILLCELL_X2 FILLER_29_367 ();
 FILLCELL_X1 FILLER_30_11 ();
 FILLCELL_X1 FILLER_30_19 ();
 FILLCELL_X2 FILLER_30_30 ();
 FILLCELL_X16 FILLER_30_39 ();
 FILLCELL_X4 FILLER_30_55 ();
 FILLCELL_X2 FILLER_30_59 ();
 FILLCELL_X1 FILLER_30_71 ();
 FILLCELL_X8 FILLER_30_76 ();
 FILLCELL_X4 FILLER_30_84 ();
 FILLCELL_X2 FILLER_30_88 ();
 FILLCELL_X1 FILLER_30_95 ();
 FILLCELL_X2 FILLER_30_144 ();
 FILLCELL_X2 FILLER_30_159 ();
 FILLCELL_X1 FILLER_30_176 ();
 FILLCELL_X8 FILLER_30_190 ();
 FILLCELL_X4 FILLER_30_202 ();
 FILLCELL_X2 FILLER_30_206 ();
 FILLCELL_X1 FILLER_30_216 ();
 FILLCELL_X1 FILLER_30_234 ();
 FILLCELL_X2 FILLER_30_249 ();
 FILLCELL_X1 FILLER_30_251 ();
 FILLCELL_X1 FILLER_30_256 ();
 FILLCELL_X1 FILLER_30_266 ();
 FILLCELL_X4 FILLER_30_271 ();
 FILLCELL_X2 FILLER_30_305 ();
 FILLCELL_X1 FILLER_30_312 ();
 FILLCELL_X4 FILLER_30_331 ();
 FILLCELL_X2 FILLER_30_362 ();
 FILLCELL_X1 FILLER_30_364 ();
 FILLCELL_X1 FILLER_30_377 ();
 FILLCELL_X1 FILLER_30_381 ();
 FILLCELL_X2 FILLER_31_4 ();
 FILLCELL_X32 FILLER_31_47 ();
 FILLCELL_X2 FILLER_31_79 ();
 FILLCELL_X1 FILLER_31_83 ();
 FILLCELL_X4 FILLER_31_96 ();
 FILLCELL_X1 FILLER_31_100 ();
 FILLCELL_X4 FILLER_31_128 ();
 FILLCELL_X1 FILLER_31_150 ();
 FILLCELL_X1 FILLER_31_160 ();
 FILLCELL_X4 FILLER_31_172 ();
 FILLCELL_X2 FILLER_31_176 ();
 FILLCELL_X4 FILLER_31_185 ();
 FILLCELL_X2 FILLER_31_189 ();
 FILLCELL_X8 FILLER_31_213 ();
 FILLCELL_X1 FILLER_31_221 ();
 FILLCELL_X1 FILLER_31_234 ();
 FILLCELL_X2 FILLER_31_239 ();
 FILLCELL_X1 FILLER_31_241 ();
 FILLCELL_X8 FILLER_31_265 ();
 FILLCELL_X2 FILLER_31_273 ();
 FILLCELL_X8 FILLER_31_290 ();
 FILLCELL_X4 FILLER_31_298 ();
 FILLCELL_X2 FILLER_31_302 ();
 FILLCELL_X1 FILLER_31_304 ();
 FILLCELL_X4 FILLER_31_310 ();
 FILLCELL_X1 FILLER_31_314 ();
 FILLCELL_X16 FILLER_31_320 ();
 FILLCELL_X4 FILLER_31_336 ();
 FILLCELL_X2 FILLER_31_340 ();
 FILLCELL_X4 FILLER_31_346 ();
 FILLCELL_X1 FILLER_31_350 ();
 FILLCELL_X16 FILLER_31_357 ();
 FILLCELL_X2 FILLER_31_383 ();
 FILLCELL_X1 FILLER_31_385 ();
 FILLCELL_X4 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_11 ();
 FILLCELL_X2 FILLER_32_19 ();
 FILLCELL_X8 FILLER_32_24 ();
 FILLCELL_X2 FILLER_32_32 ();
 FILLCELL_X16 FILLER_32_53 ();
 FILLCELL_X8 FILLER_32_69 ();
 FILLCELL_X2 FILLER_32_77 ();
 FILLCELL_X1 FILLER_32_79 ();
 FILLCELL_X2 FILLER_32_100 ();
 FILLCELL_X1 FILLER_32_102 ();
 FILLCELL_X2 FILLER_32_123 ();
 FILLCELL_X4 FILLER_32_131 ();
 FILLCELL_X1 FILLER_32_135 ();
 FILLCELL_X4 FILLER_32_141 ();
 FILLCELL_X2 FILLER_32_145 ();
 FILLCELL_X4 FILLER_32_157 ();
 FILLCELL_X1 FILLER_32_161 ();
 FILLCELL_X1 FILLER_32_179 ();
 FILLCELL_X2 FILLER_32_220 ();
 FILLCELL_X1 FILLER_32_222 ();
 FILLCELL_X4 FILLER_32_233 ();
 FILLCELL_X1 FILLER_32_237 ();
 FILLCELL_X2 FILLER_32_265 ();
 FILLCELL_X1 FILLER_32_277 ();
 FILLCELL_X2 FILLER_32_285 ();
 FILLCELL_X4 FILLER_32_293 ();
 FILLCELL_X1 FILLER_32_297 ();
 FILLCELL_X1 FILLER_32_304 ();
 FILLCELL_X4 FILLER_32_314 ();
 FILLCELL_X2 FILLER_32_318 ();
 FILLCELL_X4 FILLER_32_324 ();
 FILLCELL_X1 FILLER_32_328 ();
 FILLCELL_X4 FILLER_32_350 ();
 FILLCELL_X1 FILLER_32_354 ();
 FILLCELL_X4 FILLER_32_362 ();
 FILLCELL_X4 FILLER_32_380 ();
 FILLCELL_X2 FILLER_32_384 ();
 FILLCELL_X1 FILLER_33_4 ();
 FILLCELL_X8 FILLER_33_21 ();
 FILLCELL_X1 FILLER_33_41 ();
 FILLCELL_X2 FILLER_33_59 ();
 FILLCELL_X2 FILLER_33_95 ();
 FILLCELL_X8 FILLER_33_101 ();
 FILLCELL_X1 FILLER_33_109 ();
 FILLCELL_X8 FILLER_33_123 ();
 FILLCELL_X16 FILLER_33_145 ();
 FILLCELL_X4 FILLER_33_161 ();
 FILLCELL_X1 FILLER_33_165 ();
 FILLCELL_X4 FILLER_33_173 ();
 FILLCELL_X2 FILLER_33_188 ();
 FILLCELL_X4 FILLER_33_197 ();
 FILLCELL_X2 FILLER_33_201 ();
 FILLCELL_X8 FILLER_33_210 ();
 FILLCELL_X1 FILLER_33_218 ();
 FILLCELL_X8 FILLER_33_238 ();
 FILLCELL_X1 FILLER_33_246 ();
 FILLCELL_X1 FILLER_33_258 ();
 FILLCELL_X1 FILLER_33_270 ();
 FILLCELL_X1 FILLER_33_277 ();
 FILLCELL_X4 FILLER_33_286 ();
 FILLCELL_X1 FILLER_33_290 ();
 FILLCELL_X2 FILLER_33_302 ();
 FILLCELL_X1 FILLER_33_309 ();
 FILLCELL_X4 FILLER_33_314 ();
 FILLCELL_X1 FILLER_33_318 ();
 FILLCELL_X1 FILLER_33_328 ();
 FILLCELL_X1 FILLER_33_340 ();
 FILLCELL_X1 FILLER_33_368 ();
 FILLCELL_X1 FILLER_34_4 ();
 FILLCELL_X1 FILLER_34_48 ();
 FILLCELL_X32 FILLER_34_73 ();
 FILLCELL_X8 FILLER_34_105 ();
 FILLCELL_X2 FILLER_34_126 ();
 FILLCELL_X2 FILLER_34_131 ();
 FILLCELL_X4 FILLER_34_149 ();
 FILLCELL_X2 FILLER_34_153 ();
 FILLCELL_X1 FILLER_34_155 ();
 FILLCELL_X2 FILLER_34_159 ();
 FILLCELL_X4 FILLER_34_175 ();
 FILLCELL_X2 FILLER_34_198 ();
 FILLCELL_X1 FILLER_34_209 ();
 FILLCELL_X2 FILLER_34_213 ();
 FILLCELL_X1 FILLER_34_215 ();
 FILLCELL_X4 FILLER_34_224 ();
 FILLCELL_X16 FILLER_34_244 ();
 FILLCELL_X8 FILLER_34_260 ();
 FILLCELL_X4 FILLER_34_268 ();
 FILLCELL_X2 FILLER_34_282 ();
 FILLCELL_X1 FILLER_34_284 ();
 FILLCELL_X8 FILLER_34_301 ();
 FILLCELL_X2 FILLER_34_313 ();
 FILLCELL_X1 FILLER_34_335 ();
 FILLCELL_X2 FILLER_34_357 ();
 FILLCELL_X1 FILLER_34_359 ();
 FILLCELL_X1 FILLER_34_363 ();
 FILLCELL_X8 FILLER_34_367 ();
 FILLCELL_X1 FILLER_34_382 ();
 FILLCELL_X4 FILLER_35_25 ();
 FILLCELL_X4 FILLER_35_36 ();
 FILLCELL_X2 FILLER_35_40 ();
 FILLCELL_X4 FILLER_35_62 ();
 FILLCELL_X1 FILLER_35_66 ();
 FILLCELL_X1 FILLER_35_110 ();
 FILLCELL_X1 FILLER_35_138 ();
 FILLCELL_X2 FILLER_35_175 ();
 FILLCELL_X8 FILLER_35_181 ();
 FILLCELL_X2 FILLER_35_189 ();
 FILLCELL_X2 FILLER_35_196 ();
 FILLCELL_X1 FILLER_35_198 ();
 FILLCELL_X1 FILLER_35_203 ();
 FILLCELL_X1 FILLER_35_209 ();
 FILLCELL_X1 FILLER_35_220 ();
 FILLCELL_X4 FILLER_35_240 ();
 FILLCELL_X1 FILLER_35_244 ();
 FILLCELL_X4 FILLER_35_249 ();
 FILLCELL_X2 FILLER_35_253 ();
 FILLCELL_X2 FILLER_35_261 ();
 FILLCELL_X8 FILLER_35_269 ();
 FILLCELL_X16 FILLER_35_292 ();
 FILLCELL_X4 FILLER_35_317 ();
 FILLCELL_X2 FILLER_35_321 ();
 FILLCELL_X4 FILLER_35_332 ();
 FILLCELL_X2 FILLER_35_336 ();
 FILLCELL_X1 FILLER_35_338 ();
 FILLCELL_X4 FILLER_35_367 ();
 FILLCELL_X2 FILLER_35_371 ();
 FILLCELL_X4 FILLER_35_380 ();
 FILLCELL_X2 FILLER_35_384 ();
 FILLCELL_X2 FILLER_36_24 ();
 FILLCELL_X1 FILLER_36_26 ();
 FILLCELL_X2 FILLER_36_49 ();
 FILLCELL_X1 FILLER_36_51 ();
 FILLCELL_X2 FILLER_36_71 ();
 FILLCELL_X1 FILLER_36_73 ();
 FILLCELL_X16 FILLER_36_81 ();
 FILLCELL_X4 FILLER_36_97 ();
 FILLCELL_X2 FILLER_36_101 ();
 FILLCELL_X4 FILLER_36_110 ();
 FILLCELL_X2 FILLER_36_114 ();
 FILLCELL_X16 FILLER_36_137 ();
 FILLCELL_X2 FILLER_36_153 ();
 FILLCELL_X1 FILLER_36_155 ();
 FILLCELL_X4 FILLER_36_193 ();
 FILLCELL_X2 FILLER_36_197 ();
 FILLCELL_X1 FILLER_36_221 ();
 FILLCELL_X2 FILLER_36_228 ();
 FILLCELL_X1 FILLER_36_230 ();
 FILLCELL_X1 FILLER_36_236 ();
 FILLCELL_X1 FILLER_36_241 ();
 FILLCELL_X1 FILLER_36_250 ();
 FILLCELL_X1 FILLER_36_276 ();
 FILLCELL_X4 FILLER_36_281 ();
 FILLCELL_X1 FILLER_36_312 ();
 FILLCELL_X1 FILLER_36_322 ();
 FILLCELL_X4 FILLER_36_332 ();
 FILLCELL_X2 FILLER_36_336 ();
 FILLCELL_X1 FILLER_36_338 ();
 FILLCELL_X4 FILLER_36_342 ();
 FILLCELL_X1 FILLER_36_346 ();
 FILLCELL_X2 FILLER_36_367 ();
 FILLCELL_X1 FILLER_37_1 ();
 FILLCELL_X4 FILLER_37_12 ();
 FILLCELL_X4 FILLER_37_39 ();
 FILLCELL_X2 FILLER_37_43 ();
 FILLCELL_X16 FILLER_37_50 ();
 FILLCELL_X2 FILLER_37_81 ();
 FILLCELL_X4 FILLER_37_104 ();
 FILLCELL_X2 FILLER_37_108 ();
 FILLCELL_X2 FILLER_37_117 ();
 FILLCELL_X8 FILLER_37_122 ();
 FILLCELL_X1 FILLER_37_130 ();
 FILLCELL_X2 FILLER_37_134 ();
 FILLCELL_X1 FILLER_37_136 ();
 FILLCELL_X2 FILLER_37_140 ();
 FILLCELL_X4 FILLER_37_146 ();
 FILLCELL_X2 FILLER_37_150 ();
 FILLCELL_X2 FILLER_37_160 ();
 FILLCELL_X1 FILLER_37_162 ();
 FILLCELL_X4 FILLER_37_165 ();
 FILLCELL_X1 FILLER_37_169 ();
 FILLCELL_X8 FILLER_37_174 ();
 FILLCELL_X1 FILLER_37_187 ();
 FILLCELL_X2 FILLER_37_205 ();
 FILLCELL_X2 FILLER_37_217 ();
 FILLCELL_X2 FILLER_37_222 ();
 FILLCELL_X1 FILLER_37_242 ();
 FILLCELL_X1 FILLER_37_253 ();
 FILLCELL_X2 FILLER_37_260 ();
 FILLCELL_X1 FILLER_37_273 ();
 FILLCELL_X2 FILLER_37_313 ();
 FILLCELL_X8 FILLER_37_327 ();
 FILLCELL_X1 FILLER_37_335 ();
 FILLCELL_X4 FILLER_37_357 ();
 FILLCELL_X1 FILLER_37_375 ();
 FILLCELL_X2 FILLER_37_379 ();
 FILLCELL_X1 FILLER_37_381 ();
 FILLCELL_X4 FILLER_38_1 ();
 FILLCELL_X2 FILLER_38_5 ();
 FILLCELL_X1 FILLER_38_7 ();
 FILLCELL_X2 FILLER_38_11 ();
 FILLCELL_X1 FILLER_38_13 ();
 FILLCELL_X8 FILLER_38_24 ();
 FILLCELL_X8 FILLER_38_56 ();
 FILLCELL_X2 FILLER_38_64 ();
 FILLCELL_X1 FILLER_38_66 ();
 FILLCELL_X8 FILLER_38_84 ();
 FILLCELL_X1 FILLER_38_92 ();
 FILLCELL_X4 FILLER_38_100 ();
 FILLCELL_X2 FILLER_38_104 ();
 FILLCELL_X2 FILLER_38_113 ();
 FILLCELL_X8 FILLER_38_123 ();
 FILLCELL_X2 FILLER_38_131 ();
 FILLCELL_X1 FILLER_38_133 ();
 FILLCELL_X4 FILLER_38_180 ();
 FILLCELL_X2 FILLER_38_184 ();
 FILLCELL_X1 FILLER_38_186 ();
 FILLCELL_X8 FILLER_38_194 ();
 FILLCELL_X4 FILLER_38_202 ();
 FILLCELL_X1 FILLER_38_206 ();
 FILLCELL_X8 FILLER_38_212 ();
 FILLCELL_X1 FILLER_38_220 ();
 FILLCELL_X4 FILLER_38_230 ();
 FILLCELL_X2 FILLER_38_246 ();
 FILLCELL_X4 FILLER_38_252 ();
 FILLCELL_X2 FILLER_38_256 ();
 FILLCELL_X1 FILLER_38_258 ();
 FILLCELL_X1 FILLER_38_272 ();
 FILLCELL_X2 FILLER_38_277 ();
 FILLCELL_X2 FILLER_38_300 ();
 FILLCELL_X2 FILLER_38_312 ();
 FILLCELL_X2 FILLER_38_319 ();
 FILLCELL_X1 FILLER_38_321 ();
 FILLCELL_X4 FILLER_38_343 ();
 FILLCELL_X2 FILLER_38_347 ();
 FILLCELL_X1 FILLER_38_349 ();
 FILLCELL_X4 FILLER_38_378 ();
 FILLCELL_X1 FILLER_38_382 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X4 FILLER_39_33 ();
 FILLCELL_X8 FILLER_39_40 ();
 FILLCELL_X4 FILLER_39_48 ();
 FILLCELL_X2 FILLER_39_52 ();
 FILLCELL_X1 FILLER_39_54 ();
 FILLCELL_X8 FILLER_39_79 ();
 FILLCELL_X4 FILLER_39_87 ();
 FILLCELL_X1 FILLER_39_109 ();
 FILLCELL_X2 FILLER_39_127 ();
 FILLCELL_X1 FILLER_39_140 ();
 FILLCELL_X2 FILLER_39_145 ();
 FILLCELL_X1 FILLER_39_147 ();
 FILLCELL_X1 FILLER_39_160 ();
 FILLCELL_X8 FILLER_39_180 ();
 FILLCELL_X2 FILLER_39_188 ();
 FILLCELL_X2 FILLER_39_202 ();
 FILLCELL_X1 FILLER_39_204 ();
 FILLCELL_X1 FILLER_39_210 ();
 FILLCELL_X4 FILLER_39_217 ();
 FILLCELL_X2 FILLER_39_221 ();
 FILLCELL_X1 FILLER_39_223 ();
 FILLCELL_X1 FILLER_39_236 ();
 FILLCELL_X8 FILLER_39_241 ();
 FILLCELL_X4 FILLER_39_249 ();
 FILLCELL_X8 FILLER_39_258 ();
 FILLCELL_X4 FILLER_39_266 ();
 FILLCELL_X1 FILLER_39_270 ();
 FILLCELL_X2 FILLER_39_280 ();
 FILLCELL_X8 FILLER_39_291 ();
 FILLCELL_X2 FILLER_39_299 ();
 FILLCELL_X2 FILLER_39_329 ();
 FILLCELL_X1 FILLER_39_331 ();
 FILLCELL_X4 FILLER_39_339 ();
 FILLCELL_X2 FILLER_39_343 ();
 FILLCELL_X2 FILLER_39_352 ();
 FILLCELL_X2 FILLER_39_357 ();
 FILLCELL_X4 FILLER_40_1 ();
 FILLCELL_X2 FILLER_40_5 ();
 FILLCELL_X1 FILLER_40_10 ();
 FILLCELL_X1 FILLER_40_57 ();
 FILLCELL_X8 FILLER_40_65 ();
 FILLCELL_X4 FILLER_40_73 ();
 FILLCELL_X2 FILLER_40_77 ();
 FILLCELL_X1 FILLER_40_79 ();
 FILLCELL_X2 FILLER_40_104 ();
 FILLCELL_X1 FILLER_40_106 ();
 FILLCELL_X2 FILLER_40_122 ();
 FILLCELL_X4 FILLER_40_126 ();
 FILLCELL_X16 FILLER_40_144 ();
 FILLCELL_X8 FILLER_40_160 ();
 FILLCELL_X1 FILLER_40_168 ();
 FILLCELL_X2 FILLER_40_178 ();
 FILLCELL_X16 FILLER_40_185 ();
 FILLCELL_X2 FILLER_40_201 ();
 FILLCELL_X2 FILLER_40_211 ();
 FILLCELL_X1 FILLER_40_216 ();
 FILLCELL_X1 FILLER_40_229 ();
 FILLCELL_X2 FILLER_40_253 ();
 FILLCELL_X1 FILLER_40_255 ();
 FILLCELL_X8 FILLER_40_260 ();
 FILLCELL_X2 FILLER_40_268 ();
 FILLCELL_X32 FILLER_40_280 ();
 FILLCELL_X16 FILLER_40_312 ();
 FILLCELL_X1 FILLER_40_328 ();
 FILLCELL_X4 FILLER_40_353 ();
 FILLCELL_X2 FILLER_40_357 ();
 FILLCELL_X1 FILLER_40_359 ();
 FILLCELL_X2 FILLER_40_370 ();
 FILLCELL_X1 FILLER_40_372 ();
 FILLCELL_X4 FILLER_40_377 ();
 FILLCELL_X1 FILLER_40_385 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X2 FILLER_41_36 ();
 FILLCELL_X8 FILLER_41_45 ();
 FILLCELL_X4 FILLER_41_53 ();
 FILLCELL_X2 FILLER_41_57 ();
 FILLCELL_X16 FILLER_41_76 ();
 FILLCELL_X8 FILLER_41_92 ();
 FILLCELL_X4 FILLER_41_100 ();
 FILLCELL_X1 FILLER_41_104 ();
 FILLCELL_X4 FILLER_41_127 ();
 FILLCELL_X2 FILLER_41_131 ();
 FILLCELL_X4 FILLER_41_137 ();
 FILLCELL_X4 FILLER_41_145 ();
 FILLCELL_X1 FILLER_41_149 ();
 FILLCELL_X1 FILLER_41_153 ();
 FILLCELL_X1 FILLER_41_160 ();
 FILLCELL_X2 FILLER_41_167 ();
 FILLCELL_X1 FILLER_41_175 ();
 FILLCELL_X16 FILLER_41_180 ();
 FILLCELL_X4 FILLER_41_196 ();
 FILLCELL_X2 FILLER_41_200 ();
 FILLCELL_X1 FILLER_41_202 ();
 FILLCELL_X8 FILLER_41_207 ();
 FILLCELL_X2 FILLER_41_215 ();
 FILLCELL_X1 FILLER_41_217 ();
 FILLCELL_X2 FILLER_41_222 ();
 FILLCELL_X16 FILLER_41_227 ();
 FILLCELL_X2 FILLER_41_243 ();
 FILLCELL_X1 FILLER_41_245 ();
 FILLCELL_X1 FILLER_41_256 ();
 FILLCELL_X2 FILLER_41_273 ();
 FILLCELL_X1 FILLER_41_279 ();
 FILLCELL_X2 FILLER_41_308 ();
 FILLCELL_X1 FILLER_41_321 ();
 FILLCELL_X2 FILLER_41_343 ();
 FILLCELL_X4 FILLER_41_351 ();
 FILLCELL_X2 FILLER_41_355 ();
 FILLCELL_X1 FILLER_41_357 ();
 FILLCELL_X1 FILLER_41_361 ();
 FILLCELL_X1 FILLER_41_365 ();
 FILLCELL_X8 FILLER_42_1 ();
 FILLCELL_X4 FILLER_42_9 ();
 FILLCELL_X2 FILLER_42_16 ();
 FILLCELL_X1 FILLER_42_18 ();
 FILLCELL_X16 FILLER_42_45 ();
 FILLCELL_X8 FILLER_42_61 ();
 FILLCELL_X1 FILLER_42_69 ();
 FILLCELL_X16 FILLER_42_87 ();
 FILLCELL_X4 FILLER_42_103 ();
 FILLCELL_X1 FILLER_42_107 ();
 FILLCELL_X4 FILLER_42_112 ();
 FILLCELL_X1 FILLER_42_116 ();
 FILLCELL_X8 FILLER_42_121 ();
 FILLCELL_X1 FILLER_42_129 ();
 FILLCELL_X2 FILLER_42_133 ();
 FILLCELL_X8 FILLER_42_138 ();
 FILLCELL_X1 FILLER_42_146 ();
 FILLCELL_X4 FILLER_42_158 ();
 FILLCELL_X2 FILLER_42_162 ();
 FILLCELL_X1 FILLER_42_164 ();
 FILLCELL_X8 FILLER_42_182 ();
 FILLCELL_X2 FILLER_42_190 ();
 FILLCELL_X2 FILLER_42_201 ();
 FILLCELL_X8 FILLER_42_237 ();
 FILLCELL_X1 FILLER_42_252 ();
 FILLCELL_X4 FILLER_42_258 ();
 FILLCELL_X1 FILLER_42_262 ();
 FILLCELL_X2 FILLER_42_273 ();
 FILLCELL_X2 FILLER_42_279 ();
 FILLCELL_X1 FILLER_42_281 ();
 FILLCELL_X4 FILLER_42_327 ();
 FILLCELL_X2 FILLER_42_331 ();
 FILLCELL_X1 FILLER_42_333 ();
 FILLCELL_X16 FILLER_42_341 ();
 FILLCELL_X4 FILLER_42_357 ();
 FILLCELL_X1 FILLER_42_361 ();
 FILLCELL_X4 FILLER_42_365 ();
 FILLCELL_X2 FILLER_42_369 ();
 FILLCELL_X4 FILLER_42_377 ();
 FILLCELL_X2 FILLER_42_381 ();
 FILLCELL_X16 FILLER_43_1 ();
 FILLCELL_X8 FILLER_43_17 ();
 FILLCELL_X4 FILLER_43_25 ();
 FILLCELL_X1 FILLER_43_29 ();
 FILLCELL_X8 FILLER_43_33 ();
 FILLCELL_X4 FILLER_43_67 ();
 FILLCELL_X1 FILLER_43_71 ();
 FILLCELL_X4 FILLER_43_79 ();
 FILLCELL_X2 FILLER_43_83 ();
 FILLCELL_X1 FILLER_43_85 ();
 FILLCELL_X2 FILLER_43_103 ();
 FILLCELL_X1 FILLER_43_105 ();
 FILLCELL_X4 FILLER_43_128 ();
 FILLCELL_X4 FILLER_43_136 ();
 FILLCELL_X4 FILLER_43_142 ();
 FILLCELL_X2 FILLER_43_146 ();
 FILLCELL_X8 FILLER_43_150 ();
 FILLCELL_X2 FILLER_43_158 ();
 FILLCELL_X1 FILLER_43_160 ();
 FILLCELL_X8 FILLER_43_175 ();
 FILLCELL_X1 FILLER_43_183 ();
 FILLCELL_X4 FILLER_43_195 ();
 FILLCELL_X2 FILLER_43_199 ();
 FILLCELL_X1 FILLER_43_201 ();
 FILLCELL_X1 FILLER_43_210 ();
 FILLCELL_X4 FILLER_43_215 ();
 FILLCELL_X2 FILLER_43_219 ();
 FILLCELL_X1 FILLER_43_221 ();
 FILLCELL_X16 FILLER_43_230 ();
 FILLCELL_X1 FILLER_43_246 ();
 FILLCELL_X1 FILLER_43_257 ();
 FILLCELL_X2 FILLER_43_262 ();
 FILLCELL_X16 FILLER_43_283 ();
 FILLCELL_X8 FILLER_43_299 ();
 FILLCELL_X2 FILLER_43_307 ();
 FILLCELL_X4 FILLER_43_316 ();
 FILLCELL_X2 FILLER_43_320 ();
 FILLCELL_X32 FILLER_43_326 ();
 FILLCELL_X4 FILLER_43_358 ();
 FILLCELL_X1 FILLER_43_362 ();
 FILLCELL_X2 FILLER_43_366 ();
 FILLCELL_X2 FILLER_43_371 ();
 FILLCELL_X8 FILLER_43_376 ();
 FILLCELL_X2 FILLER_43_384 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X1 FILLER_44_9 ();
 FILLCELL_X4 FILLER_44_13 ();
 FILLCELL_X2 FILLER_44_17 ();
 FILLCELL_X1 FILLER_44_19 ();
 FILLCELL_X4 FILLER_44_46 ();
 FILLCELL_X1 FILLER_44_50 ();
 FILLCELL_X4 FILLER_44_70 ();
 FILLCELL_X8 FILLER_44_91 ();
 FILLCELL_X4 FILLER_44_99 ();
 FILLCELL_X2 FILLER_44_110 ();
 FILLCELL_X1 FILLER_44_112 ();
 FILLCELL_X1 FILLER_44_154 ();
 FILLCELL_X1 FILLER_44_166 ();
 FILLCELL_X2 FILLER_44_181 ();
 FILLCELL_X1 FILLER_44_205 ();
 FILLCELL_X2 FILLER_44_220 ();
 FILLCELL_X1 FILLER_44_226 ();
 FILLCELL_X8 FILLER_44_235 ();
 FILLCELL_X2 FILLER_44_243 ();
 FILLCELL_X1 FILLER_44_245 ();
 FILLCELL_X1 FILLER_44_275 ();
 FILLCELL_X16 FILLER_44_285 ();
 FILLCELL_X4 FILLER_44_301 ();
 FILLCELL_X2 FILLER_44_305 ();
 FILLCELL_X16 FILLER_44_324 ();
 FILLCELL_X8 FILLER_44_340 ();
 FILLCELL_X2 FILLER_44_348 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X1 FILLER_44_385 ();
 FILLCELL_X4 FILLER_45_1 ();
 FILLCELL_X2 FILLER_45_5 ();
 FILLCELL_X1 FILLER_45_7 ();
 FILLCELL_X8 FILLER_45_11 ();
 FILLCELL_X1 FILLER_45_26 ();
 FILLCELL_X1 FILLER_45_46 ();
 FILLCELL_X1 FILLER_45_73 ();
 FILLCELL_X8 FILLER_45_81 ();
 FILLCELL_X4 FILLER_45_89 ();
 FILLCELL_X1 FILLER_45_93 ();
 FILLCELL_X1 FILLER_45_111 ();
 FILLCELL_X2 FILLER_45_146 ();
 FILLCELL_X1 FILLER_45_154 ();
 FILLCELL_X2 FILLER_45_211 ();
 FILLCELL_X1 FILLER_45_213 ();
 FILLCELL_X1 FILLER_45_225 ();
 FILLCELL_X4 FILLER_45_273 ();
 FILLCELL_X1 FILLER_45_277 ();
 FILLCELL_X8 FILLER_45_310 ();
 FILLCELL_X4 FILLER_45_318 ();
 FILLCELL_X2 FILLER_45_322 ();
 FILLCELL_X32 FILLER_45_345 ();
 FILLCELL_X8 FILLER_45_377 ();
 FILLCELL_X1 FILLER_45_385 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X16 FILLER_46_33 ();
 FILLCELL_X4 FILLER_46_49 ();
 FILLCELL_X1 FILLER_46_53 ();
 FILLCELL_X8 FILLER_46_61 ();
 FILLCELL_X16 FILLER_46_93 ();
 FILLCELL_X1 FILLER_46_113 ();
 FILLCELL_X4 FILLER_46_160 ();
 FILLCELL_X1 FILLER_46_164 ();
 FILLCELL_X1 FILLER_46_191 ();
 FILLCELL_X4 FILLER_46_196 ();
 FILLCELL_X1 FILLER_46_200 ();
 FILLCELL_X2 FILLER_46_220 ();
 FILLCELL_X1 FILLER_46_239 ();
 FILLCELL_X32 FILLER_46_286 ();
 FILLCELL_X2 FILLER_46_318 ();
 FILLCELL_X32 FILLER_46_327 ();
 FILLCELL_X16 FILLER_46_359 ();
 FILLCELL_X8 FILLER_46_375 ();
 FILLCELL_X2 FILLER_46_383 ();
 FILLCELL_X1 FILLER_46_385 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X16 FILLER_47_33 ();
 FILLCELL_X8 FILLER_47_49 ();
 FILLCELL_X1 FILLER_47_57 ();
 FILLCELL_X1 FILLER_47_65 ();
 FILLCELL_X8 FILLER_47_83 ();
 FILLCELL_X4 FILLER_47_91 ();
 FILLCELL_X2 FILLER_47_95 ();
 FILLCELL_X1 FILLER_47_97 ();
 FILLCELL_X2 FILLER_47_122 ();
 FILLCELL_X1 FILLER_47_124 ();
 FILLCELL_X1 FILLER_47_132 ();
 FILLCELL_X1 FILLER_47_136 ();
 FILLCELL_X1 FILLER_47_140 ();
 FILLCELL_X1 FILLER_47_147 ();
 FILLCELL_X1 FILLER_47_159 ();
 FILLCELL_X2 FILLER_47_166 ();
 FILLCELL_X1 FILLER_47_181 ();
 FILLCELL_X4 FILLER_47_201 ();
 FILLCELL_X2 FILLER_47_205 ();
 FILLCELL_X2 FILLER_47_210 ();
 FILLCELL_X8 FILLER_47_237 ();
 FILLCELL_X2 FILLER_47_245 ();
 FILLCELL_X1 FILLER_47_247 ();
 FILLCELL_X1 FILLER_47_252 ();
 FILLCELL_X8 FILLER_47_275 ();
 FILLCELL_X1 FILLER_47_283 ();
 FILLCELL_X4 FILLER_47_301 ();
 FILLCELL_X2 FILLER_47_305 ();
 FILLCELL_X1 FILLER_47_307 ();
 FILLCELL_X32 FILLER_47_329 ();
 FILLCELL_X16 FILLER_47_361 ();
 FILLCELL_X8 FILLER_47_377 ();
 FILLCELL_X1 FILLER_47_385 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X2 FILLER_48_65 ();
 FILLCELL_X4 FILLER_48_91 ();
 FILLCELL_X16 FILLER_48_116 ();
 FILLCELL_X4 FILLER_48_132 ();
 FILLCELL_X1 FILLER_48_148 ();
 FILLCELL_X2 FILLER_48_154 ();
 FILLCELL_X8 FILLER_48_159 ();
 FILLCELL_X1 FILLER_48_167 ();
 FILLCELL_X1 FILLER_48_173 ();
 FILLCELL_X1 FILLER_48_178 ();
 FILLCELL_X2 FILLER_48_183 ();
 FILLCELL_X1 FILLER_48_202 ();
 FILLCELL_X4 FILLER_48_208 ();
 FILLCELL_X8 FILLER_48_235 ();
 FILLCELL_X2 FILLER_48_243 ();
 FILLCELL_X4 FILLER_48_258 ();
 FILLCELL_X2 FILLER_48_262 ();
 FILLCELL_X1 FILLER_48_264 ();
 FILLCELL_X1 FILLER_48_274 ();
 FILLCELL_X4 FILLER_48_289 ();
 FILLCELL_X2 FILLER_48_293 ();
 FILLCELL_X2 FILLER_48_299 ();
 FILLCELL_X1 FILLER_48_301 ();
 FILLCELL_X2 FILLER_48_316 ();
 FILLCELL_X1 FILLER_48_318 ();
 FILLCELL_X1 FILLER_48_322 ();
 FILLCELL_X32 FILLER_48_344 ();
 FILLCELL_X8 FILLER_48_376 ();
 FILLCELL_X2 FILLER_48_384 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X16 FILLER_49_33 ();
 FILLCELL_X8 FILLER_49_49 ();
 FILLCELL_X2 FILLER_49_57 ();
 FILLCELL_X1 FILLER_49_59 ();
 FILLCELL_X4 FILLER_49_67 ();
 FILLCELL_X4 FILLER_49_91 ();
 FILLCELL_X2 FILLER_49_95 ();
 FILLCELL_X1 FILLER_49_107 ();
 FILLCELL_X1 FILLER_49_129 ();
 FILLCELL_X1 FILLER_49_134 ();
 FILLCELL_X2 FILLER_49_139 ();
 FILLCELL_X1 FILLER_49_141 ();
 FILLCELL_X2 FILLER_49_148 ();
 FILLCELL_X4 FILLER_49_186 ();
 FILLCELL_X1 FILLER_49_190 ();
 FILLCELL_X4 FILLER_49_195 ();
 FILLCELL_X8 FILLER_49_203 ();
 FILLCELL_X4 FILLER_49_222 ();
 FILLCELL_X1 FILLER_49_226 ();
 FILLCELL_X4 FILLER_49_234 ();
 FILLCELL_X2 FILLER_49_238 ();
 FILLCELL_X1 FILLER_49_240 ();
 FILLCELL_X1 FILLER_49_245 ();
 FILLCELL_X4 FILLER_49_260 ();
 FILLCELL_X2 FILLER_49_264 ();
 FILLCELL_X4 FILLER_49_273 ();
 FILLCELL_X2 FILLER_49_277 ();
 FILLCELL_X8 FILLER_49_310 ();
 FILLCELL_X1 FILLER_49_318 ();
 FILLCELL_X32 FILLER_49_332 ();
 FILLCELL_X16 FILLER_49_364 ();
 FILLCELL_X4 FILLER_49_380 ();
 FILLCELL_X2 FILLER_49_384 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X8 FILLER_50_65 ();
 FILLCELL_X4 FILLER_50_73 ();
 FILLCELL_X2 FILLER_50_77 ();
 FILLCELL_X2 FILLER_50_109 ();
 FILLCELL_X2 FILLER_50_118 ();
 FILLCELL_X2 FILLER_50_154 ();
 FILLCELL_X1 FILLER_50_156 ();
 FILLCELL_X1 FILLER_50_172 ();
 FILLCELL_X1 FILLER_50_229 ();
 FILLCELL_X2 FILLER_50_296 ();
 FILLCELL_X2 FILLER_50_319 ();
 FILLCELL_X1 FILLER_50_342 ();
 FILLCELL_X32 FILLER_50_350 ();
 FILLCELL_X4 FILLER_50_382 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X8 FILLER_51_33 ();
 FILLCELL_X4 FILLER_51_41 ();
 FILLCELL_X2 FILLER_51_45 ();
 FILLCELL_X4 FILLER_51_50 ();
 FILLCELL_X1 FILLER_51_54 ();
 FILLCELL_X2 FILLER_51_64 ();
 FILLCELL_X1 FILLER_51_66 ();
 FILLCELL_X2 FILLER_51_92 ();
 FILLCELL_X1 FILLER_51_94 ();
 FILLCELL_X1 FILLER_51_107 ();
 FILLCELL_X2 FILLER_51_120 ();
 FILLCELL_X1 FILLER_51_122 ();
 FILLCELL_X1 FILLER_51_135 ();
 FILLCELL_X1 FILLER_51_145 ();
 FILLCELL_X1 FILLER_51_149 ();
 FILLCELL_X1 FILLER_51_153 ();
 FILLCELL_X1 FILLER_51_178 ();
 FILLCELL_X2 FILLER_51_206 ();
 FILLCELL_X1 FILLER_51_208 ();
 FILLCELL_X1 FILLER_51_218 ();
 FILLCELL_X1 FILLER_51_259 ();
 FILLCELL_X1 FILLER_51_269 ();
 FILLCELL_X1 FILLER_51_307 ();
 FILLCELL_X1 FILLER_51_317 ();
 FILLCELL_X1 FILLER_51_321 ();
 FILLCELL_X1 FILLER_51_341 ();
 FILLCELL_X32 FILLER_51_345 ();
 FILLCELL_X8 FILLER_51_377 ();
 FILLCELL_X1 FILLER_51_385 ();
endmodule
