module fixed_point_sqrt (clk,
    enable,
    reset,
    x,
    y);
 input clk;
 input enable;
 input reset;
 input [15:0] x;
 output [15:0] y;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__buf_2 _105_ (.A(enable),
    .X(_045_));
 sky130_fd_sc_hd__nor4_4 _106_ (.A(net6),
    .B(net5),
    .C(net7),
    .D(net8),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _107_ (.A(net15),
    .B(_045_),
    .Y(_047_));
 sky130_fd_sc_hd__a211oi_1 _108_ (.A1(_045_),
    .A2(_046_),
    .B1(_047_),
    .C1(net1),
    .Y(_000_));
 sky130_fd_sc_hd__buf_2 _109_ (.A(x[3]),
    .X(_048_));
 sky130_fd_sc_hd__nor3_1 _110_ (.A(net2),
    .B(_048_),
    .C(net10),
    .Y(_049_));
 sky130_fd_sc_hd__clkbuf_2 _111_ (.A(x[2]),
    .X(_050_));
 sky130_fd_sc_hd__buf_4 _112_ (.A(x[5]),
    .X(_051_));
 sky130_fd_sc_hd__nor3_1 _113_ (.A(net9),
    .B(_050_),
    .C(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__buf_4 _114_ (.A(x[6]),
    .X(_053_));
 sky130_fd_sc_hd__nor3_1 _115_ (.A(net11),
    .B(_053_),
    .C(net13),
    .Y(_054_));
 sky130_fd_sc_hd__nand3_2 _116_ (.A(_049_),
    .B(_052_),
    .C(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__buf_2 _117_ (.A(net12),
    .X(_056_));
 sky130_fd_sc_hd__nor2_1 _118_ (.A(net3),
    .B(net4),
    .Y(_057_));
 sky130_fd_sc_hd__nand3_1 _119_ (.A(_056_),
    .B(_046_),
    .C(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__o21a_1 _120_ (.A1(_055_),
    .A2(_058_),
    .B1(_045_),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _121_ (.A(_046_),
    .B(_057_),
    .Y(_060_));
 sky130_fd_sc_hd__nor4bb_1 _122_ (.A(_053_),
    .B(_056_),
    .C_N(net13),
    .D_N(net11),
    .Y(_061_));
 sky130_fd_sc_hd__nand3_1 _123_ (.A(_049_),
    .B(_052_),
    .C(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__nand4_1 _124_ (.A(net10),
    .B(net5),
    .C(net7),
    .D(net8),
    .Y(_063_));
 sky130_fd_sc_hd__nand4_1 _125_ (.A(_056_),
    .B(net3),
    .C(net4),
    .D(net6),
    .Y(_064_));
 sky130_fd_sc_hd__buf_4 _126_ (.A(net2),
    .X(_065_));
 sky130_fd_sc_hd__nand4_1 _127_ (.A(_065_),
    .B(net9),
    .C(_048_),
    .D(_053_),
    .Y(_066_));
 sky130_fd_sc_hd__nand4_1 _128_ (.A(_050_),
    .B(_051_),
    .C(net11),
    .D(net13),
    .Y(_067_));
 sky130_fd_sc_hd__or4_2 _129_ (.A(_063_),
    .B(_064_),
    .C(_066_),
    .D(_067_),
    .X(_068_));
 sky130_fd_sc_hd__o21ai_2 _130_ (.A1(_060_),
    .A2(_062_),
    .B1(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2b_1 _131_ (.A(_045_),
    .B_N(net17),
    .Y(_070_));
 sky130_fd_sc_hd__a21oi_1 _132_ (.A1(_059_),
    .A2(_069_),
    .B1(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__nor2_1 _133_ (.A(net1),
    .B(_071_),
    .Y(_001_));
 sky130_fd_sc_hd__nor4_1 _134_ (.A(_063_),
    .B(_064_),
    .C(_066_),
    .D(_067_),
    .Y(_072_));
 sky130_fd_sc_hd__nor2b_1 _135_ (.A(_045_),
    .B_N(net16),
    .Y(_073_));
 sky130_fd_sc_hd__a21oi_1 _136_ (.A1(_059_),
    .A2(_072_),
    .B1(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2_1 _137_ (.A(net1),
    .B(_074_),
    .Y(_002_));
 sky130_fd_sc_hd__nor2_1 _138_ (.A(_050_),
    .B(_051_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _139_ (.A(net13),
    .B(_056_),
    .Y(_076_));
 sky130_fd_sc_hd__nand3_2 _140_ (.A(_046_),
    .B(_057_),
    .C(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__nor4_1 _141_ (.A(net9),
    .B(net11),
    .C(_053_),
    .D(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__a41o_1 _142_ (.A1(_065_),
    .A2(_048_),
    .A3(_075_),
    .A4(_078_),
    .B1(_069_),
    .X(_079_));
 sky130_fd_sc_hd__nor2b_1 _143_ (.A(_045_),
    .B_N(net20),
    .Y(_080_));
 sky130_fd_sc_hd__a21oi_1 _144_ (.A1(_059_),
    .A2(_079_),
    .B1(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _145_ (.A(net1),
    .B(_081_),
    .Y(_003_));
 sky130_fd_sc_hd__nor2b_1 _146_ (.A(net1),
    .B_N(_059_),
    .Y(_082_));
 sky130_fd_sc_hd__nor3_1 _147_ (.A(net11),
    .B(_053_),
    .C(_077_),
    .Y(_083_));
 sky130_fd_sc_hd__nand2b_1 _148_ (.A_N(_048_),
    .B(net10),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(_065_),
    .B(_048_),
    .Y(_085_));
 sky130_fd_sc_hd__a21oi_1 _150_ (.A1(_065_),
    .A2(_084_),
    .B1(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__nor4bb_1 _151_ (.A(_048_),
    .B(net10),
    .C_N(_051_),
    .D_N(_050_),
    .Y(_087_));
 sky130_fd_sc_hd__nor4_1 _152_ (.A(_065_),
    .B(_048_),
    .C(_051_),
    .D(net10),
    .Y(_088_));
 sky130_fd_sc_hd__a21oi_1 _153_ (.A1(_065_),
    .A2(_087_),
    .B1(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__o31ai_1 _154_ (.A1(_050_),
    .A2(_051_),
    .A3(_086_),
    .B1(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__nor2_1 _155_ (.A(net9),
    .B(net11),
    .Y(_091_));
 sky130_fd_sc_hd__xnor2_1 _156_ (.A(_050_),
    .B(_051_),
    .Y(_092_));
 sky130_fd_sc_hd__nand4_1 _157_ (.A(_053_),
    .B(_049_),
    .C(_091_),
    .D(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__nor2_1 _158_ (.A(_077_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__nor2_1 _159_ (.A(_056_),
    .B(net6),
    .Y(_095_));
 sky130_fd_sc_hd__nand3_1 _160_ (.A(net5),
    .B(_057_),
    .C(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__nand2b_1 _161_ (.A_N(net4),
    .B(net3),
    .Y(_097_));
 sky130_fd_sc_hd__or4_1 _162_ (.A(net12),
    .B(net6),
    .C(net5),
    .D(_097_),
    .X(_098_));
 sky130_fd_sc_hd__and3b_1 _163_ (.A_N(net4),
    .B(net6),
    .C(net3),
    .X(_099_));
 sky130_fd_sc_hd__nor3b_1 _164_ (.A(net3),
    .B(net6),
    .C_N(net4),
    .Y(_100_));
 sky130_fd_sc_hd__nor2b_1 _165_ (.A(net5),
    .B_N(_056_),
    .Y(_101_));
 sky130_fd_sc_hd__o21ai_1 _166_ (.A1(_099_),
    .A2(_100_),
    .B1(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__or2_2 _167_ (.A(net7),
    .B(net8),
    .X(_103_));
 sky130_fd_sc_hd__a311oi_4 _168_ (.A1(_096_),
    .A2(_098_),
    .A3(_102_),
    .B1(_055_),
    .C1(_103_),
    .Y(_009_));
 sky130_fd_sc_hd__a211oi_2 _169_ (.A1(_078_),
    .A2(_090_),
    .B1(_094_),
    .C1(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__nand3_1 _170_ (.A(_082_),
    .B(_083_),
    .C(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _171_ (.A(_045_),
    .B(net1),
    .Y(_012_));
 sky130_fd_sc_hd__xor2_1 _172_ (.A(_065_),
    .B(_053_),
    .X(_013_));
 sky130_fd_sc_hd__nand3b_1 _173_ (.A_N(_050_),
    .B(_048_),
    .C(_065_),
    .Y(_014_));
 sky130_fd_sc_hd__or3b_1 _174_ (.A(_065_),
    .B(_048_),
    .C_N(_050_),
    .X(_015_));
 sky130_fd_sc_hd__or4_1 _175_ (.A(net9),
    .B(net10),
    .C(net11),
    .D(_053_),
    .X(_016_));
 sky130_fd_sc_hd__a211oi_1 _176_ (.A1(_014_),
    .A2(_015_),
    .B1(_051_),
    .C1(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__a31oi_1 _177_ (.A1(_087_),
    .A2(_091_),
    .A3(_013_),
    .B1(_017_),
    .Y(_018_));
 sky130_fd_sc_hd__o21ai_0 _178_ (.A1(_077_),
    .A2(_018_),
    .B1(_068_),
    .Y(_019_));
 sky130_fd_sc_hd__a22oi_1 _179_ (.A1(net21),
    .A2(_012_),
    .B1(_082_),
    .B2(_019_),
    .Y(_020_));
 sky130_fd_sc_hd__nand2_1 _180_ (.A(_011_),
    .B(_020_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2_1 _181_ (.A(_069_),
    .B(_009_),
    .Y(_021_));
 sky130_fd_sc_hd__a21boi_0 _182_ (.A1(_077_),
    .A2(_021_),
    .B1_N(_082_),
    .Y(_022_));
 sky130_fd_sc_hd__or2_0 _183_ (.A(_060_),
    .B(_062_),
    .X(_023_));
 sky130_fd_sc_hd__a31o_1 _184_ (.A1(_048_),
    .A2(net10),
    .A3(_075_),
    .B1(_087_),
    .X(_024_));
 sky130_fd_sc_hd__a32o_1 _185_ (.A1(net10),
    .A2(_075_),
    .A3(_085_),
    .B1(_024_),
    .B2(_065_),
    .X(_025_));
 sky130_fd_sc_hd__a221o_1 _186_ (.A1(_023_),
    .A2(_010_),
    .B1(_025_),
    .B2(_078_),
    .C1(_072_),
    .X(_026_));
 sky130_fd_sc_hd__a22o_1 _187_ (.A1(net22),
    .A2(_012_),
    .B1(_022_),
    .B2(_026_),
    .X(_005_));
 sky130_fd_sc_hd__nor2_1 _188_ (.A(net4),
    .B(net5),
    .Y(_027_));
 sky130_fd_sc_hd__o21ai_0 _189_ (.A1(net13),
    .A2(_056_),
    .B1(net3),
    .Y(_028_));
 sky130_fd_sc_hd__a21boi_1 _190_ (.A1(_027_),
    .A2(_028_),
    .B1_N(net6),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _191_ (.A(_069_),
    .B(_094_),
    .Y(_030_));
 sky130_fd_sc_hd__o41ai_1 _192_ (.A1(_103_),
    .A2(_083_),
    .A3(_009_),
    .A4(_029_),
    .B1(_030_),
    .Y(_031_));
 sky130_fd_sc_hd__a22o_1 _193_ (.A1(net23),
    .A2(_012_),
    .B1(_082_),
    .B2(_031_),
    .X(_006_));
 sky130_fd_sc_hd__nor2_1 _194_ (.A(_103_),
    .B(_055_),
    .Y(_032_));
 sky130_fd_sc_hd__o21bai_1 _195_ (.A1(net3),
    .A2(net6),
    .B1_N(_099_),
    .Y(_033_));
 sky130_fd_sc_hd__a31oi_1 _196_ (.A1(_101_),
    .A2(_032_),
    .A3(_033_),
    .B1(_069_),
    .Y(_034_));
 sky130_fd_sc_hd__or3_1 _197_ (.A(net13),
    .B(_056_),
    .C(net3),
    .X(_035_));
 sky130_fd_sc_hd__nand4_1 _198_ (.A(_046_),
    .B(_097_),
    .C(_010_),
    .D(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _199_ (.A(_045_),
    .B(net24),
    .Y(_037_));
 sky130_fd_sc_hd__a311oi_1 _200_ (.A1(_045_),
    .A2(_034_),
    .A3(_036_),
    .B1(_037_),
    .C1(net1),
    .Y(_007_));
 sky130_fd_sc_hd__o311a_1 _201_ (.A1(_103_),
    .A2(_046_),
    .A3(_029_),
    .B1(_068_),
    .C1(_060_),
    .X(_038_));
 sky130_fd_sc_hd__nand3_1 _202_ (.A(_082_),
    .B(_010_),
    .C(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__nand3b_1 _203_ (.A_N(net3),
    .B(net4),
    .C(_056_),
    .Y(_040_));
 sky130_fd_sc_hd__o21ai_0 _204_ (.A1(_056_),
    .A2(_097_),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_1 _205_ (.A(_046_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__o21ai_0 _206_ (.A1(_055_),
    .A2(_042_),
    .B1(_068_),
    .Y(_043_));
 sky130_fd_sc_hd__a22oi_1 _207_ (.A1(net25),
    .A2(_012_),
    .B1(_082_),
    .B2(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _208_ (.A(_039_),
    .B(_044_),
    .Y(_008_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _210_ (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(net16),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 _212_ (.A(net16),
    .X(net19));
 sky130_fd_sc_hd__buf_4 _213_ (.A(net26),
    .X(y[12]));
 sky130_fd_sc_hd__buf_4 _214_ (.A(net27),
    .X(y[13]));
 sky130_fd_sc_hd__buf_4 _215_ (.A(net28),
    .X(y[14]));
 sky130_fd_sc_hd__buf_4 _216_ (.A(net29),
    .X(y[15]));
 sky130_fd_sc_hd__dfxtp_1 \y[10]$_SDFFE_PP0P_  (.D(_000_),
    .Q(net15),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[1]$_SDFFE_PP0P_  (.D(_001_),
    .Q(net17),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[3]$_SDFFE_PP0P_  (.D(_002_),
    .Q(net16),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[4]$_SDFFE_PP0P_  (.D(_003_),
    .Q(net20),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[5]$_SDFFE_PP0P_  (.D(_004_),
    .Q(net21),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[6]$_SDFFE_PP0P_  (.D(_005_),
    .Q(net22),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[7]$_SDFFE_PP0P_  (.D(_006_),
    .Q(net23),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[8]$_SDFFE_PP0P_  (.D(_007_),
    .Q(net24),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \y[9]$_SDFFE_PP0P_  (.D(_008_),
    .Q(net25),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_74 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(reset),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(x[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(x[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(x[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(x[12]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(x[13]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(x[14]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(x[15]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(x[1]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(x[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(x[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(x[8]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(x[9]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(y[0]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(y[10]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(y[11]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(y[1]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(y[2]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(y[3]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(y[4]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(y[5]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(y[6]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(y[7]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(y[8]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(y[9]));
 sky130_fd_sc_hd__conb_1 _213__26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 _214__27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 _215__28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 _216__29 (.LO(net29));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_167 ();
endmodule
