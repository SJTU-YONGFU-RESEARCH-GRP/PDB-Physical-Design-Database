module ddr_controller (clk,
    cmd_ready,
    cmd_valid,
    cmd_write,
    init_done,
    phy_cas_n,
    phy_cke,
    phy_clk,
    phy_cs_n,
    phy_odt,
    phy_ras_n,
    phy_reset_n,
    phy_we_n,
    rd_ready,
    rd_valid,
    rst_n,
    wr_ready,
    wr_valid,
    cmd_addr,
    cmd_burst_len,
    phy_addr,
    phy_bank,
    phy_bank_group,
    phy_dm,
    phy_dq,
    phy_dqs_n,
    phy_dqs_p,
    rd_data,
    state,
    wr_data,
    wr_mask);
 input clk;
 output cmd_ready;
 input cmd_valid;
 input cmd_write;
 output init_done;
 output phy_cas_n;
 output phy_cke;
 input phy_clk;
 output phy_cs_n;
 output phy_odt;
 output phy_ras_n;
 output phy_reset_n;
 output phy_we_n;
 input rd_ready;
 output rd_valid;
 input rst_n;
 output wr_ready;
 input wr_valid;
 input [27:0] cmd_addr;
 input [3:0] cmd_burst_len;
 output [13:0] phy_addr;
 output [2:0] phy_bank;
 output [1:0] phy_bank_group;
 output [7:0] phy_dm;
 inout [63:0] phy_dq;
 inout [7:0] phy_dqs_n;
 inout [7:0] phy_dqs_p;
 output [63:0] rd_data;
 output [1:0] state;
 input [63:0] wr_data;
 input [7:0] wr_mask;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire clknet_0_clk;
 wire net209;
 wire \active_row[0][0] ;
 wire \active_row[0][10] ;
 wire \active_row[0][11] ;
 wire \active_row[0][12] ;
 wire \active_row[0][13] ;
 wire \active_row[0][1] ;
 wire \active_row[0][2] ;
 wire \active_row[0][3] ;
 wire \active_row[0][4] ;
 wire \active_row[0][5] ;
 wire \active_row[0][6] ;
 wire \active_row[0][7] ;
 wire \active_row[0][8] ;
 wire \active_row[0][9] ;
 wire \active_row[1][0] ;
 wire \active_row[1][10] ;
 wire \active_row[1][11] ;
 wire \active_row[1][12] ;
 wire \active_row[1][13] ;
 wire \active_row[1][1] ;
 wire \active_row[1][2] ;
 wire \active_row[1][3] ;
 wire \active_row[1][4] ;
 wire \active_row[1][5] ;
 wire \active_row[1][6] ;
 wire \active_row[1][7] ;
 wire \active_row[1][8] ;
 wire \active_row[1][9] ;
 wire \active_row[2][0] ;
 wire \active_row[2][10] ;
 wire \active_row[2][11] ;
 wire \active_row[2][12] ;
 wire \active_row[2][13] ;
 wire \active_row[2][1] ;
 wire \active_row[2][2] ;
 wire \active_row[2][3] ;
 wire \active_row[2][4] ;
 wire \active_row[2][5] ;
 wire \active_row[2][6] ;
 wire \active_row[2][7] ;
 wire \active_row[2][8] ;
 wire \active_row[2][9] ;
 wire \active_row[3][0] ;
 wire \active_row[3][10] ;
 wire \active_row[3][11] ;
 wire \active_row[3][12] ;
 wire \active_row[3][13] ;
 wire \active_row[3][1] ;
 wire \active_row[3][2] ;
 wire \active_row[3][3] ;
 wire \active_row[3][4] ;
 wire \active_row[3][5] ;
 wire \active_row[3][6] ;
 wire \active_row[3][7] ;
 wire \active_row[3][8] ;
 wire \active_row[3][9] ;
 wire \active_row[4][0] ;
 wire \active_row[4][10] ;
 wire \active_row[4][11] ;
 wire \active_row[4][12] ;
 wire \active_row[4][13] ;
 wire \active_row[4][1] ;
 wire \active_row[4][2] ;
 wire \active_row[4][3] ;
 wire \active_row[4][4] ;
 wire \active_row[4][5] ;
 wire \active_row[4][6] ;
 wire \active_row[4][7] ;
 wire \active_row[4][8] ;
 wire \active_row[4][9] ;
 wire \active_row[5][0] ;
 wire \active_row[5][10] ;
 wire \active_row[5][11] ;
 wire \active_row[5][12] ;
 wire \active_row[5][13] ;
 wire \active_row[5][1] ;
 wire \active_row[5][2] ;
 wire \active_row[5][3] ;
 wire \active_row[5][4] ;
 wire \active_row[5][5] ;
 wire \active_row[5][6] ;
 wire \active_row[5][7] ;
 wire \active_row[5][8] ;
 wire \active_row[5][9] ;
 wire \active_row[6][0] ;
 wire \active_row[6][10] ;
 wire \active_row[6][11] ;
 wire \active_row[6][12] ;
 wire \active_row[6][13] ;
 wire \active_row[6][1] ;
 wire \active_row[6][2] ;
 wire \active_row[6][3] ;
 wire \active_row[6][4] ;
 wire \active_row[6][5] ;
 wire \active_row[6][6] ;
 wire \active_row[6][7] ;
 wire \active_row[6][8] ;
 wire \active_row[6][9] ;
 wire \active_row[7][0] ;
 wire \active_row[7][10] ;
 wire \active_row[7][11] ;
 wire \active_row[7][12] ;
 wire \active_row[7][13] ;
 wire \active_row[7][1] ;
 wire \active_row[7][2] ;
 wire \active_row[7][3] ;
 wire \active_row[7][4] ;
 wire \active_row[7][5] ;
 wire \active_row[7][6] ;
 wire \active_row[7][7] ;
 wire \active_row[7][8] ;
 wire \active_row[7][9] ;
 wire \bank_active[0] ;
 wire \bank_active[1] ;
 wire \bank_active[2] ;
 wire \bank_active[3] ;
 wire \bank_active[4] ;
 wire \bank_active[5] ;
 wire \bank_active[6] ;
 wire \bank_active[7] ;
 wire \burst_counter[0] ;
 wire \burst_counter[1] ;
 wire \burst_counter[2] ;
 wire \burst_counter[3] ;
 wire cmd_reg_valid;
 wire \init_state[0] ;
 wire \init_state[1] ;
 wire \init_state[2] ;
 wire \init_state[3] ;
 wire \init_state[4] ;
 wire \init_state[5] ;
 wire \init_state[6] ;
 wire \init_state[7] ;
 wire \refresh_counter[0] ;
 wire \refresh_counter[10] ;
 wire \refresh_counter[11] ;
 wire \refresh_counter[12] ;
 wire \refresh_counter[13] ;
 wire \refresh_counter[14] ;
 wire \refresh_counter[15] ;
 wire \refresh_counter[1] ;
 wire \refresh_counter[2] ;
 wire \refresh_counter[3] ;
 wire \refresh_counter[4] ;
 wire \refresh_counter[5] ;
 wire \refresh_counter[6] ;
 wire \refresh_counter[7] ;
 wire \refresh_counter[8] ;
 wire \refresh_counter[9] ;
 wire \timer[0] ;
 wire \timer[10] ;
 wire \timer[11] ;
 wire \timer[12] ;
 wire \timer[13] ;
 wire \timer[14] ;
 wire \timer[15] ;
 wire \timer[1] ;
 wire \timer[2] ;
 wire \timer[3] ;
 wire \timer[4] ;
 wire \timer[5] ;
 wire \timer[6] ;
 wire \timer[7] ;
 wire \timer[8] ;
 wire \timer[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 BUF_X4 _1192_ (.A(net33),
    .Z(_0801_));
 CLKBUF_X3 _1193_ (.A(_0801_),
    .Z(_0802_));
 BUF_X2 _1194_ (.A(_0802_),
    .Z(_0803_));
 CLKBUF_X2 _1195_ (.A(_1182_),
    .Z(_0804_));
 INV_X1 _1196_ (.A(_0804_),
    .ZN(_0805_));
 BUF_X4 _1197_ (.A(_0805_),
    .Z(_0806_));
 CLKBUF_X2 _1198_ (.A(_1176_),
    .Z(_0807_));
 BUF_X1 _1199_ (.A(\timer[3] ),
    .Z(_0808_));
 NOR2_X2 _1200_ (.A1(\timer[2] ),
    .A2(_0808_),
    .ZN(_0809_));
 NAND2_X4 _1201_ (.A1(_0807_),
    .A2(_0809_),
    .ZN(_0810_));
 OR3_X2 _1202_ (.A1(\timer[11] ),
    .A2(\timer[10] ),
    .A3(\timer[12] ),
    .ZN(_0811_));
 OR3_X1 _1203_ (.A1(\timer[13] ),
    .A2(\timer[14] ),
    .A3(\timer[15] ),
    .ZN(_0812_));
 OR3_X1 _1204_ (.A1(\timer[7] ),
    .A2(\timer[6] ),
    .A3(\timer[8] ),
    .ZN(_0813_));
 OR3_X1 _1205_ (.A1(\timer[5] ),
    .A2(\timer[4] ),
    .A3(\timer[9] ),
    .ZN(_0814_));
 OR4_X1 _1206_ (.A1(_0811_),
    .A2(_0812_),
    .A3(_0813_),
    .A4(_0814_),
    .ZN(_0815_));
 BUF_X4 _1207_ (.A(_0815_),
    .Z(_0816_));
 NOR2_X4 _1208_ (.A1(_0810_),
    .A2(_0816_),
    .ZN(_0817_));
 INV_X1 _1209_ (.A(_0817_),
    .ZN(_0818_));
 BUF_X4 _1210_ (.A(_0818_),
    .Z(_0819_));
 BUF_X4 _1211_ (.A(_0819_),
    .Z(_0820_));
 NOR2_X4 _1212_ (.A1(_0806_),
    .A2(_0820_),
    .ZN(_0821_));
 MUX2_X1 _1213_ (.A(\init_state[2] ),
    .B(\init_state[4] ),
    .S(_0821_),
    .Z(_0822_));
 AND2_X1 _1214_ (.A1(_0803_),
    .A2(_0822_),
    .ZN(_0002_));
 BUF_X1 _1215_ (.A(\init_state[3] ),
    .Z(_0823_));
 CLKBUF_X3 _1216_ (.A(\init_state[5] ),
    .Z(_0824_));
 MUX2_X1 _1217_ (.A(_0823_),
    .B(_0824_),
    .S(_0821_),
    .Z(_0825_));
 AND2_X1 _1218_ (.A1(_0803_),
    .A2(_0825_),
    .ZN(_0003_));
 BUF_X1 _1219_ (.A(\init_state[0] ),
    .Z(_0826_));
 MUX2_X1 _1220_ (.A(\init_state[4] ),
    .B(_0826_),
    .S(_0821_),
    .Z(_0827_));
 AND2_X1 _1221_ (.A1(_0803_),
    .A2(_0827_),
    .ZN(_0004_));
 CLKBUF_X3 _1222_ (.A(\init_state[1] ),
    .Z(_0828_));
 MUX2_X1 _1223_ (.A(_0824_),
    .B(_0828_),
    .S(_0821_),
    .Z(_0829_));
 AND2_X1 _1224_ (.A1(_0803_),
    .A2(_0829_),
    .ZN(_0005_));
 MUX2_X1 _1225_ (.A(\init_state[6] ),
    .B(\init_state[2] ),
    .S(_0821_),
    .Z(_0830_));
 AND2_X1 _1226_ (.A1(_0803_),
    .A2(_0830_),
    .ZN(_0006_));
 INV_X1 _1227_ (.A(_0826_),
    .ZN(_0831_));
 OAI21_X1 _1228_ (.A(_0803_),
    .B1(_0831_),
    .B2(_0821_),
    .ZN(_0000_));
 MUX2_X1 _1229_ (.A(_0828_),
    .B(\init_state[6] ),
    .S(_0821_),
    .Z(_0832_));
 AND2_X1 _1230_ (.A1(_0803_),
    .A2(_0832_),
    .ZN(_0001_));
 INV_X4 _1231_ (.A(_0801_),
    .ZN(_0833_));
 CLKBUF_X3 _1232_ (.A(_0833_),
    .Z(_0834_));
 CLKBUF_X3 _1233_ (.A(_0834_),
    .Z(_0835_));
 BUF_X1 _1234_ (.A(\init_state[7] ),
    .Z(_0836_));
 AOI21_X1 _1235_ (.A(_0836_),
    .B1(_0821_),
    .B2(_0823_),
    .ZN(_0837_));
 NOR2_X1 _1236_ (.A1(_0835_),
    .A2(_0837_),
    .ZN(_0007_));
 OR2_X1 _1237_ (.A1(\refresh_counter[13] ),
    .A2(\refresh_counter[12] ),
    .ZN(_0838_));
 OR4_X2 _1238_ (.A1(\refresh_counter[15] ),
    .A2(\refresh_counter[14] ),
    .A3(\refresh_counter[11] ),
    .A4(_0838_),
    .ZN(_0839_));
 BUF_X1 _1239_ (.A(\refresh_counter[5] ),
    .Z(_0840_));
 NOR2_X1 _1240_ (.A1(\refresh_counter[6] ),
    .A2(_0840_),
    .ZN(_0841_));
 NAND3_X1 _1241_ (.A1(\refresh_counter[3] ),
    .A2(\refresh_counter[2] ),
    .A3(\refresh_counter[4] ),
    .ZN(_0842_));
 NOR2_X1 _1242_ (.A1(_1167_),
    .A2(_1165_),
    .ZN(_0843_));
 OAI21_X2 _1243_ (.A(_0841_),
    .B1(_0842_),
    .B2(_0843_),
    .ZN(_0844_));
 AND4_X1 _1244_ (.A1(\refresh_counter[7] ),
    .A2(\refresh_counter[10] ),
    .A3(\refresh_counter[9] ),
    .A4(\refresh_counter[8] ),
    .ZN(_0845_));
 AOI21_X4 _1245_ (.A(_0839_),
    .B1(_0844_),
    .B2(_0845_),
    .ZN(_1162_));
 BUF_X4 _1246_ (.A(_0820_),
    .Z(_1170_));
 BUF_X2 _1247_ (.A(net101),
    .Z(_0846_));
 BUF_X4 _1248_ (.A(net117),
    .Z(_0847_));
 INV_X4 _1249_ (.A(_0847_),
    .ZN(_0848_));
 INV_X2 _1250_ (.A(net115),
    .ZN(_0849_));
 BUF_X4 _1251_ (.A(_1184_),
    .Z(_0850_));
 INV_X4 _1252_ (.A(_0850_),
    .ZN(_0851_));
 BUF_X2 _1253_ (.A(net116),
    .Z(_0852_));
 NOR4_X4 _1254_ (.A1(_0833_),
    .A2(_0851_),
    .A3(_0852_),
    .A4(_0819_),
    .ZN(_0853_));
 NAND3_X4 _1255_ (.A1(_0848_),
    .A2(_0849_),
    .A3(_0853_),
    .ZN(_0854_));
 BUF_X4 _1256_ (.A(_0854_),
    .Z(_0855_));
 MUX2_X1 _1257_ (.A(_0846_),
    .B(\active_row[0][0] ),
    .S(_0855_),
    .Z(_0046_));
 BUF_X2 _1258_ (.A(net102),
    .Z(_0856_));
 MUX2_X1 _1259_ (.A(_0856_),
    .B(\active_row[0][10] ),
    .S(_0855_),
    .Z(_0047_));
 BUF_X2 _1260_ (.A(net103),
    .Z(_0857_));
 MUX2_X1 _1261_ (.A(_0857_),
    .B(\active_row[0][11] ),
    .S(_0855_),
    .Z(_0048_));
 BUF_X2 _1262_ (.A(net104),
    .Z(_0858_));
 MUX2_X1 _1263_ (.A(_0858_),
    .B(\active_row[0][12] ),
    .S(_0855_),
    .Z(_0049_));
 BUF_X2 _1264_ (.A(net105),
    .Z(_0859_));
 MUX2_X1 _1265_ (.A(_0859_),
    .B(\active_row[0][13] ),
    .S(_0855_),
    .Z(_0050_));
 BUF_X2 _1266_ (.A(net106),
    .Z(_0860_));
 MUX2_X1 _1267_ (.A(_0860_),
    .B(\active_row[0][1] ),
    .S(_0855_),
    .Z(_0051_));
 BUF_X2 _1268_ (.A(net107),
    .Z(_0861_));
 MUX2_X1 _1269_ (.A(_0861_),
    .B(\active_row[0][2] ),
    .S(_0855_),
    .Z(_0052_));
 CLKBUF_X2 _1270_ (.A(net108),
    .Z(_0862_));
 MUX2_X1 _1271_ (.A(_0862_),
    .B(\active_row[0][3] ),
    .S(_0855_),
    .Z(_0053_));
 BUF_X2 _1272_ (.A(net109),
    .Z(_0863_));
 MUX2_X1 _1273_ (.A(_0863_),
    .B(\active_row[0][4] ),
    .S(_0855_),
    .Z(_0054_));
 BUF_X2 _1274_ (.A(net110),
    .Z(_0864_));
 MUX2_X1 _1275_ (.A(_0864_),
    .B(\active_row[0][5] ),
    .S(_0855_),
    .Z(_0055_));
 BUF_X2 _1276_ (.A(net111),
    .Z(_0865_));
 MUX2_X1 _1277_ (.A(_0865_),
    .B(\active_row[0][6] ),
    .S(_0854_),
    .Z(_0056_));
 BUF_X2 _1278_ (.A(net112),
    .Z(_0866_));
 MUX2_X1 _1279_ (.A(_0866_),
    .B(\active_row[0][7] ),
    .S(_0854_),
    .Z(_0057_));
 BUF_X2 _1280_ (.A(net113),
    .Z(_0867_));
 MUX2_X1 _1281_ (.A(_0867_),
    .B(\active_row[0][8] ),
    .S(_0854_),
    .Z(_0058_));
 CLKBUF_X2 _1282_ (.A(net114),
    .Z(_0868_));
 MUX2_X1 _1283_ (.A(_0868_),
    .B(\active_row[0][9] ),
    .S(_0854_),
    .Z(_0059_));
 INV_X4 _1284_ (.A(_1145_),
    .ZN(_0869_));
 NAND3_X4 _1285_ (.A1(_0848_),
    .A2(_0869_),
    .A3(_0853_),
    .ZN(_0870_));
 BUF_X4 _1286_ (.A(_0870_),
    .Z(_0871_));
 MUX2_X1 _1287_ (.A(_0846_),
    .B(\active_row[1][0] ),
    .S(_0871_),
    .Z(_0060_));
 MUX2_X1 _1288_ (.A(_0856_),
    .B(\active_row[1][10] ),
    .S(_0871_),
    .Z(_0061_));
 MUX2_X1 _1289_ (.A(_0857_),
    .B(\active_row[1][11] ),
    .S(_0871_),
    .Z(_0062_));
 MUX2_X1 _1290_ (.A(_0858_),
    .B(\active_row[1][12] ),
    .S(_0871_),
    .Z(_0063_));
 MUX2_X1 _1291_ (.A(_0859_),
    .B(\active_row[1][13] ),
    .S(_0871_),
    .Z(_0064_));
 MUX2_X1 _1292_ (.A(_0860_),
    .B(\active_row[1][1] ),
    .S(_0871_),
    .Z(_0065_));
 MUX2_X1 _1293_ (.A(_0861_),
    .B(\active_row[1][2] ),
    .S(_0871_),
    .Z(_0066_));
 MUX2_X1 _1294_ (.A(_0862_),
    .B(\active_row[1][3] ),
    .S(_0871_),
    .Z(_0067_));
 MUX2_X1 _1295_ (.A(_0863_),
    .B(\active_row[1][4] ),
    .S(_0871_),
    .Z(_0068_));
 MUX2_X1 _1296_ (.A(_0864_),
    .B(\active_row[1][5] ),
    .S(_0871_),
    .Z(_0069_));
 MUX2_X1 _1297_ (.A(_0865_),
    .B(\active_row[1][6] ),
    .S(_0870_),
    .Z(_0070_));
 MUX2_X1 _1298_ (.A(_0866_),
    .B(\active_row[1][7] ),
    .S(_0870_),
    .Z(_0071_));
 MUX2_X1 _1299_ (.A(_0867_),
    .B(\active_row[1][8] ),
    .S(_0870_),
    .Z(_0072_));
 MUX2_X1 _1300_ (.A(_0868_),
    .B(\active_row[1][9] ),
    .S(_0870_),
    .Z(_0073_));
 BUF_X4 _1301_ (.A(_0817_),
    .Z(_0872_));
 NAND4_X4 _1302_ (.A1(_0801_),
    .A2(_0850_),
    .A3(_0852_),
    .A4(_0872_),
    .ZN(_0873_));
 NOR3_X4 _1303_ (.A1(_0847_),
    .A2(_0869_),
    .A3(_0873_),
    .ZN(_0874_));
 BUF_X4 _1304_ (.A(_0874_),
    .Z(_0875_));
 MUX2_X1 _1305_ (.A(\active_row[2][0] ),
    .B(_0846_),
    .S(_0875_),
    .Z(_0074_));
 MUX2_X1 _1306_ (.A(\active_row[2][10] ),
    .B(_0856_),
    .S(_0875_),
    .Z(_0075_));
 MUX2_X1 _1307_ (.A(\active_row[2][11] ),
    .B(_0857_),
    .S(_0875_),
    .Z(_0076_));
 MUX2_X1 _1308_ (.A(\active_row[2][12] ),
    .B(_0858_),
    .S(_0875_),
    .Z(_0077_));
 MUX2_X1 _1309_ (.A(\active_row[2][13] ),
    .B(_0859_),
    .S(_0875_),
    .Z(_0078_));
 MUX2_X1 _1310_ (.A(\active_row[2][1] ),
    .B(_0860_),
    .S(_0875_),
    .Z(_0079_));
 MUX2_X1 _1311_ (.A(\active_row[2][2] ),
    .B(_0861_),
    .S(_0875_),
    .Z(_0080_));
 MUX2_X1 _1312_ (.A(\active_row[2][3] ),
    .B(_0862_),
    .S(_0875_),
    .Z(_0081_));
 MUX2_X1 _1313_ (.A(\active_row[2][4] ),
    .B(_0863_),
    .S(_0875_),
    .Z(_0082_));
 MUX2_X1 _1314_ (.A(\active_row[2][5] ),
    .B(_0864_),
    .S(_0875_),
    .Z(_0083_));
 MUX2_X1 _1315_ (.A(\active_row[2][6] ),
    .B(_0865_),
    .S(_0874_),
    .Z(_0084_));
 MUX2_X1 _1316_ (.A(\active_row[2][7] ),
    .B(_0866_),
    .S(_0874_),
    .Z(_0085_));
 MUX2_X1 _1317_ (.A(\active_row[2][8] ),
    .B(_0867_),
    .S(_0874_),
    .Z(_0086_));
 MUX2_X1 _1318_ (.A(\active_row[2][9] ),
    .B(_0868_),
    .S(_0874_),
    .Z(_0087_));
 OR3_X4 _1319_ (.A1(_0847_),
    .A2(_1145_),
    .A3(_0873_),
    .ZN(_0876_));
 BUF_X4 _1320_ (.A(_0876_),
    .Z(_0877_));
 MUX2_X1 _1321_ (.A(_0846_),
    .B(\active_row[3][0] ),
    .S(_0877_),
    .Z(_0088_));
 MUX2_X1 _1322_ (.A(_0856_),
    .B(\active_row[3][10] ),
    .S(_0877_),
    .Z(_0089_));
 MUX2_X1 _1323_ (.A(_0857_),
    .B(\active_row[3][11] ),
    .S(_0877_),
    .Z(_0090_));
 MUX2_X1 _1324_ (.A(_0858_),
    .B(\active_row[3][12] ),
    .S(_0877_),
    .Z(_0091_));
 MUX2_X1 _1325_ (.A(_0859_),
    .B(\active_row[3][13] ),
    .S(_0877_),
    .Z(_0092_));
 MUX2_X1 _1326_ (.A(_0860_),
    .B(\active_row[3][1] ),
    .S(_0877_),
    .Z(_0093_));
 MUX2_X1 _1327_ (.A(_0861_),
    .B(\active_row[3][2] ),
    .S(_0877_),
    .Z(_0094_));
 MUX2_X1 _1328_ (.A(_0862_),
    .B(\active_row[3][3] ),
    .S(_0877_),
    .Z(_0095_));
 MUX2_X1 _1329_ (.A(_0863_),
    .B(\active_row[3][4] ),
    .S(_0877_),
    .Z(_0096_));
 MUX2_X1 _1330_ (.A(_0864_),
    .B(\active_row[3][5] ),
    .S(_0877_),
    .Z(_0097_));
 MUX2_X1 _1331_ (.A(_0865_),
    .B(\active_row[3][6] ),
    .S(_0876_),
    .Z(_0098_));
 MUX2_X1 _1332_ (.A(_0866_),
    .B(\active_row[3][7] ),
    .S(_0876_),
    .Z(_0099_));
 MUX2_X1 _1333_ (.A(_0867_),
    .B(\active_row[3][8] ),
    .S(_0876_),
    .Z(_0100_));
 MUX2_X1 _1334_ (.A(_0868_),
    .B(\active_row[3][9] ),
    .S(_0876_),
    .Z(_0101_));
 NAND3_X4 _1335_ (.A1(_0847_),
    .A2(_0849_),
    .A3(_0853_),
    .ZN(_0878_));
 BUF_X4 _1336_ (.A(_0878_),
    .Z(_0879_));
 MUX2_X1 _1337_ (.A(_0846_),
    .B(\active_row[4][0] ),
    .S(_0879_),
    .Z(_0102_));
 MUX2_X1 _1338_ (.A(_0856_),
    .B(\active_row[4][10] ),
    .S(_0879_),
    .Z(_0103_));
 MUX2_X1 _1339_ (.A(_0857_),
    .B(\active_row[4][11] ),
    .S(_0879_),
    .Z(_0104_));
 MUX2_X1 _1340_ (.A(_0858_),
    .B(\active_row[4][12] ),
    .S(_0879_),
    .Z(_0105_));
 MUX2_X1 _1341_ (.A(_0859_),
    .B(\active_row[4][13] ),
    .S(_0879_),
    .Z(_0106_));
 MUX2_X1 _1342_ (.A(_0860_),
    .B(\active_row[4][1] ),
    .S(_0879_),
    .Z(_0107_));
 MUX2_X1 _1343_ (.A(_0861_),
    .B(\active_row[4][2] ),
    .S(_0879_),
    .Z(_0108_));
 MUX2_X1 _1344_ (.A(_0862_),
    .B(\active_row[4][3] ),
    .S(_0879_),
    .Z(_0109_));
 MUX2_X1 _1345_ (.A(_0863_),
    .B(\active_row[4][4] ),
    .S(_0879_),
    .Z(_0110_));
 MUX2_X1 _1346_ (.A(_0864_),
    .B(\active_row[4][5] ),
    .S(_0879_),
    .Z(_0111_));
 MUX2_X1 _1347_ (.A(_0865_),
    .B(\active_row[4][6] ),
    .S(_0878_),
    .Z(_0112_));
 MUX2_X1 _1348_ (.A(_0866_),
    .B(\active_row[4][7] ),
    .S(_0878_),
    .Z(_0113_));
 MUX2_X1 _1349_ (.A(_0867_),
    .B(\active_row[4][8] ),
    .S(_0878_),
    .Z(_0114_));
 MUX2_X1 _1350_ (.A(_0868_),
    .B(\active_row[4][9] ),
    .S(_0878_),
    .Z(_0115_));
 NAND3_X4 _1351_ (.A1(_0847_),
    .A2(_0869_),
    .A3(_0853_),
    .ZN(_0880_));
 BUF_X4 _1352_ (.A(_0880_),
    .Z(_0881_));
 MUX2_X1 _1353_ (.A(_0846_),
    .B(\active_row[5][0] ),
    .S(_0881_),
    .Z(_0116_));
 MUX2_X1 _1354_ (.A(_0856_),
    .B(\active_row[5][10] ),
    .S(_0881_),
    .Z(_0117_));
 MUX2_X1 _1355_ (.A(_0857_),
    .B(\active_row[5][11] ),
    .S(_0881_),
    .Z(_0118_));
 MUX2_X1 _1356_ (.A(_0858_),
    .B(\active_row[5][12] ),
    .S(_0881_),
    .Z(_0119_));
 MUX2_X1 _1357_ (.A(_0859_),
    .B(\active_row[5][13] ),
    .S(_0881_),
    .Z(_0120_));
 MUX2_X1 _1358_ (.A(_0860_),
    .B(\active_row[5][1] ),
    .S(_0881_),
    .Z(_0121_));
 MUX2_X1 _1359_ (.A(_0861_),
    .B(\active_row[5][2] ),
    .S(_0881_),
    .Z(_0122_));
 MUX2_X1 _1360_ (.A(_0862_),
    .B(\active_row[5][3] ),
    .S(_0881_),
    .Z(_0123_));
 MUX2_X1 _1361_ (.A(_0863_),
    .B(\active_row[5][4] ),
    .S(_0881_),
    .Z(_0124_));
 MUX2_X1 _1362_ (.A(_0864_),
    .B(\active_row[5][5] ),
    .S(_0881_),
    .Z(_0125_));
 MUX2_X1 _1363_ (.A(_0865_),
    .B(\active_row[5][6] ),
    .S(_0880_),
    .Z(_0126_));
 MUX2_X1 _1364_ (.A(_0866_),
    .B(\active_row[5][7] ),
    .S(_0880_),
    .Z(_0127_));
 MUX2_X1 _1365_ (.A(_0867_),
    .B(\active_row[5][8] ),
    .S(_0880_),
    .Z(_0128_));
 MUX2_X1 _1366_ (.A(_0868_),
    .B(\active_row[5][9] ),
    .S(_0880_),
    .Z(_0129_));
 NOR3_X4 _1367_ (.A1(_0848_),
    .A2(net115),
    .A3(_0873_),
    .ZN(_0882_));
 BUF_X4 _1368_ (.A(_0882_),
    .Z(_0883_));
 MUX2_X1 _1369_ (.A(\active_row[6][0] ),
    .B(_0846_),
    .S(_0883_),
    .Z(_0130_));
 MUX2_X1 _1370_ (.A(\active_row[6][10] ),
    .B(_0856_),
    .S(_0883_),
    .Z(_0131_));
 MUX2_X1 _1371_ (.A(\active_row[6][11] ),
    .B(_0857_),
    .S(_0883_),
    .Z(_0132_));
 MUX2_X1 _1372_ (.A(\active_row[6][12] ),
    .B(_0858_),
    .S(_0883_),
    .Z(_0133_));
 MUX2_X1 _1373_ (.A(\active_row[6][13] ),
    .B(_0859_),
    .S(_0883_),
    .Z(_0134_));
 MUX2_X1 _1374_ (.A(\active_row[6][1] ),
    .B(_0860_),
    .S(_0883_),
    .Z(_0135_));
 MUX2_X1 _1375_ (.A(\active_row[6][2] ),
    .B(_0861_),
    .S(_0883_),
    .Z(_0136_));
 MUX2_X1 _1376_ (.A(\active_row[6][3] ),
    .B(_0862_),
    .S(_0883_),
    .Z(_0137_));
 MUX2_X1 _1377_ (.A(\active_row[6][4] ),
    .B(_0863_),
    .S(_0883_),
    .Z(_0138_));
 MUX2_X1 _1378_ (.A(\active_row[6][5] ),
    .B(_0864_),
    .S(_0883_),
    .Z(_0139_));
 MUX2_X1 _1379_ (.A(\active_row[6][6] ),
    .B(_0865_),
    .S(_0882_),
    .Z(_0140_));
 MUX2_X1 _1380_ (.A(\active_row[6][7] ),
    .B(_0866_),
    .S(_0882_),
    .Z(_0141_));
 MUX2_X1 _1381_ (.A(\active_row[6][8] ),
    .B(_0867_),
    .S(_0882_),
    .Z(_0142_));
 MUX2_X1 _1382_ (.A(\active_row[6][9] ),
    .B(_0868_),
    .S(_0882_),
    .Z(_0143_));
 NOR3_X4 _1383_ (.A1(_0848_),
    .A2(_1145_),
    .A3(_0873_),
    .ZN(_0884_));
 BUF_X4 _1384_ (.A(_0884_),
    .Z(_0885_));
 MUX2_X1 _1385_ (.A(\active_row[7][0] ),
    .B(_0846_),
    .S(_0885_),
    .Z(_0144_));
 MUX2_X1 _1386_ (.A(\active_row[7][10] ),
    .B(_0856_),
    .S(_0885_),
    .Z(_0145_));
 MUX2_X1 _1387_ (.A(\active_row[7][11] ),
    .B(_0857_),
    .S(_0885_),
    .Z(_0146_));
 MUX2_X1 _1388_ (.A(\active_row[7][12] ),
    .B(_0858_),
    .S(_0885_),
    .Z(_0147_));
 MUX2_X1 _1389_ (.A(\active_row[7][13] ),
    .B(_0859_),
    .S(_0885_),
    .Z(_0148_));
 MUX2_X1 _1390_ (.A(\active_row[7][1] ),
    .B(_0860_),
    .S(_0885_),
    .Z(_0149_));
 MUX2_X1 _1391_ (.A(\active_row[7][2] ),
    .B(_0861_),
    .S(_0885_),
    .Z(_0150_));
 MUX2_X1 _1392_ (.A(\active_row[7][3] ),
    .B(_0862_),
    .S(_0885_),
    .Z(_0151_));
 MUX2_X1 _1393_ (.A(\active_row[7][4] ),
    .B(_0863_),
    .S(_0885_),
    .Z(_0152_));
 MUX2_X1 _1394_ (.A(\active_row[7][5] ),
    .B(_0864_),
    .S(_0885_),
    .Z(_0153_));
 MUX2_X1 _1395_ (.A(\active_row[7][6] ),
    .B(_0865_),
    .S(_0884_),
    .Z(_0154_));
 MUX2_X1 _1396_ (.A(\active_row[7][7] ),
    .B(_0866_),
    .S(_0884_),
    .Z(_0155_));
 MUX2_X1 _1397_ (.A(\active_row[7][8] ),
    .B(_0867_),
    .S(_0884_),
    .Z(_0156_));
 MUX2_X1 _1398_ (.A(\active_row[7][9] ),
    .B(_0868_),
    .S(_0884_),
    .Z(_0157_));
 BUF_X4 _1399_ (.A(_1188_),
    .Z(_0886_));
 INV_X2 _1400_ (.A(_0886_),
    .ZN(_0887_));
 CLKBUF_X3 _1401_ (.A(_0887_),
    .Z(_0888_));
 INV_X1 _1402_ (.A(net118),
    .ZN(_0889_));
 CLKBUF_X2 _1403_ (.A(net130),
    .Z(_0890_));
 NAND3_X2 _1404_ (.A1(_0889_),
    .A2(_0890_),
    .A3(net128),
    .ZN(_0891_));
 OR2_X1 _1405_ (.A1(_0888_),
    .A2(_0891_),
    .ZN(_0892_));
 CLKBUF_X3 _1406_ (.A(_0892_),
    .Z(_0893_));
 CLKBUF_X3 _1407_ (.A(_0893_),
    .Z(_0894_));
 MUX2_X1 _1408_ (.A(net34),
    .B(net131),
    .S(_0894_),
    .Z(_0193_));
 MUX2_X1 _1409_ (.A(net35),
    .B(net132),
    .S(_0894_),
    .Z(_0194_));
 MUX2_X1 _1410_ (.A(net36),
    .B(net133),
    .S(_0894_),
    .Z(_0195_));
 MUX2_X1 _1411_ (.A(net37),
    .B(net134),
    .S(_0894_),
    .Z(_0196_));
 MUX2_X1 _1412_ (.A(net38),
    .B(net135),
    .S(_0894_),
    .Z(_0197_));
 MUX2_X1 _1413_ (.A(net39),
    .B(net136),
    .S(_0894_),
    .Z(_0198_));
 MUX2_X1 _1414_ (.A(net40),
    .B(net137),
    .S(_0894_),
    .Z(_0199_));
 MUX2_X1 _1415_ (.A(net41),
    .B(net138),
    .S(_0894_),
    .Z(_0200_));
 MUX2_X1 _1416_ (.A(net42),
    .B(net139),
    .S(_0894_),
    .Z(_0201_));
 MUX2_X1 _1417_ (.A(net43),
    .B(net140),
    .S(_0894_),
    .Z(_0202_));
 CLKBUF_X3 _1418_ (.A(_0893_),
    .Z(_0895_));
 MUX2_X1 _1419_ (.A(net44),
    .B(net141),
    .S(_0895_),
    .Z(_0203_));
 MUX2_X1 _1420_ (.A(net45),
    .B(net142),
    .S(_0895_),
    .Z(_0204_));
 MUX2_X1 _1421_ (.A(net46),
    .B(net143),
    .S(_0895_),
    .Z(_0205_));
 MUX2_X1 _1422_ (.A(net47),
    .B(net144),
    .S(_0895_),
    .Z(_0206_));
 MUX2_X1 _1423_ (.A(net48),
    .B(net145),
    .S(_0895_),
    .Z(_0207_));
 MUX2_X1 _1424_ (.A(net49),
    .B(net146),
    .S(_0895_),
    .Z(_0208_));
 MUX2_X1 _1425_ (.A(net50),
    .B(net147),
    .S(_0895_),
    .Z(_0209_));
 MUX2_X1 _1426_ (.A(net51),
    .B(net148),
    .S(_0895_),
    .Z(_0210_));
 MUX2_X1 _1427_ (.A(net52),
    .B(net149),
    .S(_0895_),
    .Z(_0211_));
 MUX2_X1 _1428_ (.A(net53),
    .B(net150),
    .S(_0895_),
    .Z(_0212_));
 CLKBUF_X3 _1429_ (.A(_0893_),
    .Z(_0896_));
 MUX2_X1 _1430_ (.A(net54),
    .B(net151),
    .S(_0896_),
    .Z(_0213_));
 MUX2_X1 _1431_ (.A(net55),
    .B(net152),
    .S(_0896_),
    .Z(_0214_));
 MUX2_X1 _1432_ (.A(net56),
    .B(net153),
    .S(_0896_),
    .Z(_0215_));
 MUX2_X1 _1433_ (.A(net57),
    .B(net154),
    .S(_0896_),
    .Z(_0216_));
 MUX2_X1 _1434_ (.A(net58),
    .B(net155),
    .S(_0896_),
    .Z(_0217_));
 MUX2_X1 _1435_ (.A(net59),
    .B(net156),
    .S(_0896_),
    .Z(_0218_));
 MUX2_X1 _1436_ (.A(net60),
    .B(net157),
    .S(_0896_),
    .Z(_0219_));
 MUX2_X1 _1437_ (.A(net61),
    .B(net158),
    .S(_0896_),
    .Z(_0220_));
 MUX2_X1 _1438_ (.A(net62),
    .B(net159),
    .S(_0896_),
    .Z(_0221_));
 MUX2_X1 _1439_ (.A(net63),
    .B(net160),
    .S(_0896_),
    .Z(_0222_));
 CLKBUF_X3 _1440_ (.A(_0893_),
    .Z(_0897_));
 MUX2_X1 _1441_ (.A(net64),
    .B(net161),
    .S(_0897_),
    .Z(_0223_));
 MUX2_X1 _1442_ (.A(net65),
    .B(net162),
    .S(_0897_),
    .Z(_0224_));
 MUX2_X1 _1443_ (.A(net66),
    .B(net163),
    .S(_0897_),
    .Z(_0225_));
 MUX2_X1 _1444_ (.A(net67),
    .B(net164),
    .S(_0897_),
    .Z(_0226_));
 MUX2_X1 _1445_ (.A(net68),
    .B(net165),
    .S(_0897_),
    .Z(_0227_));
 MUX2_X1 _1446_ (.A(net69),
    .B(net166),
    .S(_0897_),
    .Z(_0228_));
 MUX2_X1 _1447_ (.A(net70),
    .B(net167),
    .S(_0897_),
    .Z(_0229_));
 MUX2_X1 _1448_ (.A(net71),
    .B(net168),
    .S(_0897_),
    .Z(_0230_));
 MUX2_X1 _1449_ (.A(net72),
    .B(net169),
    .S(_0897_),
    .Z(_0231_));
 MUX2_X1 _1450_ (.A(net73),
    .B(net170),
    .S(_0897_),
    .Z(_0232_));
 CLKBUF_X3 _1451_ (.A(_0893_),
    .Z(_0898_));
 MUX2_X1 _1452_ (.A(net74),
    .B(net171),
    .S(_0898_),
    .Z(_0233_));
 MUX2_X1 _1453_ (.A(net75),
    .B(net172),
    .S(_0898_),
    .Z(_0234_));
 MUX2_X1 _1454_ (.A(net76),
    .B(net173),
    .S(_0898_),
    .Z(_0235_));
 MUX2_X1 _1455_ (.A(net77),
    .B(net174),
    .S(_0898_),
    .Z(_0236_));
 MUX2_X1 _1456_ (.A(net78),
    .B(net175),
    .S(_0898_),
    .Z(_0237_));
 MUX2_X1 _1457_ (.A(net79),
    .B(net176),
    .S(_0898_),
    .Z(_0238_));
 MUX2_X1 _1458_ (.A(net80),
    .B(net177),
    .S(_0898_),
    .Z(_0239_));
 MUX2_X1 _1459_ (.A(net81),
    .B(net178),
    .S(_0898_),
    .Z(_0240_));
 MUX2_X1 _1460_ (.A(net82),
    .B(net179),
    .S(_0898_),
    .Z(_0241_));
 MUX2_X1 _1461_ (.A(net83),
    .B(net180),
    .S(_0898_),
    .Z(_0242_));
 CLKBUF_X3 _1462_ (.A(_0893_),
    .Z(_0899_));
 MUX2_X1 _1463_ (.A(net84),
    .B(net181),
    .S(_0899_),
    .Z(_0243_));
 MUX2_X1 _1464_ (.A(net85),
    .B(net182),
    .S(_0899_),
    .Z(_0244_));
 MUX2_X1 _1465_ (.A(net86),
    .B(net183),
    .S(_0899_),
    .Z(_0245_));
 MUX2_X1 _1466_ (.A(net87),
    .B(net184),
    .S(_0899_),
    .Z(_0246_));
 MUX2_X1 _1467_ (.A(net88),
    .B(net185),
    .S(_0899_),
    .Z(_0247_));
 MUX2_X1 _1468_ (.A(net89),
    .B(net186),
    .S(_0899_),
    .Z(_0248_));
 MUX2_X1 _1469_ (.A(net90),
    .B(net187),
    .S(_0899_),
    .Z(_0249_));
 MUX2_X1 _1470_ (.A(net91),
    .B(net188),
    .S(_0899_),
    .Z(_0250_));
 MUX2_X1 _1471_ (.A(net92),
    .B(net189),
    .S(_0899_),
    .Z(_0251_));
 MUX2_X1 _1472_ (.A(net93),
    .B(net190),
    .S(_0899_),
    .Z(_0252_));
 MUX2_X1 _1473_ (.A(net94),
    .B(net191),
    .S(_0893_),
    .Z(_0253_));
 MUX2_X1 _1474_ (.A(net95),
    .B(net192),
    .S(_0893_),
    .Z(_0254_));
 MUX2_X1 _1475_ (.A(net96),
    .B(net193),
    .S(_0893_),
    .Z(_0255_));
 MUX2_X1 _1476_ (.A(net97),
    .B(net194),
    .S(_0893_),
    .Z(_0256_));
 OR3_X1 _1477_ (.A1(_0824_),
    .A2(_0828_),
    .A3(\init_state[6] ),
    .ZN(_0900_));
 AOI21_X2 _1478_ (.A(_0805_),
    .B1(_0817_),
    .B2(_0900_),
    .ZN(_0901_));
 BUF_X4 _1479_ (.A(_1186_),
    .Z(_0902_));
 INV_X2 _1480_ (.A(_0902_),
    .ZN(_0903_));
 CLKBUF_X2 _1481_ (.A(cmd_valid),
    .Z(_0904_));
 INV_X1 _1482_ (.A(_0904_),
    .ZN(_0905_));
 NOR3_X4 _1483_ (.A1(_0905_),
    .A2(_0810_),
    .A3(_0816_),
    .ZN(_0906_));
 AOI21_X4 _1484_ (.A(_0903_),
    .B1(_1162_),
    .B2(_0906_),
    .ZN(_0907_));
 NOR2_X4 _1485_ (.A1(_0901_),
    .A2(_0907_),
    .ZN(_0908_));
 NOR4_X4 _1486_ (.A1(_0804_),
    .A2(_0902_),
    .A3(_0886_),
    .A4(_0850_),
    .ZN(_0909_));
 NOR2_X4 _1487_ (.A1(_0851_),
    .A2(_0817_),
    .ZN(_0910_));
 INV_X1 _1488_ (.A(\burst_counter[3] ),
    .ZN(_0911_));
 INV_X1 _1489_ (.A(\burst_counter[2] ),
    .ZN(_0912_));
 NAND3_X4 _1490_ (.A1(_0911_),
    .A2(_0912_),
    .A3(_1157_),
    .ZN(_0913_));
 INV_X2 _1491_ (.A(_0913_),
    .ZN(_0914_));
 AOI21_X4 _1492_ (.A(_0887_),
    .B1(_0817_),
    .B2(_0914_),
    .ZN(_0915_));
 NOR3_X4 _1493_ (.A1(_0909_),
    .A2(_0910_),
    .A3(_0915_),
    .ZN(_0916_));
 AOI21_X4 _1494_ (.A(_0833_),
    .B1(_0908_),
    .B2(_0916_),
    .ZN(_0917_));
 NAND2_X1 _1495_ (.A1(_0846_),
    .A2(_0917_),
    .ZN(_0918_));
 NAND2_X2 _1496_ (.A1(_0908_),
    .A2(_0916_),
    .ZN(_0919_));
 CLKBUF_X3 _1497_ (.A(_0919_),
    .Z(_0920_));
 NOR2_X1 _1498_ (.A1(_0833_),
    .A2(_0920_),
    .ZN(_0921_));
 BUF_X4 _1499_ (.A(_0804_),
    .Z(_0922_));
 CLKBUF_X3 _1500_ (.A(_0922_),
    .Z(_0923_));
 OAI21_X1 _1501_ (.A(_0923_),
    .B1(_0824_),
    .B2(_0828_),
    .ZN(_0924_));
 NAND2_X1 _1502_ (.A1(_0921_),
    .A2(_0924_),
    .ZN(_0925_));
 NAND2_X1 _1503_ (.A1(_0806_),
    .A2(_0888_),
    .ZN(_0926_));
 BUF_X4 _1504_ (.A(cmd_addr[12]),
    .Z(_0927_));
 BUF_X8 _1505_ (.A(_0927_),
    .Z(_0928_));
 BUF_X4 _1506_ (.A(_0928_),
    .Z(_0929_));
 BUF_X4 _1507_ (.A(_0929_),
    .Z(_0930_));
 MUX2_X1 _1508_ (.A(_0028_),
    .B(_0030_),
    .S(_0930_),
    .Z(_0931_));
 MUX2_X1 _1509_ (.A(_0029_),
    .B(_0031_),
    .S(_0930_),
    .Z(_0932_));
 BUF_X4 _1510_ (.A(cmd_addr[11]),
    .Z(_0933_));
 BUF_X4 _1511_ (.A(_0933_),
    .Z(_0934_));
 MUX2_X1 _1512_ (.A(_0931_),
    .B(_0932_),
    .S(_0934_),
    .Z(_0935_));
 MUX2_X1 _1513_ (.A(_0024_),
    .B(_0026_),
    .S(_0930_),
    .Z(_0936_));
 MUX2_X1 _1514_ (.A(_0025_),
    .B(_0027_),
    .S(_0930_),
    .Z(_0937_));
 MUX2_X1 _1515_ (.A(_0936_),
    .B(_0937_),
    .S(_0934_),
    .Z(_0938_));
 BUF_X4 _1516_ (.A(net2),
    .Z(_0291_));
 INV_X2 _1517_ (.A(_0291_),
    .ZN(_0292_));
 BUF_X4 _1518_ (.A(_0292_),
    .Z(_0293_));
 MUX2_X1 _1519_ (.A(_0935_),
    .B(_0938_),
    .S(_0293_),
    .Z(_0294_));
 CLKBUF_X3 _1520_ (.A(_0291_),
    .Z(_0295_));
 INV_X1 _1521_ (.A(_0933_),
    .ZN(_0296_));
 CLKBUF_X3 _1522_ (.A(_0296_),
    .Z(_0297_));
 MUX2_X1 _1523_ (.A(\active_row[1][11] ),
    .B(\active_row[3][11] ),
    .S(_0929_),
    .Z(_0298_));
 NOR3_X1 _1524_ (.A1(_0295_),
    .A2(_0297_),
    .A3(_0298_),
    .ZN(_0299_));
 OR2_X1 _1525_ (.A1(net2),
    .A2(_0933_),
    .ZN(_0300_));
 CLKBUF_X3 _1526_ (.A(_0300_),
    .Z(_0301_));
 MUX2_X1 _1527_ (.A(\active_row[0][11] ),
    .B(\active_row[2][11] ),
    .S(_0929_),
    .Z(_0302_));
 NOR2_X1 _1528_ (.A1(_0301_),
    .A2(_0302_),
    .ZN(_0303_));
 NAND2_X4 _1529_ (.A1(_0291_),
    .A2(_0933_),
    .ZN(_0304_));
 MUX2_X1 _1530_ (.A(\active_row[5][11] ),
    .B(\active_row[7][11] ),
    .S(_0929_),
    .Z(_0305_));
 NOR2_X1 _1531_ (.A1(_0304_),
    .A2(_0305_),
    .ZN(_0306_));
 BUF_X4 _1532_ (.A(_0927_),
    .Z(_0307_));
 MUX2_X1 _1533_ (.A(\active_row[4][11] ),
    .B(\active_row[6][11] ),
    .S(_0307_),
    .Z(_0308_));
 NOR3_X1 _1534_ (.A1(_0292_),
    .A2(_0934_),
    .A3(_0308_),
    .ZN(_0309_));
 NOR4_X2 _1535_ (.A1(_0299_),
    .A2(_0303_),
    .A3(_0306_),
    .A4(_0309_),
    .ZN(_0310_));
 XOR2_X2 _1536_ (.A(net15),
    .B(_0310_),
    .Z(_0311_));
 CLKBUF_X3 _1537_ (.A(_0933_),
    .Z(_0312_));
 MUX2_X1 _1538_ (.A(\active_row[6][5] ),
    .B(\active_row[7][5] ),
    .S(_0312_),
    .Z(_0313_));
 NAND3_X1 _1539_ (.A1(_0295_),
    .A2(_0930_),
    .A3(_0313_),
    .ZN(_0314_));
 INV_X1 _1540_ (.A(_0930_),
    .ZN(_0315_));
 MUX2_X1 _1541_ (.A(\active_row[4][5] ),
    .B(\active_row[5][5] ),
    .S(_0933_),
    .Z(_0316_));
 NAND3_X1 _1542_ (.A1(_0295_),
    .A2(_0315_),
    .A3(_0316_),
    .ZN(_0317_));
 BUF_X4 _1543_ (.A(_0928_),
    .Z(_0318_));
 MUX2_X1 _1544_ (.A(\active_row[1][5] ),
    .B(\active_row[3][5] ),
    .S(_0318_),
    .Z(_0319_));
 NAND3_X1 _1545_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0319_),
    .ZN(_0320_));
 NOR2_X1 _1546_ (.A1(_0291_),
    .A2(_0312_),
    .ZN(_0321_));
 MUX2_X1 _1547_ (.A(\active_row[0][5] ),
    .B(\active_row[2][5] ),
    .S(_0318_),
    .Z(_0322_));
 NAND2_X1 _1548_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0323_));
 NAND4_X2 _1549_ (.A1(_0314_),
    .A2(_0317_),
    .A3(_0320_),
    .A4(_0323_),
    .ZN(_0324_));
 XOR2_X2 _1550_ (.A(net8),
    .B(_0324_),
    .Z(_0325_));
 MUX2_X1 _1551_ (.A(\active_row[1][0] ),
    .B(\active_row[3][0] ),
    .S(_0307_),
    .Z(_0326_));
 NOR3_X1 _1552_ (.A1(_0295_),
    .A2(_0297_),
    .A3(_0326_),
    .ZN(_0327_));
 MUX2_X1 _1553_ (.A(\active_row[0][0] ),
    .B(\active_row[2][0] ),
    .S(_0929_),
    .Z(_0328_));
 NOR2_X1 _1554_ (.A1(_0301_),
    .A2(_0328_),
    .ZN(_0329_));
 MUX2_X1 _1555_ (.A(\active_row[5][0] ),
    .B(\active_row[7][0] ),
    .S(_0307_),
    .Z(_0330_));
 NOR2_X1 _1556_ (.A1(_0304_),
    .A2(_0330_),
    .ZN(_0331_));
 BUF_X4 _1557_ (.A(_0927_),
    .Z(_0332_));
 MUX2_X1 _1558_ (.A(\active_row[4][0] ),
    .B(\active_row[6][0] ),
    .S(_0332_),
    .Z(_0333_));
 NOR3_X1 _1559_ (.A1(_0292_),
    .A2(_0312_),
    .A3(_0333_),
    .ZN(_0334_));
 NOR4_X2 _1560_ (.A1(_0327_),
    .A2(_0329_),
    .A3(_0331_),
    .A4(_0334_),
    .ZN(_0335_));
 XOR2_X2 _1561_ (.A(net3),
    .B(_0335_),
    .Z(_0336_));
 NOR4_X2 _1562_ (.A1(_0294_),
    .A2(_0311_),
    .A3(_0325_),
    .A4(_0336_),
    .ZN(_0337_));
 MUX2_X1 _1563_ (.A(\active_row[4][13] ),
    .B(\active_row[5][13] ),
    .S(_0312_),
    .Z(_0338_));
 NAND3_X1 _1564_ (.A1(_0295_),
    .A2(_0315_),
    .A3(_0338_),
    .ZN(_0339_));
 MUX2_X1 _1565_ (.A(\active_row[6][13] ),
    .B(\active_row[7][13] ),
    .S(_0312_),
    .Z(_0340_));
 NAND3_X1 _1566_ (.A1(_0295_),
    .A2(_0930_),
    .A3(_0340_),
    .ZN(_0341_));
 MUX2_X1 _1567_ (.A(\active_row[1][13] ),
    .B(\active_row[3][13] ),
    .S(_0318_),
    .Z(_0342_));
 NAND3_X1 _1568_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0342_),
    .ZN(_0343_));
 MUX2_X1 _1569_ (.A(\active_row[0][13] ),
    .B(\active_row[2][13] ),
    .S(_0930_),
    .Z(_0344_));
 NAND2_X1 _1570_ (.A1(_0321_),
    .A2(_0344_),
    .ZN(_0345_));
 NAND4_X2 _1571_ (.A1(_0339_),
    .A2(_0341_),
    .A3(_0343_),
    .A4(_0345_),
    .ZN(_0346_));
 XOR2_X2 _1572_ (.A(net17),
    .B(_0346_),
    .Z(_0347_));
 MUX2_X1 _1573_ (.A(\active_row[6][12] ),
    .B(\active_row[7][12] ),
    .S(_0312_),
    .Z(_0348_));
 NAND3_X1 _1574_ (.A1(_0295_),
    .A2(_0930_),
    .A3(_0348_),
    .ZN(_0349_));
 MUX2_X1 _1575_ (.A(\active_row[4][12] ),
    .B(\active_row[5][12] ),
    .S(_0312_),
    .Z(_0350_));
 NAND3_X1 _1576_ (.A1(_0295_),
    .A2(_0315_),
    .A3(_0350_),
    .ZN(_0351_));
 MUX2_X1 _1577_ (.A(\active_row[1][12] ),
    .B(\active_row[3][12] ),
    .S(_0318_),
    .Z(_0352_));
 NAND3_X1 _1578_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0352_),
    .ZN(_0353_));
 MUX2_X1 _1579_ (.A(\active_row[0][12] ),
    .B(\active_row[2][12] ),
    .S(_0318_),
    .Z(_0354_));
 NAND2_X1 _1580_ (.A1(_0321_),
    .A2(_0354_),
    .ZN(_0355_));
 NAND4_X2 _1581_ (.A1(_0349_),
    .A2(_0351_),
    .A3(_0353_),
    .A4(_0355_),
    .ZN(_0356_));
 XOR2_X2 _1582_ (.A(net16),
    .B(_0356_),
    .Z(_0357_));
 MUX2_X1 _1583_ (.A(\active_row[1][6] ),
    .B(\active_row[3][6] ),
    .S(_0318_),
    .Z(_0358_));
 NOR3_X1 _1584_ (.A1(_0295_),
    .A2(_0297_),
    .A3(_0358_),
    .ZN(_0359_));
 MUX2_X1 _1585_ (.A(\active_row[0][6] ),
    .B(\active_row[2][6] ),
    .S(_0318_),
    .Z(_0360_));
 NOR2_X1 _1586_ (.A1(_0301_),
    .A2(_0360_),
    .ZN(_0361_));
 MUX2_X1 _1587_ (.A(\active_row[5][6] ),
    .B(\active_row[7][6] ),
    .S(_0929_),
    .Z(_0362_));
 NOR2_X1 _1588_ (.A1(_0304_),
    .A2(_0362_),
    .ZN(_0363_));
 MUX2_X1 _1589_ (.A(\active_row[4][6] ),
    .B(\active_row[6][6] ),
    .S(_0307_),
    .Z(_0364_));
 NOR3_X1 _1590_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0364_),
    .ZN(_0365_));
 NOR4_X2 _1591_ (.A1(_0359_),
    .A2(_0361_),
    .A3(_0363_),
    .A4(_0365_),
    .ZN(_0366_));
 XOR2_X2 _1592_ (.A(net10),
    .B(_0366_),
    .Z(_0367_));
 NOR3_X2 _1593_ (.A1(_0347_),
    .A2(_0357_),
    .A3(_0367_),
    .ZN(_0368_));
 MUX2_X1 _1594_ (.A(\active_row[5][2] ),
    .B(\active_row[7][2] ),
    .S(_0928_),
    .Z(_0369_));
 MUX2_X1 _1595_ (.A(\active_row[4][2] ),
    .B(\active_row[6][2] ),
    .S(_0928_),
    .Z(_0370_));
 MUX2_X1 _1596_ (.A(_0369_),
    .B(_0370_),
    .S(_0296_),
    .Z(_0371_));
 MUX2_X1 _1597_ (.A(\active_row[1][2] ),
    .B(\active_row[3][2] ),
    .S(_0332_),
    .Z(_0372_));
 MUX2_X1 _1598_ (.A(\active_row[0][2] ),
    .B(\active_row[2][2] ),
    .S(_0332_),
    .Z(_0373_));
 MUX2_X1 _1599_ (.A(_0372_),
    .B(_0373_),
    .S(_0297_),
    .Z(_0374_));
 MUX2_X1 _1600_ (.A(_0371_),
    .B(_0374_),
    .S(_0293_),
    .Z(_0375_));
 XOR2_X2 _1601_ (.A(net5),
    .B(_0375_),
    .Z(_0376_));
 MUX2_X1 _1602_ (.A(\active_row[0][10] ),
    .B(\active_row[2][10] ),
    .S(_0929_),
    .Z(_0377_));
 NOR2_X1 _1603_ (.A1(_0301_),
    .A2(_0377_),
    .ZN(_0378_));
 MUX2_X1 _1604_ (.A(\active_row[1][10] ),
    .B(\active_row[3][10] ),
    .S(_0332_),
    .Z(_0379_));
 NOR3_X1 _1605_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0379_),
    .ZN(_0380_));
 MUX2_X1 _1606_ (.A(\active_row[4][10] ),
    .B(\active_row[6][10] ),
    .S(_0332_),
    .Z(_0381_));
 NOR3_X1 _1607_ (.A1(_0292_),
    .A2(_0312_),
    .A3(_0381_),
    .ZN(_0382_));
 MUX2_X1 _1608_ (.A(\active_row[5][10] ),
    .B(\active_row[7][10] ),
    .S(_0307_),
    .Z(_0383_));
 NOR2_X1 _1609_ (.A1(_0304_),
    .A2(_0383_),
    .ZN(_0384_));
 NOR4_X2 _1610_ (.A1(_0378_),
    .A2(_0380_),
    .A3(_0382_),
    .A4(_0384_),
    .ZN(_0385_));
 XOR2_X2 _1611_ (.A(net14),
    .B(_0385_),
    .Z(_0386_));
 MUX2_X1 _1612_ (.A(\active_row[0][7] ),
    .B(\active_row[2][7] ),
    .S(_0929_),
    .Z(_0387_));
 NOR2_X1 _1613_ (.A1(_0301_),
    .A2(_0387_),
    .ZN(_0388_));
 MUX2_X1 _1614_ (.A(\active_row[1][7] ),
    .B(\active_row[3][7] ),
    .S(_0332_),
    .Z(_0389_));
 NOR3_X1 _1615_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0389_),
    .ZN(_0390_));
 MUX2_X1 _1616_ (.A(\active_row[4][7] ),
    .B(\active_row[6][7] ),
    .S(_0928_),
    .Z(_0391_));
 NOR3_X1 _1617_ (.A1(_0292_),
    .A2(_0312_),
    .A3(_0391_),
    .ZN(_0392_));
 MUX2_X1 _1618_ (.A(\active_row[5][7] ),
    .B(\active_row[7][7] ),
    .S(_0332_),
    .Z(_0393_));
 NOR2_X1 _1619_ (.A1(_0304_),
    .A2(_0393_),
    .ZN(_0394_));
 NOR4_X2 _1620_ (.A1(_0388_),
    .A2(_0390_),
    .A3(_0392_),
    .A4(_0394_),
    .ZN(_0395_));
 XOR2_X2 _1621_ (.A(net11),
    .B(_0395_),
    .Z(_0396_));
 MUX2_X1 _1622_ (.A(\active_row[0][1] ),
    .B(\active_row[2][1] ),
    .S(_0929_),
    .Z(_0397_));
 NOR2_X1 _1623_ (.A1(_0301_),
    .A2(_0397_),
    .ZN(_0398_));
 MUX2_X1 _1624_ (.A(\active_row[1][1] ),
    .B(\active_row[3][1] ),
    .S(_0332_),
    .Z(_0399_));
 NOR3_X1 _1625_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0399_),
    .ZN(_0400_));
 MUX2_X1 _1626_ (.A(\active_row[4][1] ),
    .B(\active_row[6][1] ),
    .S(_0928_),
    .Z(_0401_));
 NOR3_X1 _1627_ (.A1(_0292_),
    .A2(_0312_),
    .A3(_0401_),
    .ZN(_0402_));
 MUX2_X1 _1628_ (.A(\active_row[5][1] ),
    .B(\active_row[7][1] ),
    .S(_0332_),
    .Z(_0403_));
 NOR2_X1 _1629_ (.A1(_0304_),
    .A2(_0403_),
    .ZN(_0404_));
 NOR4_X2 _1630_ (.A1(_0398_),
    .A2(_0400_),
    .A3(_0402_),
    .A4(_0404_),
    .ZN(_0405_));
 XOR2_X2 _1631_ (.A(net4),
    .B(_0405_),
    .Z(_0406_));
 NOR4_X4 _1632_ (.A1(_0376_),
    .A2(_0386_),
    .A3(_0396_),
    .A4(_0406_),
    .ZN(_0407_));
 MUX2_X1 _1633_ (.A(\active_row[0][9] ),
    .B(\active_row[2][9] ),
    .S(_0318_),
    .Z(_0408_));
 NOR2_X1 _1634_ (.A1(_0301_),
    .A2(_0408_),
    .ZN(_0409_));
 MUX2_X1 _1635_ (.A(\active_row[1][9] ),
    .B(\active_row[3][9] ),
    .S(_0307_),
    .Z(_0410_));
 NOR3_X1 _1636_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0410_),
    .ZN(_0411_));
 MUX2_X1 _1637_ (.A(\active_row[4][9] ),
    .B(\active_row[6][9] ),
    .S(_0307_),
    .Z(_0412_));
 NOR3_X1 _1638_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0412_),
    .ZN(_0413_));
 MUX2_X1 _1639_ (.A(\active_row[5][9] ),
    .B(\active_row[7][9] ),
    .S(_0929_),
    .Z(_0414_));
 NOR2_X1 _1640_ (.A1(_0304_),
    .A2(_0414_),
    .ZN(_0415_));
 NOR4_X2 _1641_ (.A1(_0409_),
    .A2(_0411_),
    .A3(_0413_),
    .A4(_0415_),
    .ZN(_0416_));
 XOR2_X2 _1642_ (.A(net13),
    .B(_0416_),
    .Z(_0417_));
 MUX2_X1 _1643_ (.A(\active_row[4][4] ),
    .B(\active_row[6][4] ),
    .S(_0307_),
    .Z(_0418_));
 NOR3_X1 _1644_ (.A1(_0293_),
    .A2(_0934_),
    .A3(_0418_),
    .ZN(_0419_));
 MUX2_X1 _1645_ (.A(\active_row[5][4] ),
    .B(\active_row[7][4] ),
    .S(_0307_),
    .Z(_0420_));
 NOR2_X1 _1646_ (.A1(_0304_),
    .A2(_0420_),
    .ZN(_0421_));
 MUX2_X1 _1647_ (.A(\active_row[0][4] ),
    .B(\active_row[2][4] ),
    .S(_0307_),
    .Z(_0422_));
 NOR2_X1 _1648_ (.A1(_0301_),
    .A2(_0422_),
    .ZN(_0423_));
 MUX2_X1 _1649_ (.A(\active_row[1][4] ),
    .B(\active_row[3][4] ),
    .S(_0928_),
    .Z(_0424_));
 NOR3_X1 _1650_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0424_),
    .ZN(_0425_));
 NOR4_X2 _1651_ (.A1(_0419_),
    .A2(_0421_),
    .A3(_0423_),
    .A4(_0425_),
    .ZN(_0426_));
 XOR2_X2 _1652_ (.A(net7),
    .B(_0426_),
    .Z(_0427_));
 MUX2_X1 _1653_ (.A(\active_row[4][8] ),
    .B(\active_row[6][8] ),
    .S(_0927_),
    .Z(_0428_));
 MUX2_X1 _1654_ (.A(\active_row[5][8] ),
    .B(\active_row[7][8] ),
    .S(_0928_),
    .Z(_0429_));
 MUX2_X1 _1655_ (.A(_0428_),
    .B(_0429_),
    .S(_0933_),
    .Z(_0430_));
 MUX2_X1 _1656_ (.A(\active_row[0][8] ),
    .B(\active_row[2][8] ),
    .S(_0928_),
    .Z(_0431_));
 MUX2_X1 _1657_ (.A(\active_row[1][8] ),
    .B(\active_row[3][8] ),
    .S(_0928_),
    .Z(_0432_));
 MUX2_X1 _1658_ (.A(_0431_),
    .B(_0432_),
    .S(_0933_),
    .Z(_0433_));
 MUX2_X1 _1659_ (.A(_0430_),
    .B(_0433_),
    .S(_0293_),
    .Z(_0434_));
 XOR2_X2 _1660_ (.A(net12),
    .B(_0434_),
    .Z(_0435_));
 MUX2_X1 _1661_ (.A(\active_row[1][3] ),
    .B(\active_row[3][3] ),
    .S(_0332_),
    .Z(_0436_));
 OR3_X1 _1662_ (.A1(_0291_),
    .A2(_0297_),
    .A3(_0436_),
    .ZN(_0437_));
 MUX2_X1 _1663_ (.A(\active_row[0][3] ),
    .B(\active_row[2][3] ),
    .S(_0318_),
    .Z(_0438_));
 MUX2_X1 _1664_ (.A(\active_row[4][3] ),
    .B(\active_row[5][3] ),
    .S(_0933_),
    .Z(_0439_));
 MUX2_X1 _1665_ (.A(\active_row[6][3] ),
    .B(\active_row[7][3] ),
    .S(_0933_),
    .Z(_0440_));
 MUX2_X1 _1666_ (.A(_0439_),
    .B(_0440_),
    .S(_0318_),
    .Z(_0441_));
 OAI221_X2 _1667_ (.A(_0437_),
    .B1(_0438_),
    .B2(_0301_),
    .C1(_0441_),
    .C2(_0293_),
    .ZN(_0442_));
 XNOR2_X2 _1668_ (.A(net6),
    .B(_0442_),
    .ZN(_0443_));
 NOR4_X4 _1669_ (.A1(_0417_),
    .A2(_0427_),
    .A3(_0435_),
    .A4(_0443_),
    .ZN(_0444_));
 NAND4_X4 _1670_ (.A1(_0337_),
    .A2(_0368_),
    .A3(_0407_),
    .A4(_0444_),
    .ZN(_0445_));
 MUX2_X1 _1671_ (.A(net1),
    .B(net3),
    .S(_0445_),
    .Z(_0446_));
 BUF_X4 _1672_ (.A(_0902_),
    .Z(_0447_));
 BUF_X4 _1673_ (.A(_0850_),
    .Z(_0448_));
 AOI221_X2 _1674_ (.A(_0926_),
    .B1(_0446_),
    .B2(_0447_),
    .C1(_0448_),
    .C2(net1),
    .ZN(_0449_));
 OAI21_X1 _1675_ (.A(_0918_),
    .B1(_0925_),
    .B2(_0449_),
    .ZN(_0158_));
 NAND2_X1 _1676_ (.A1(_0856_),
    .A2(_0917_),
    .ZN(_0450_));
 NAND2_X1 _1677_ (.A1(_0806_),
    .A2(_0921_),
    .ZN(_0451_));
 CLKBUF_X3 _1678_ (.A(_0886_),
    .Z(_0452_));
 BUF_X4 _1679_ (.A(_0452_),
    .Z(_0453_));
 AND2_X2 _1680_ (.A1(_0447_),
    .A2(_0445_),
    .ZN(_0454_));
 AOI21_X1 _1681_ (.A(_0453_),
    .B1(net14),
    .B2(_0454_),
    .ZN(_0455_));
 OAI21_X1 _1682_ (.A(_0450_),
    .B1(_0451_),
    .B2(_0455_),
    .ZN(_0159_));
 NOR2_X4 _1683_ (.A1(_0806_),
    .A2(_0824_),
    .ZN(_0456_));
 NAND2_X1 _1684_ (.A1(_0828_),
    .A2(_0456_),
    .ZN(_0457_));
 OAI21_X1 _1685_ (.A(_0801_),
    .B1(_0920_),
    .B2(_0457_),
    .ZN(_0458_));
 NAND2_X1 _1686_ (.A1(net15),
    .A2(_0454_),
    .ZN(_0459_));
 INV_X1 _1687_ (.A(_0824_),
    .ZN(_0460_));
 AOI21_X1 _1688_ (.A(_0806_),
    .B1(_0460_),
    .B2(_0828_),
    .ZN(_0461_));
 NOR3_X1 _1689_ (.A1(_0886_),
    .A2(_0919_),
    .A3(_0461_),
    .ZN(_0462_));
 INV_X1 _1690_ (.A(_0857_),
    .ZN(_0463_));
 AOI221_X1 _1691_ (.A(_0458_),
    .B1(_0459_),
    .B2(_0462_),
    .C1(_0463_),
    .C2(_0920_),
    .ZN(_0160_));
 NAND2_X1 _1692_ (.A1(_0858_),
    .A2(_0917_),
    .ZN(_0464_));
 AOI21_X1 _1693_ (.A(_0453_),
    .B1(net16),
    .B2(_0454_),
    .ZN(_0465_));
 OAI21_X1 _1694_ (.A(_0464_),
    .B1(_0465_),
    .B2(_0451_),
    .ZN(_0161_));
 NAND2_X1 _1695_ (.A1(_0859_),
    .A2(_0917_),
    .ZN(_0466_));
 AOI21_X1 _1696_ (.A(_0453_),
    .B1(net17),
    .B2(_0454_),
    .ZN(_0467_));
 OAI21_X1 _1697_ (.A(_0466_),
    .B1(_0467_),
    .B2(_0451_),
    .ZN(_0162_));
 NOR2_X2 _1698_ (.A1(_0922_),
    .A2(_0886_),
    .ZN(_0468_));
 NAND3_X2 _1699_ (.A1(_0908_),
    .A2(_0916_),
    .A3(_0468_),
    .ZN(_0469_));
 BUF_X4 _1700_ (.A(_0447_),
    .Z(_0470_));
 MUX2_X1 _1701_ (.A(net9),
    .B(net4),
    .S(_0445_),
    .Z(_0471_));
 AOI221_X2 _1702_ (.A(_0469_),
    .B1(net9),
    .B2(_0448_),
    .C1(_0470_),
    .C2(_0471_),
    .ZN(_0472_));
 NAND2_X1 _1703_ (.A1(_0860_),
    .A2(_0917_),
    .ZN(_0473_));
 AOI21_X1 _1704_ (.A(_0472_),
    .B1(_0473_),
    .B2(_0925_),
    .ZN(_0163_));
 NAND2_X1 _1705_ (.A1(_0861_),
    .A2(_0917_),
    .ZN(_0474_));
 OAI21_X1 _1706_ (.A(_0921_),
    .B1(_0828_),
    .B2(_0806_),
    .ZN(_0475_));
 MUX2_X1 _1707_ (.A(net18),
    .B(net5),
    .S(_0445_),
    .Z(_0476_));
 AOI221_X1 _1708_ (.A(_0926_),
    .B1(_0476_),
    .B2(_0447_),
    .C1(_0448_),
    .C2(net18),
    .ZN(_0477_));
 OAI21_X1 _1709_ (.A(_0474_),
    .B1(_0475_),
    .B2(_0477_),
    .ZN(_0164_));
 CLKBUF_X3 _1710_ (.A(_0802_),
    .Z(_0478_));
 AOI21_X1 _1711_ (.A(_0452_),
    .B1(_0448_),
    .B2(net19),
    .ZN(_0479_));
 NOR2_X1 _1712_ (.A1(_0923_),
    .A2(_0479_),
    .ZN(_0480_));
 MUX2_X1 _1713_ (.A(_0480_),
    .B(_0862_),
    .S(_0920_),
    .Z(_0481_));
 NAND2_X1 _1714_ (.A1(_0478_),
    .A2(_0481_),
    .ZN(_0482_));
 NOR3_X1 _1715_ (.A1(_0833_),
    .A2(_0923_),
    .A3(_0920_),
    .ZN(_0483_));
 BUF_X4 _1716_ (.A(_0445_),
    .Z(_0484_));
 MUX2_X1 _1717_ (.A(net19),
    .B(net6),
    .S(_0484_),
    .Z(_0485_));
 NAND3_X1 _1718_ (.A1(_0470_),
    .A2(_0483_),
    .A3(_0485_),
    .ZN(_0486_));
 NAND2_X1 _1719_ (.A1(_0482_),
    .A2(_0486_),
    .ZN(_0165_));
 NAND2_X1 _1720_ (.A1(_0448_),
    .A2(net20),
    .ZN(_0487_));
 AOI21_X1 _1721_ (.A(_0456_),
    .B1(_0487_),
    .B2(_0468_),
    .ZN(_0488_));
 MUX2_X1 _1722_ (.A(_0488_),
    .B(_0863_),
    .S(_0920_),
    .Z(_0489_));
 NOR4_X4 _1723_ (.A1(_0833_),
    .A2(_0903_),
    .A3(_0919_),
    .A4(_0456_),
    .ZN(_0490_));
 MUX2_X1 _1724_ (.A(net20),
    .B(net7),
    .S(_0484_),
    .Z(_0491_));
 AOI22_X1 _1725_ (.A1(_0478_),
    .A2(_0489_),
    .B1(_0490_),
    .B2(_0491_),
    .ZN(_0492_));
 INV_X1 _1726_ (.A(_0492_),
    .ZN(_0166_));
 MUX2_X1 _1727_ (.A(net21),
    .B(net8),
    .S(_0445_),
    .Z(_0493_));
 AOI221_X1 _1728_ (.A(_0469_),
    .B1(_0493_),
    .B2(_0447_),
    .C1(_0448_),
    .C2(net21),
    .ZN(_0494_));
 NAND2_X1 _1729_ (.A1(_0864_),
    .A2(_0917_),
    .ZN(_0495_));
 AOI21_X1 _1730_ (.A(_0494_),
    .B1(_0495_),
    .B2(_0925_),
    .ZN(_0167_));
 NAND2_X1 _1731_ (.A1(_0850_),
    .A2(net22),
    .ZN(_0496_));
 AOI21_X1 _1732_ (.A(_0456_),
    .B1(_0496_),
    .B2(_0468_),
    .ZN(_0497_));
 MUX2_X1 _1733_ (.A(_0497_),
    .B(_0865_),
    .S(_0920_),
    .Z(_0498_));
 MUX2_X1 _1734_ (.A(net22),
    .B(net10),
    .S(_0484_),
    .Z(_0499_));
 AOI22_X1 _1735_ (.A1(_0478_),
    .A2(_0498_),
    .B1(_0499_),
    .B2(_0490_),
    .ZN(_0500_));
 INV_X1 _1736_ (.A(_0500_),
    .ZN(_0168_));
 AOI21_X1 _1737_ (.A(_0452_),
    .B1(_0448_),
    .B2(net23),
    .ZN(_0501_));
 NOR2_X1 _1738_ (.A1(_0923_),
    .A2(_0501_),
    .ZN(_0502_));
 MUX2_X1 _1739_ (.A(_0502_),
    .B(_0866_),
    .S(_0920_),
    .Z(_0503_));
 NAND2_X1 _1740_ (.A1(_0478_),
    .A2(_0503_),
    .ZN(_0504_));
 MUX2_X1 _1741_ (.A(net23),
    .B(net11),
    .S(_0484_),
    .Z(_0505_));
 NAND3_X1 _1742_ (.A1(_0470_),
    .A2(_0483_),
    .A3(_0505_),
    .ZN(_0506_));
 NAND2_X1 _1743_ (.A1(_0504_),
    .A2(_0506_),
    .ZN(_0169_));
 MUX2_X1 _1744_ (.A(net24),
    .B(net12),
    .S(_0445_),
    .Z(_0507_));
 NAND2_X1 _1745_ (.A1(_0470_),
    .A2(_0507_),
    .ZN(_0508_));
 NAND2_X1 _1746_ (.A1(_0850_),
    .A2(net24),
    .ZN(_0509_));
 AND2_X1 _1747_ (.A1(_0462_),
    .A2(_0509_),
    .ZN(_0510_));
 INV_X1 _1748_ (.A(_0867_),
    .ZN(_0511_));
 AOI221_X2 _1749_ (.A(_0458_),
    .B1(_0508_),
    .B2(_0510_),
    .C1(_0920_),
    .C2(_0511_),
    .ZN(_0170_));
 NAND2_X1 _1750_ (.A1(_0850_),
    .A2(net25),
    .ZN(_0512_));
 AOI21_X1 _1751_ (.A(_0456_),
    .B1(_0512_),
    .B2(_0468_),
    .ZN(_0513_));
 MUX2_X1 _1752_ (.A(_0513_),
    .B(_0868_),
    .S(_0920_),
    .Z(_0514_));
 MUX2_X1 _1753_ (.A(net25),
    .B(net13),
    .S(_0484_),
    .Z(_0515_));
 AOI22_X1 _1754_ (.A1(_0802_),
    .A2(_0514_),
    .B1(_0515_),
    .B2(_0490_),
    .ZN(_0516_));
 INV_X1 _1755_ (.A(_0516_),
    .ZN(_0171_));
 BUF_X2 _1756_ (.A(_1147_),
    .Z(_0517_));
 INV_X1 _1757_ (.A(_0517_),
    .ZN(_0518_));
 NOR4_X1 _1758_ (.A1(_0852_),
    .A2(_0869_),
    .A3(_1148_),
    .A4(_0518_),
    .ZN(_0519_));
 NAND2_X1 _1759_ (.A1(_0848_),
    .A2(_0519_),
    .ZN(_0520_));
 AOI21_X1 _1760_ (.A(_0452_),
    .B1(_0024_),
    .B2(_0520_),
    .ZN(_0521_));
 NOR2_X2 _1761_ (.A1(_0922_),
    .A2(_0902_),
    .ZN(_0522_));
 NAND2_X1 _1762_ (.A1(_0850_),
    .A2(_0818_),
    .ZN(_0523_));
 OAI21_X2 _1763_ (.A(_0886_),
    .B1(_0819_),
    .B2(_0913_),
    .ZN(_0524_));
 NAND3_X2 _1764_ (.A1(_0522_),
    .A2(_0523_),
    .A3(_0524_),
    .ZN(_0525_));
 MUX2_X1 _1765_ (.A(_0521_),
    .B(\bank_active[0] ),
    .S(_0525_),
    .Z(_0526_));
 AND2_X1 _1766_ (.A1(_0803_),
    .A2(_0526_),
    .ZN(_0172_));
 BUF_X2 _1767_ (.A(_0525_),
    .Z(_0527_));
 INV_X1 _1768_ (.A(_0025_),
    .ZN(_0528_));
 XNOR2_X2 _1769_ (.A(_0847_),
    .B(_0517_),
    .ZN(_0529_));
 AOI21_X1 _1770_ (.A(_0528_),
    .B1(_1151_),
    .B2(_0529_),
    .ZN(_0530_));
 NOR3_X1 _1771_ (.A1(_0453_),
    .A2(_0527_),
    .A3(_0530_),
    .ZN(_0531_));
 AOI21_X1 _1772_ (.A(_0531_),
    .B1(_0527_),
    .B2(\bank_active[1] ),
    .ZN(_0532_));
 NOR2_X1 _1773_ (.A1(_0835_),
    .A2(_0532_),
    .ZN(_0173_));
 INV_X1 _1774_ (.A(_0026_),
    .ZN(_0533_));
 AOI21_X1 _1775_ (.A(_0533_),
    .B1(_1149_),
    .B2(_0529_),
    .ZN(_0534_));
 NOR3_X1 _1776_ (.A1(_0453_),
    .A2(_0527_),
    .A3(_0534_),
    .ZN(_0535_));
 AOI21_X1 _1777_ (.A(_0535_),
    .B1(_0527_),
    .B2(\bank_active[2] ),
    .ZN(_0536_));
 NOR2_X1 _1778_ (.A1(_0835_),
    .A2(_0536_),
    .ZN(_0174_));
 INV_X1 _1779_ (.A(_0027_),
    .ZN(_0537_));
 AOI21_X1 _1780_ (.A(_0537_),
    .B1(_1153_),
    .B2(_0529_),
    .ZN(_0538_));
 NOR3_X1 _1781_ (.A1(_0453_),
    .A2(_0527_),
    .A3(_0538_),
    .ZN(_0539_));
 AOI21_X1 _1782_ (.A(_0539_),
    .B1(_0527_),
    .B2(\bank_active[3] ),
    .ZN(_0540_));
 NOR2_X1 _1783_ (.A1(_0835_),
    .A2(_0540_),
    .ZN(_0175_));
 AND3_X1 _1784_ (.A1(_0848_),
    .A2(_0852_),
    .A3(_0518_),
    .ZN(_0541_));
 AOI21_X1 _1785_ (.A(_0541_),
    .B1(_0517_),
    .B2(_0847_),
    .ZN(_0542_));
 OR3_X1 _1786_ (.A1(_0869_),
    .A2(_1148_),
    .A3(_0542_),
    .ZN(_0543_));
 AOI21_X1 _1787_ (.A(_0452_),
    .B1(_0028_),
    .B2(_0543_),
    .ZN(_0544_));
 MUX2_X1 _1788_ (.A(_0544_),
    .B(\bank_active[4] ),
    .S(_0525_),
    .Z(_0545_));
 AND2_X1 _1789_ (.A1(_0803_),
    .A2(_0545_),
    .ZN(_0176_));
 INV_X1 _1790_ (.A(_0029_),
    .ZN(_0546_));
 XOR2_X2 _1791_ (.A(_0847_),
    .B(_0517_),
    .Z(_0547_));
 AOI21_X1 _1792_ (.A(_0546_),
    .B1(_1151_),
    .B2(_0547_),
    .ZN(_0548_));
 NOR3_X1 _1793_ (.A1(_0453_),
    .A2(_0527_),
    .A3(_0548_),
    .ZN(_0549_));
 AOI21_X1 _1794_ (.A(_0549_),
    .B1(_0527_),
    .B2(\bank_active[5] ),
    .ZN(_0550_));
 NOR2_X1 _1795_ (.A1(_0835_),
    .A2(_0550_),
    .ZN(_0177_));
 INV_X1 _1796_ (.A(_0030_),
    .ZN(_0551_));
 AOI21_X1 _1797_ (.A(_0551_),
    .B1(_1149_),
    .B2(_0547_),
    .ZN(_0552_));
 NOR3_X1 _1798_ (.A1(_0452_),
    .A2(_0525_),
    .A3(_0552_),
    .ZN(_0553_));
 AOI21_X1 _1799_ (.A(_0553_),
    .B1(_0527_),
    .B2(\bank_active[6] ),
    .ZN(_0554_));
 NOR2_X1 _1800_ (.A1(_0835_),
    .A2(_0554_),
    .ZN(_0178_));
 INV_X1 _1801_ (.A(_0031_),
    .ZN(_0555_));
 AOI21_X1 _1802_ (.A(_0555_),
    .B1(_1153_),
    .B2(_0547_),
    .ZN(_0556_));
 NOR3_X1 _1803_ (.A1(_0452_),
    .A2(_0525_),
    .A3(_0556_),
    .ZN(_0557_));
 AOI21_X1 _1804_ (.A(_0557_),
    .B1(_0527_),
    .B2(\bank_active[7] ),
    .ZN(_0558_));
 NOR2_X1 _1805_ (.A1(_0835_),
    .A2(_0558_),
    .ZN(_0179_));
 MUX2_X1 _1806_ (.A(_0828_),
    .B(_0934_),
    .S(_0447_),
    .Z(_0559_));
 OAI21_X2 _1807_ (.A(_0908_),
    .B1(_0447_),
    .B2(_0923_),
    .ZN(_0560_));
 MUX2_X1 _1808_ (.A(_0559_),
    .B(net115),
    .S(_0560_),
    .Z(_0561_));
 AND2_X1 _1809_ (.A1(_0803_),
    .A2(_0561_),
    .ZN(_0180_));
 NAND2_X1 _1810_ (.A1(_0852_),
    .A2(_0560_),
    .ZN(_0562_));
 NOR3_X1 _1811_ (.A1(_0824_),
    .A2(_0447_),
    .A3(_0828_),
    .ZN(_0563_));
 AOI21_X1 _1812_ (.A(_0563_),
    .B1(_0930_),
    .B2(_0470_),
    .ZN(_0564_));
 OR2_X1 _1813_ (.A1(_0560_),
    .A2(_0564_),
    .ZN(_0565_));
 AOI21_X1 _1814_ (.A(_0834_),
    .B1(_0562_),
    .B2(_0565_),
    .ZN(_0181_));
 NAND2_X1 _1815_ (.A1(_0847_),
    .A2(_0560_),
    .ZN(_0566_));
 NAND3_X1 _1816_ (.A1(_0470_),
    .A2(_0295_),
    .A3(_0908_),
    .ZN(_0567_));
 AOI21_X1 _1817_ (.A(_0834_),
    .B1(_0566_),
    .B2(_0567_),
    .ZN(_0182_));
 MUX2_X1 _1818_ (.A(net26),
    .B(_1155_),
    .S(_0886_),
    .Z(_0568_));
 AOI22_X1 _1819_ (.A1(_0887_),
    .A2(_0523_),
    .B1(_0913_),
    .B2(_0872_),
    .ZN(_0569_));
 OR3_X2 _1820_ (.A1(_0922_),
    .A2(_0907_),
    .A3(_0569_),
    .ZN(_0570_));
 AOI21_X2 _1821_ (.A(_0570_),
    .B1(_0484_),
    .B2(_0447_),
    .ZN(_0571_));
 MUX2_X1 _1822_ (.A(\burst_counter[0] ),
    .B(_0568_),
    .S(_0571_),
    .Z(_0572_));
 AND2_X1 _1823_ (.A1(_0478_),
    .A2(_0572_),
    .ZN(_0183_));
 NOR2_X1 _1824_ (.A1(_0452_),
    .A2(net27),
    .ZN(_0573_));
 AOI21_X1 _1825_ (.A(_0573_),
    .B1(_1158_),
    .B2(_0452_),
    .ZN(_0574_));
 MUX2_X1 _1826_ (.A(\burst_counter[1] ),
    .B(_0574_),
    .S(_0571_),
    .Z(_0575_));
 AND2_X1 _1827_ (.A1(_0478_),
    .A2(_0575_),
    .ZN(_0184_));
 INV_X1 _1828_ (.A(_1159_),
    .ZN(_0576_));
 AOI221_X1 _1829_ (.A(_0570_),
    .B1(_0576_),
    .B2(_0886_),
    .C1(_0447_),
    .C2(_0484_),
    .ZN(_0577_));
 AND2_X1 _1830_ (.A1(_0888_),
    .A2(net28),
    .ZN(_0578_));
 NOR3_X1 _1831_ (.A1(_0888_),
    .A2(\burst_counter[2] ),
    .A3(_0576_),
    .ZN(_0579_));
 OAI21_X1 _1832_ (.A(_0802_),
    .B1(_0578_),
    .B2(_0579_),
    .ZN(_0580_));
 OAI33_X1 _1833_ (.A1(_0834_),
    .A2(_0912_),
    .A3(_0577_),
    .B1(_0580_),
    .B2(_0454_),
    .B3(_0570_),
    .ZN(_0185_));
 NAND2_X1 _1834_ (.A1(_0802_),
    .A2(\burst_counter[3] ),
    .ZN(_0581_));
 NOR3_X2 _1835_ (.A1(\burst_counter[2] ),
    .A2(\burst_counter[1] ),
    .A3(\burst_counter[0] ),
    .ZN(_0582_));
 NAND4_X1 _1836_ (.A1(_0802_),
    .A2(_0452_),
    .A3(_0911_),
    .A4(_0582_),
    .ZN(_0583_));
 MUX2_X1 _1837_ (.A(_0581_),
    .B(_0583_),
    .S(_0571_),
    .Z(_0584_));
 NAND4_X1 _1838_ (.A1(_0802_),
    .A2(_0888_),
    .A3(net29),
    .A4(_0571_),
    .ZN(_0585_));
 NAND3_X1 _1839_ (.A1(_0802_),
    .A2(_0453_),
    .A3(\burst_counter[3] ),
    .ZN(_0586_));
 OAI211_X2 _1840_ (.A(_0584_),
    .B(_0585_),
    .C1(_0586_),
    .C2(_0582_),
    .ZN(_0186_));
 INV_X1 _1841_ (.A(net30),
    .ZN(_0587_));
 NAND2_X1 _1842_ (.A1(_0904_),
    .A2(_0872_),
    .ZN(_0588_));
 NOR3_X2 _1843_ (.A1(_0587_),
    .A2(_0588_),
    .A3(_0445_),
    .ZN(_0589_));
 AOI21_X1 _1844_ (.A(_0903_),
    .B1(_1162_),
    .B2(_0589_),
    .ZN(_0590_));
 OAI21_X2 _1845_ (.A(_0850_),
    .B1(_0587_),
    .B2(_0819_),
    .ZN(_0591_));
 INV_X1 _1846_ (.A(_0591_),
    .ZN(_0592_));
 NAND3_X2 _1847_ (.A1(_0887_),
    .A2(_0851_),
    .A3(_0522_),
    .ZN(_0593_));
 NAND2_X1 _1848_ (.A1(_0801_),
    .A2(_0593_),
    .ZN(_0594_));
 OR2_X1 _1849_ (.A1(_0901_),
    .A2(_0594_),
    .ZN(_0595_));
 OR4_X1 _1850_ (.A1(_0915_),
    .A2(_0590_),
    .A3(_0592_),
    .A4(_0595_),
    .ZN(_0187_));
 NOR3_X1 _1851_ (.A1(_0453_),
    .A2(_0910_),
    .A3(_0595_),
    .ZN(_0596_));
 NOR4_X4 _1852_ (.A1(\refresh_counter[15] ),
    .A2(\refresh_counter[14] ),
    .A3(\refresh_counter[11] ),
    .A4(_0838_),
    .ZN(_0597_));
 OR2_X1 _1853_ (.A1(\refresh_counter[6] ),
    .A2(_0840_),
    .ZN(_0598_));
 AND3_X1 _1854_ (.A1(\refresh_counter[3] ),
    .A2(\refresh_counter[2] ),
    .A3(\refresh_counter[4] ),
    .ZN(_0599_));
 OR2_X1 _1855_ (.A1(_1167_),
    .A2(_1165_),
    .ZN(_0600_));
 AOI21_X2 _1856_ (.A(_0598_),
    .B1(_0599_),
    .B2(_0600_),
    .ZN(_0601_));
 NAND4_X2 _1857_ (.A1(\refresh_counter[7] ),
    .A2(\refresh_counter[10] ),
    .A3(\refresh_counter[9] ),
    .A4(\refresh_counter[8] ),
    .ZN(_0602_));
 OAI211_X4 _1858_ (.A(_0902_),
    .B(_0597_),
    .C1(_0601_),
    .C2(_0602_),
    .ZN(_0603_));
 NOR2_X1 _1859_ (.A1(_0588_),
    .A2(_0484_),
    .ZN(_0604_));
 OAI21_X1 _1860_ (.A(_0596_),
    .B1(_0603_),
    .B2(_0604_),
    .ZN(_0188_));
 AOI21_X1 _1861_ (.A(_0603_),
    .B1(_0484_),
    .B2(_0906_),
    .ZN(_0605_));
 OR4_X1 _1862_ (.A1(_0448_),
    .A2(_0915_),
    .A3(_0595_),
    .A4(_0605_),
    .ZN(_0189_));
 AND2_X1 _1863_ (.A1(_0851_),
    .A2(_1183_),
    .ZN(_0606_));
 OAI21_X1 _1864_ (.A(_0606_),
    .B1(_0484_),
    .B2(_0903_),
    .ZN(_0607_));
 OAI21_X1 _1865_ (.A(_0836_),
    .B1(_0032_),
    .B2(_0872_),
    .ZN(_0608_));
 AOI21_X1 _1866_ (.A(_0907_),
    .B1(_0608_),
    .B2(_0922_),
    .ZN(_0609_));
 NAND2_X1 _1867_ (.A1(_0916_),
    .A2(_0609_),
    .ZN(_0610_));
 MUX2_X1 _1868_ (.A(_0607_),
    .B(net196),
    .S(_0610_),
    .Z(_0611_));
 AND2_X1 _1869_ (.A1(_0478_),
    .A2(_0611_),
    .ZN(_0190_));
 MUX2_X1 _1870_ (.A(_1183_),
    .B(net197),
    .S(_0610_),
    .Z(_0612_));
 AND2_X1 _1871_ (.A1(_0478_),
    .A2(_0612_),
    .ZN(_0191_));
 AOI21_X1 _1872_ (.A(net100),
    .B1(_0821_),
    .B2(_0836_),
    .ZN(_0613_));
 NOR2_X1 _1873_ (.A1(_0835_),
    .A2(_0613_),
    .ZN(_0192_));
 NAND2_X1 _1874_ (.A1(_0478_),
    .A2(_0453_),
    .ZN(_0614_));
 CLKBUF_X3 _1875_ (.A(_0872_),
    .Z(_0615_));
 AOI21_X1 _1876_ (.A(_0891_),
    .B1(_0913_),
    .B2(net32),
    .ZN(_0616_));
 OR3_X2 _1877_ (.A1(\timer[2] ),
    .A2(_0808_),
    .A3(_0816_),
    .ZN(_0617_));
 NAND4_X1 _1878_ (.A1(_0889_),
    .A2(_0890_),
    .A3(net128),
    .A4(_1178_),
    .ZN(_0618_));
 NOR2_X1 _1879_ (.A1(_0617_),
    .A2(_0618_),
    .ZN(_0619_));
 BUF_X1 _1880_ (.A(_1175_),
    .Z(_0620_));
 AND2_X1 _1881_ (.A1(_0620_),
    .A2(_0809_),
    .ZN(_0621_));
 OR3_X2 _1882_ (.A1(_0816_),
    .A2(_0891_),
    .A3(_0621_),
    .ZN(_0622_));
 AND2_X1 _1883_ (.A1(_0810_),
    .A2(_0622_),
    .ZN(_0623_));
 AOI22_X1 _1884_ (.A1(_0615_),
    .A2(_0616_),
    .B1(_0619_),
    .B2(_0623_),
    .ZN(_0624_));
 NOR2_X1 _1885_ (.A1(_0614_),
    .A2(_0624_),
    .ZN(_0257_));
 AOI21_X1 _1886_ (.A(_0806_),
    .B1(_0836_),
    .B2(_0872_),
    .ZN(_0625_));
 NOR2_X1 _1887_ (.A1(_0522_),
    .A2(_0625_),
    .ZN(_0626_));
 NOR2_X1 _1888_ (.A1(_1164_),
    .A2(_0626_),
    .ZN(_0627_));
 AOI21_X1 _1889_ (.A(_0627_),
    .B1(_1163_),
    .B2(_0470_),
    .ZN(_0628_));
 NOR2_X1 _1890_ (.A1(_0835_),
    .A2(_0628_),
    .ZN(_0258_));
 NAND2_X1 _1891_ (.A1(_0603_),
    .A2(_0626_),
    .ZN(_0629_));
 NAND2_X2 _1892_ (.A1(_0801_),
    .A2(_0629_),
    .ZN(_0630_));
 CLKBUF_X3 _1893_ (.A(_0630_),
    .Z(_0631_));
 AND2_X1 _1894_ (.A1(_1167_),
    .A2(_1162_),
    .ZN(_0632_));
 AND4_X1 _1895_ (.A1(\refresh_counter[7] ),
    .A2(\refresh_counter[6] ),
    .A3(_0840_),
    .A4(_0599_),
    .ZN(_0633_));
 AND2_X1 _1896_ (.A1(_0632_),
    .A2(_0633_),
    .ZN(_0634_));
 NAND3_X1 _1897_ (.A1(\refresh_counter[9] ),
    .A2(\refresh_counter[8] ),
    .A3(_0634_),
    .ZN(_0635_));
 XNOR2_X1 _1898_ (.A(_0042_),
    .B(_0635_),
    .ZN(_0636_));
 NOR2_X1 _1899_ (.A1(_0631_),
    .A2(_0636_),
    .ZN(_0259_));
 NOR2_X1 _1900_ (.A1(_0043_),
    .A2(_0631_),
    .ZN(_0260_));
 NOR2_X1 _1901_ (.A1(_0044_),
    .A2(_0630_),
    .ZN(_0261_));
 NOR2_X1 _1902_ (.A1(_0045_),
    .A2(_0630_),
    .ZN(_0262_));
 NOR2_X1 _1903_ (.A1(_0008_),
    .A2(_0630_),
    .ZN(_0263_));
 NOR2_X1 _1904_ (.A1(_0009_),
    .A2(_0630_),
    .ZN(_0264_));
 MUX2_X1 _1905_ (.A(_0033_),
    .B(_1166_),
    .S(_1162_),
    .Z(_0637_));
 NOR2_X1 _1906_ (.A1(_0631_),
    .A2(_0637_),
    .ZN(_0265_));
 OR2_X1 _1907_ (.A1(_0034_),
    .A2(_0632_),
    .ZN(_0638_));
 NAND2_X1 _1908_ (.A1(_0034_),
    .A2(_0632_),
    .ZN(_0639_));
 AOI21_X1 _1909_ (.A(_0630_),
    .B1(_0638_),
    .B2(_0639_),
    .ZN(_0266_));
 AND3_X1 _1910_ (.A1(\refresh_counter[1] ),
    .A2(\refresh_counter[0] ),
    .A3(_1162_),
    .ZN(_0640_));
 NAND2_X1 _1911_ (.A1(\refresh_counter[2] ),
    .A2(_0640_),
    .ZN(_0641_));
 XNOR2_X1 _1912_ (.A(_0035_),
    .B(_0641_),
    .ZN(_0642_));
 NOR2_X1 _1913_ (.A1(_0631_),
    .A2(_0642_),
    .ZN(_0267_));
 NAND3_X1 _1914_ (.A1(\refresh_counter[3] ),
    .A2(\refresh_counter[2] ),
    .A3(_0632_),
    .ZN(_0643_));
 XNOR2_X1 _1915_ (.A(_0036_),
    .B(_0643_),
    .ZN(_0644_));
 NOR2_X1 _1916_ (.A1(_0631_),
    .A2(_0644_),
    .ZN(_0268_));
 NAND2_X1 _1917_ (.A1(_0599_),
    .A2(_0640_),
    .ZN(_0645_));
 XNOR2_X1 _1918_ (.A(_0037_),
    .B(_0645_),
    .ZN(_0646_));
 NOR2_X1 _1919_ (.A1(_0631_),
    .A2(_0646_),
    .ZN(_0269_));
 NAND3_X1 _1920_ (.A1(_0840_),
    .A2(_0599_),
    .A3(_0632_),
    .ZN(_0647_));
 XNOR2_X1 _1921_ (.A(_0038_),
    .B(_0647_),
    .ZN(_0648_));
 NOR2_X1 _1922_ (.A1(_0631_),
    .A2(_0648_),
    .ZN(_0270_));
 NAND4_X1 _1923_ (.A1(\refresh_counter[6] ),
    .A2(_0840_),
    .A3(_0599_),
    .A4(_0640_),
    .ZN(_0649_));
 XNOR2_X1 _1924_ (.A(_0039_),
    .B(_0649_),
    .ZN(_0650_));
 NOR2_X1 _1925_ (.A1(_0631_),
    .A2(_0650_),
    .ZN(_0271_));
 XOR2_X1 _1926_ (.A(_0040_),
    .B(_0634_),
    .Z(_0651_));
 NOR2_X1 _1927_ (.A1(_0631_),
    .A2(_0651_),
    .ZN(_0272_));
 NAND3_X1 _1928_ (.A1(\refresh_counter[8] ),
    .A2(_0633_),
    .A3(_0640_),
    .ZN(_0652_));
 XNOR2_X1 _1929_ (.A(_0041_),
    .B(_0652_),
    .ZN(_0653_));
 NOR2_X1 _1930_ (.A1(_0631_),
    .A2(_0653_),
    .ZN(_0273_));
 NOR2_X1 _1931_ (.A1(\init_state[4] ),
    .A2(_0823_),
    .ZN(_0654_));
 NOR4_X4 _1932_ (.A1(\init_state[2] ),
    .A2(_0824_),
    .A3(_0828_),
    .A4(\init_state[6] ),
    .ZN(_0655_));
 NAND2_X2 _1933_ (.A1(_0654_),
    .A2(_0655_),
    .ZN(_0656_));
 NOR2_X1 _1934_ (.A1(_0826_),
    .A2(_0656_),
    .ZN(_0657_));
 NAND2_X1 _1935_ (.A1(_0922_),
    .A2(_1171_),
    .ZN(_0658_));
 OAI221_X1 _1936_ (.A(_0593_),
    .B1(_0657_),
    .B2(_0658_),
    .C1(_1173_),
    .C2(_0851_),
    .ZN(_0659_));
 NOR3_X2 _1937_ (.A1(_0816_),
    .A2(_0891_),
    .A3(_0621_),
    .ZN(_0660_));
 NAND2_X1 _1938_ (.A1(_0889_),
    .A2(net128),
    .ZN(_0661_));
 INV_X1 _1939_ (.A(_0890_),
    .ZN(_0662_));
 NAND2_X1 _1940_ (.A1(_0662_),
    .A2(net98),
    .ZN(_0663_));
 NAND3_X2 _1941_ (.A1(_0890_),
    .A2(net32),
    .A3(net195),
    .ZN(_0664_));
 AOI21_X4 _1942_ (.A(_0661_),
    .B1(_0663_),
    .B2(_0664_),
    .ZN(_0665_));
 MUX2_X1 _1943_ (.A(_1172_),
    .B(_0914_),
    .S(_0665_),
    .Z(_0666_));
 OR3_X1 _1944_ (.A1(_0619_),
    .A2(_0660_),
    .A3(_0666_),
    .ZN(_0667_));
 OAI21_X1 _1945_ (.A(_0667_),
    .B1(_0622_),
    .B2(\timer[0] ),
    .ZN(_0668_));
 NOR2_X1 _1946_ (.A1(_0888_),
    .A2(_0872_),
    .ZN(_0669_));
 OAI33_X1 _1947_ (.A1(_0888_),
    .A2(_0819_),
    .A3(_0914_),
    .B1(_0656_),
    .B2(_0826_),
    .B3(_0805_),
    .ZN(_0670_));
 INV_X1 _1948_ (.A(_1172_),
    .ZN(_0671_));
 AOI221_X1 _1949_ (.A(_0659_),
    .B1(_0668_),
    .B2(_0669_),
    .C1(_0670_),
    .C2(_0671_),
    .ZN(_0672_));
 OAI21_X1 _1950_ (.A(_0605_),
    .B1(_0906_),
    .B2(_0671_),
    .ZN(_0673_));
 AOI221_X1 _1951_ (.A(_0834_),
    .B1(_1172_),
    .B2(_0909_),
    .C1(_0672_),
    .C2(_0673_),
    .ZN(_0274_));
 AOI21_X2 _1952_ (.A(_0909_),
    .B1(_0657_),
    .B2(_0922_),
    .ZN(_0674_));
 AND2_X1 _1953_ (.A1(_0902_),
    .A2(_1162_),
    .ZN(_0675_));
 NOR2_X1 _1954_ (.A1(_0904_),
    .A2(_0603_),
    .ZN(_0676_));
 OAI22_X1 _1955_ (.A1(_0922_),
    .A2(_0675_),
    .B1(_0676_),
    .B2(_0818_),
    .ZN(_0677_));
 NAND2_X1 _1956_ (.A1(_0674_),
    .A2(_0677_),
    .ZN(_0678_));
 NOR2_X1 _1957_ (.A1(_0816_),
    .A2(_0618_),
    .ZN(_0679_));
 OAI221_X2 _1958_ (.A(_0622_),
    .B1(_0665_),
    .B2(_0679_),
    .C1(_0816_),
    .C2(_0810_),
    .ZN(_0680_));
 AND2_X1 _1959_ (.A1(_0915_),
    .A2(_0680_),
    .ZN(_0681_));
 OR2_X1 _1960_ (.A1(_0678_),
    .A2(_0681_),
    .ZN(_0682_));
 OAI21_X4 _1961_ (.A(_0801_),
    .B1(_0910_),
    .B2(_0682_),
    .ZN(_0683_));
 OR2_X1 _1962_ (.A1(_0813_),
    .A2(_0814_),
    .ZN(_0684_));
 NOR2_X1 _1963_ (.A1(_0810_),
    .A2(_0684_),
    .ZN(_0685_));
 OAI21_X2 _1964_ (.A(_0685_),
    .B1(_0812_),
    .B2(_0811_),
    .ZN(_0686_));
 XNOR2_X1 _1965_ (.A(_0018_),
    .B(_0686_),
    .ZN(_0687_));
 NOR2_X1 _1966_ (.A1(_0683_),
    .A2(_0687_),
    .ZN(_0275_));
 INV_X1 _1967_ (.A(_0808_),
    .ZN(_0688_));
 NOR3_X2 _1968_ (.A1(\timer[2] ),
    .A2(\timer[0] ),
    .A3(\timer[1] ),
    .ZN(_0689_));
 NAND2_X2 _1969_ (.A1(_0688_),
    .A2(_0689_),
    .ZN(_0690_));
 NOR4_X1 _1970_ (.A1(\timer[10] ),
    .A2(_0684_),
    .A3(_0615_),
    .A4(_0690_),
    .ZN(_0691_));
 XOR2_X1 _1971_ (.A(_0019_),
    .B(_0691_),
    .Z(_0692_));
 NOR2_X1 _1972_ (.A1(_0683_),
    .A2(_0692_),
    .ZN(_0276_));
 NOR3_X1 _1973_ (.A1(\timer[11] ),
    .A2(\timer[10] ),
    .A3(_0686_),
    .ZN(_0693_));
 XOR2_X1 _1974_ (.A(_0020_),
    .B(_0693_),
    .Z(_0694_));
 NOR2_X1 _1975_ (.A1(_0683_),
    .A2(_0694_),
    .ZN(_0277_));
 OAI21_X1 _1976_ (.A(_0615_),
    .B1(_0915_),
    .B2(_0678_),
    .ZN(_0695_));
 NOR4_X1 _1977_ (.A1(_0021_),
    .A2(_0811_),
    .A3(_0684_),
    .A4(_0690_),
    .ZN(_0696_));
 OR4_X1 _1978_ (.A1(_0811_),
    .A2(_0684_),
    .A3(_0872_),
    .A4(_0690_),
    .ZN(_0697_));
 AOI221_X1 _1979_ (.A(_0683_),
    .B1(_0695_),
    .B2(_0696_),
    .C1(_0697_),
    .C2(_0021_),
    .ZN(_0278_));
 NOR3_X1 _1980_ (.A1(\timer[13] ),
    .A2(_0811_),
    .A3(_0686_),
    .ZN(_0698_));
 XOR2_X1 _1981_ (.A(_0022_),
    .B(_0698_),
    .Z(_0699_));
 NOR2_X1 _1982_ (.A1(_0683_),
    .A2(_0699_),
    .ZN(_0279_));
 NOR3_X1 _1983_ (.A1(\timer[13] ),
    .A2(\timer[14] ),
    .A3(_0697_),
    .ZN(_0700_));
 XOR2_X1 _1984_ (.A(_0023_),
    .B(_0700_),
    .Z(_0701_));
 NOR2_X1 _1985_ (.A1(_0683_),
    .A2(_0701_),
    .ZN(_0280_));
 MUX2_X1 _1986_ (.A(_0620_),
    .B(_1177_),
    .S(_0820_),
    .Z(_0702_));
 AOI21_X1 _1987_ (.A(_0834_),
    .B1(_0909_),
    .B2(_0702_),
    .ZN(_0703_));
 NAND2_X1 _1988_ (.A1(_0831_),
    .A2(_0654_),
    .ZN(_0704_));
 OAI21_X1 _1989_ (.A(_0655_),
    .B1(_0704_),
    .B2(_0620_),
    .ZN(_0705_));
 OAI21_X1 _1990_ (.A(_0922_),
    .B1(_0820_),
    .B2(_0705_),
    .ZN(_0706_));
 AOI22_X1 _1991_ (.A1(_1177_),
    .A2(_0820_),
    .B1(_0591_),
    .B2(_0706_),
    .ZN(_0707_));
 NOR2_X1 _1992_ (.A1(_0909_),
    .A2(_0707_),
    .ZN(_0708_));
 NOR2_X1 _1993_ (.A1(_0904_),
    .A2(_0819_),
    .ZN(_0709_));
 AOI221_X1 _1994_ (.A(_0603_),
    .B1(_0709_),
    .B2(_0620_),
    .C1(_1177_),
    .C2(_0819_),
    .ZN(_0710_));
 INV_X1 _1995_ (.A(_0710_),
    .ZN(_0711_));
 NOR2_X1 _1996_ (.A1(_0665_),
    .A2(_0679_),
    .ZN(_0712_));
 NOR2_X1 _1997_ (.A1(_0660_),
    .A2(_0712_),
    .ZN(_0713_));
 OAI21_X1 _1998_ (.A(_1170_),
    .B1(_0713_),
    .B2(_1177_),
    .ZN(_0714_));
 NAND3_X1 _1999_ (.A1(_0620_),
    .A2(_0615_),
    .A3(_0913_),
    .ZN(_0715_));
 NAND2_X1 _2000_ (.A1(_0714_),
    .A2(_0715_),
    .ZN(_0716_));
 OAI221_X1 _2001_ (.A(_0708_),
    .B1(_0711_),
    .B2(_0589_),
    .C1(_0888_),
    .C2(_0716_),
    .ZN(_0717_));
 AND2_X1 _2002_ (.A1(_0703_),
    .A2(_0717_),
    .ZN(_0281_));
 NAND3_X1 _2003_ (.A1(_0470_),
    .A2(_0587_),
    .A3(_0604_),
    .ZN(_0718_));
 INV_X1 _2004_ (.A(_0010_),
    .ZN(_0719_));
 OAI21_X1 _2005_ (.A(_0807_),
    .B1(_0593_),
    .B2(_0617_),
    .ZN(_0720_));
 NOR2_X1 _2006_ (.A1(_0719_),
    .A2(_0720_),
    .ZN(_0721_));
 NAND2_X1 _2007_ (.A1(_0807_),
    .A2(_0617_),
    .ZN(_0722_));
 AOI21_X1 _2008_ (.A(_0721_),
    .B1(_0722_),
    .B2(_0719_),
    .ZN(_0723_));
 NAND2_X1 _2009_ (.A1(_0593_),
    .A2(_0591_),
    .ZN(_0724_));
 NAND2_X1 _2010_ (.A1(_0010_),
    .A2(_0615_),
    .ZN(_0725_));
 AOI21_X1 _2011_ (.A(_0724_),
    .B1(_0725_),
    .B2(_0681_),
    .ZN(_0726_));
 NOR3_X1 _2012_ (.A1(_0719_),
    .A2(_0617_),
    .A3(_0656_),
    .ZN(_0727_));
 AOI21_X1 _2013_ (.A(_0727_),
    .B1(_0656_),
    .B2(_0872_),
    .ZN(_0728_));
 OAI21_X1 _2014_ (.A(_0923_),
    .B1(_0826_),
    .B2(_0728_),
    .ZN(_0729_));
 AOI21_X1 _2015_ (.A(_0723_),
    .B1(_0726_),
    .B2(_0729_),
    .ZN(_0730_));
 NAND2_X1 _2016_ (.A1(_0010_),
    .A2(_0722_),
    .ZN(_0731_));
 OAI21_X1 _2017_ (.A(_0807_),
    .B1(_0904_),
    .B2(_0617_),
    .ZN(_0732_));
 OAI21_X1 _2018_ (.A(_0731_),
    .B1(_0732_),
    .B2(_0010_),
    .ZN(_0733_));
 NAND2_X1 _2019_ (.A1(_1162_),
    .A2(_0733_),
    .ZN(_0734_));
 AOI21_X1 _2020_ (.A(_0730_),
    .B1(_0734_),
    .B2(_0470_),
    .ZN(_0735_));
 AOI21_X1 _2021_ (.A(_0834_),
    .B1(_0718_),
    .B2(_0735_),
    .ZN(_0282_));
 AOI21_X1 _2022_ (.A(_0922_),
    .B1(_0819_),
    .B2(_0909_),
    .ZN(_0736_));
 NOR2_X1 _2023_ (.A1(_0819_),
    .A2(_0656_),
    .ZN(_0737_));
 OAI221_X1 _2024_ (.A(_0591_),
    .B1(_0736_),
    .B2(_0737_),
    .C1(_0674_),
    .C2(_0011_),
    .ZN(_0738_));
 NAND3_X1 _2025_ (.A1(_0011_),
    .A2(_0872_),
    .A3(_0913_),
    .ZN(_0739_));
 AND2_X1 _2026_ (.A1(_0886_),
    .A2(_0739_),
    .ZN(_0740_));
 AOI21_X1 _2027_ (.A(_0738_),
    .B1(_0740_),
    .B2(_0680_),
    .ZN(_0741_));
 OAI21_X1 _2028_ (.A(_0011_),
    .B1(_0909_),
    .B2(_0905_),
    .ZN(_0742_));
 OAI21_X1 _2029_ (.A(_0675_),
    .B1(_0742_),
    .B2(_0820_),
    .ZN(_0743_));
 OR2_X1 _2030_ (.A1(_0589_),
    .A2(_0743_),
    .ZN(_0744_));
 XNOR2_X1 _2031_ (.A(_0808_),
    .B(_0689_),
    .ZN(_0745_));
 AOI221_X1 _2032_ (.A(_0834_),
    .B1(_0741_),
    .B2(_0744_),
    .C1(_0745_),
    .C2(_1170_),
    .ZN(_0283_));
 XOR2_X1 _2033_ (.A(_0012_),
    .B(_0810_),
    .Z(_0746_));
 NAND2_X1 _2034_ (.A1(_0522_),
    .A2(_0674_),
    .ZN(_0747_));
 OAI21_X1 _2035_ (.A(_0851_),
    .B1(_0524_),
    .B2(_0713_),
    .ZN(_0748_));
 OAI221_X1 _2036_ (.A(_0746_),
    .B1(_0747_),
    .B2(_0748_),
    .C1(_0810_),
    .C2(_0816_),
    .ZN(_0749_));
 OR2_X1 _2037_ (.A1(_0012_),
    .A2(_0820_),
    .ZN(_0750_));
 AOI21_X1 _2038_ (.A(_0750_),
    .B1(_0674_),
    .B2(_0524_),
    .ZN(_0751_));
 OAI21_X1 _2039_ (.A(_1162_),
    .B1(_0750_),
    .B2(_0904_),
    .ZN(_0752_));
 AOI21_X1 _2040_ (.A(_0751_),
    .B1(_0752_),
    .B2(_0470_),
    .ZN(_0753_));
 AOI21_X1 _2041_ (.A(_0834_),
    .B1(_0749_),
    .B2(_0753_),
    .ZN(_0284_));
 NOR2_X1 _2042_ (.A1(\timer[4] ),
    .A2(_0690_),
    .ZN(_0754_));
 XNOR2_X1 _2043_ (.A(_0013_),
    .B(_0754_),
    .ZN(_0755_));
 NAND3_X1 _2044_ (.A1(_0806_),
    .A2(_0593_),
    .A3(_0603_),
    .ZN(_0756_));
 OAI21_X1 _2045_ (.A(_0755_),
    .B1(_0756_),
    .B2(_0748_),
    .ZN(_0757_));
 OAI21_X1 _2046_ (.A(_0831_),
    .B1(_0013_),
    .B2(_0656_),
    .ZN(_0758_));
 AOI21_X1 _2047_ (.A(_1170_),
    .B1(_0758_),
    .B2(_0923_),
    .ZN(_0759_));
 NOR3_X1 _2048_ (.A1(_0909_),
    .A2(_0915_),
    .A3(_0676_),
    .ZN(_0760_));
 OR2_X1 _2049_ (.A1(_0013_),
    .A2(_0760_),
    .ZN(_0761_));
 AOI221_X1 _2050_ (.A(_0833_),
    .B1(_1170_),
    .B2(_0757_),
    .C1(_0759_),
    .C2(_0761_),
    .ZN(_0285_));
 NAND2_X1 _2051_ (.A1(_0819_),
    .A2(_0660_),
    .ZN(_0762_));
 OAI21_X1 _2052_ (.A(_0762_),
    .B1(_0820_),
    .B2(_0014_),
    .ZN(_0763_));
 AOI22_X1 _2053_ (.A1(_0923_),
    .A2(_0704_),
    .B1(_0763_),
    .B2(_0915_),
    .ZN(_0764_));
 NOR2_X1 _2054_ (.A1(_0594_),
    .A2(_0764_),
    .ZN(_0765_));
 OAI21_X1 _2055_ (.A(_0851_),
    .B1(_0655_),
    .B2(_0806_),
    .ZN(_0766_));
 NAND2_X1 _2056_ (.A1(_0820_),
    .A2(_0766_),
    .ZN(_0767_));
 NOR4_X1 _2057_ (.A1(_0524_),
    .A2(_0619_),
    .A3(_0660_),
    .A4(_0665_),
    .ZN(_0768_));
 AOI21_X1 _2058_ (.A(_0768_),
    .B1(_0675_),
    .B2(_0588_),
    .ZN(_0769_));
 NAND3_X1 _2059_ (.A1(_0674_),
    .A2(_0767_),
    .A3(_0769_),
    .ZN(_0770_));
 AOI21_X1 _2060_ (.A(_0765_),
    .B1(_0770_),
    .B2(_0802_),
    .ZN(_0771_));
 NOR3_X1 _2061_ (.A1(\timer[5] ),
    .A2(\timer[4] ),
    .A3(_0810_),
    .ZN(_0772_));
 NAND2_X1 _2062_ (.A1(_1170_),
    .A2(_0772_),
    .ZN(_0773_));
 NAND2_X1 _2063_ (.A1(_0014_),
    .A2(_0773_),
    .ZN(_0774_));
 AOI21_X1 _2064_ (.A(_0774_),
    .B1(_0765_),
    .B2(_0615_),
    .ZN(_0775_));
 NOR2_X1 _2065_ (.A1(_0014_),
    .A2(_0773_),
    .ZN(_0776_));
 NOR3_X1 _2066_ (.A1(_0771_),
    .A2(_0775_),
    .A3(_0776_),
    .ZN(_0286_));
 OR3_X1 _2067_ (.A1(\timer[5] ),
    .A2(\timer[4] ),
    .A3(_0690_),
    .ZN(_0777_));
 NOR2_X1 _2068_ (.A1(\timer[6] ),
    .A2(_0777_),
    .ZN(_0778_));
 XOR2_X1 _2069_ (.A(_0015_),
    .B(_0778_),
    .Z(_0779_));
 NOR3_X1 _2070_ (.A1(_0806_),
    .A2(_0831_),
    .A3(_0615_),
    .ZN(_0780_));
 NAND2_X1 _2071_ (.A1(_0015_),
    .A2(_0615_),
    .ZN(_0781_));
 AOI21_X1 _2072_ (.A(_0780_),
    .B1(_0781_),
    .B2(_0770_),
    .ZN(_0782_));
 OR2_X1 _2073_ (.A1(\init_state[4] ),
    .A2(_0823_),
    .ZN(_0783_));
 OAI21_X1 _2074_ (.A(_0762_),
    .B1(_0820_),
    .B2(_0015_),
    .ZN(_0784_));
 AOI22_X1 _2075_ (.A1(_0923_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0915_),
    .ZN(_0785_));
 AOI221_X1 _2076_ (.A(_0833_),
    .B1(_1170_),
    .B2(_0779_),
    .C1(_0782_),
    .C2(_0785_),
    .ZN(_0287_));
 NOR2_X1 _2077_ (.A1(\timer[7] ),
    .A2(\timer[6] ),
    .ZN(_0786_));
 NAND2_X1 _2078_ (.A1(_0786_),
    .A2(_0772_),
    .ZN(_0787_));
 XOR2_X1 _2079_ (.A(_0016_),
    .B(_0787_),
    .Z(_0788_));
 OAI21_X1 _2080_ (.A(_0788_),
    .B1(_0748_),
    .B2(_0678_),
    .ZN(_0789_));
 OAI22_X1 _2081_ (.A1(_0016_),
    .A2(_0695_),
    .B1(_0789_),
    .B2(_0615_),
    .ZN(_0790_));
 AND2_X1 _2082_ (.A1(_0478_),
    .A2(_0790_),
    .ZN(_0288_));
 OAI21_X1 _2083_ (.A(_0802_),
    .B1(_0448_),
    .B2(_0682_),
    .ZN(_0791_));
 NOR2_X1 _2084_ (.A1(_0813_),
    .A2(_0777_),
    .ZN(_0792_));
 NAND2_X1 _2085_ (.A1(_1170_),
    .A2(_0792_),
    .ZN(_0793_));
 NOR2_X1 _2086_ (.A1(_0615_),
    .A2(_0792_),
    .ZN(_0794_));
 NOR2_X1 _2087_ (.A1(_0017_),
    .A2(_0794_),
    .ZN(_0795_));
 AOI221_X1 _2088_ (.A(_0791_),
    .B1(_0793_),
    .B2(_0017_),
    .C1(_0795_),
    .C2(_0695_),
    .ZN(_0289_));
 NAND3_X1 _2089_ (.A1(_0888_),
    .A2(_0448_),
    .A3(net30),
    .ZN(_0796_));
 OR4_X1 _2090_ (.A1(_0888_),
    .A2(_0890_),
    .A3(_0661_),
    .A4(_0914_),
    .ZN(_0797_));
 AOI21_X1 _2091_ (.A(_1170_),
    .B1(_0796_),
    .B2(_0797_),
    .ZN(_0798_));
 AOI21_X1 _2092_ (.A(_0798_),
    .B1(_0675_),
    .B2(_0589_),
    .ZN(_0799_));
 NOR3_X1 _2093_ (.A1(_0835_),
    .A2(_0923_),
    .A3(_0799_),
    .ZN(_0290_));
 NOR2_X1 _2094_ (.A1(_1170_),
    .A2(_0603_),
    .ZN(net99));
 NOR2_X1 _2095_ (.A1(_0823_),
    .A2(_0836_),
    .ZN(_0800_));
 AOI21_X1 _2096_ (.A(_0834_),
    .B1(_0655_),
    .B2(_0800_),
    .ZN(net129));
 HA_X1 _2097_ (.A(_1145_),
    .B(_1146_),
    .CO(_1147_),
    .S(_1148_));
 HA_X1 _2098_ (.A(_1145_),
    .B(net116),
    .CO(_1149_),
    .S(_1150_));
 HA_X1 _2099_ (.A(net115),
    .B(_1146_),
    .CO(_1151_),
    .S(_1152_));
 HA_X1 _2100_ (.A(net115),
    .B(net116),
    .CO(_1153_),
    .S(_1154_));
 HA_X1 _2101_ (.A(_1155_),
    .B(_1156_),
    .CO(_1157_),
    .S(_1158_));
 HA_X1 _2102_ (.A(_1155_),
    .B(_1156_),
    .CO(_1159_),
    .S(_1160_));
 HA_X1 _2103_ (.A(_1161_),
    .B(_1162_),
    .CO(_1163_),
    .S(_1164_));
 HA_X1 _2104_ (.A(_1161_),
    .B(\refresh_counter[1] ),
    .CO(_1165_),
    .S(_1166_));
 HA_X1 _2105_ (.A(\refresh_counter[0] ),
    .B(\refresh_counter[1] ),
    .CO(_1167_),
    .S(_1168_));
 HA_X1 _2106_ (.A(_1169_),
    .B(_1170_),
    .CO(_1171_),
    .S(_1172_));
 HA_X1 _2107_ (.A(\timer[0] ),
    .B(_1170_),
    .CO(_1173_),
    .S(_1174_));
 HA_X1 _2108_ (.A(_1169_),
    .B(_1175_),
    .CO(_1176_),
    .S(_1177_));
 HA_X1 _2109_ (.A(\timer[0] ),
    .B(_1175_),
    .CO(_1178_),
    .S(_1179_));
 HA_X1 _2110_ (.A(_1180_),
    .B(_1181_),
    .CO(_1182_),
    .S(_1183_));
 HA_X1 _2111_ (.A(_1180_),
    .B(net197),
    .CO(_1184_),
    .S(_1185_));
 HA_X1 _2112_ (.A(net196),
    .B(_1181_),
    .CO(_1186_),
    .S(_1187_));
 HA_X1 _2113_ (.A(net196),
    .B(net197),
    .CO(_1188_),
    .S(_1189_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 LOGIC1_X1 _2118__209 (.Z(net209));
 BUF_X1 _2116_ (.A(net199),
    .Z(phy_bank_group[0]));
 BUF_X1 _2117_ (.A(net200),
    .Z(phy_bank_group[1]));
 BUF_X1 _2118_ (.A(net209),
    .Z(phy_cke));
 BUF_X1 _2119_ (.A(wr_mask[0]),
    .Z(net120));
 BUF_X1 _2120_ (.A(wr_mask[1]),
    .Z(net121));
 BUF_X1 _2121_ (.A(wr_mask[2]),
    .Z(net122));
 BUF_X1 _2122_ (.A(wr_mask[3]),
    .Z(net123));
 BUF_X1 _2123_ (.A(wr_mask[4]),
    .Z(net124));
 BUF_X1 _2124_ (.A(wr_mask[5]),
    .Z(net125));
 BUF_X1 _2125_ (.A(wr_mask[6]),
    .Z(net126));
 BUF_X1 _2126_ (.A(wr_mask[7]),
    .Z(net127));
 BUF_X1 _2127_ (.A(net34),
    .Z(phy_dq[0]));
 BUF_X1 _2128_ (.A(net45),
    .Z(phy_dq[1]));
 BUF_X1 _2129_ (.A(net56),
    .Z(phy_dq[2]));
 BUF_X1 _2130_ (.A(net67),
    .Z(phy_dq[3]));
 BUF_X1 _2131_ (.A(net78),
    .Z(phy_dq[4]));
 BUF_X1 _2132_ (.A(net89),
    .Z(phy_dq[5]));
 BUF_X1 _2133_ (.A(net94),
    .Z(phy_dq[6]));
 BUF_X1 _2134_ (.A(net95),
    .Z(phy_dq[7]));
 BUF_X1 _2135_ (.A(net96),
    .Z(phy_dq[8]));
 BUF_X1 _2136_ (.A(net97),
    .Z(phy_dq[9]));
 BUF_X1 _2137_ (.A(net35),
    .Z(phy_dq[10]));
 BUF_X1 _2138_ (.A(net36),
    .Z(phy_dq[11]));
 BUF_X1 _2139_ (.A(net37),
    .Z(phy_dq[12]));
 BUF_X1 _2140_ (.A(net38),
    .Z(phy_dq[13]));
 BUF_X1 _2141_ (.A(net39),
    .Z(phy_dq[14]));
 BUF_X1 _2142_ (.A(net40),
    .Z(phy_dq[15]));
 BUF_X1 _2143_ (.A(net41),
    .Z(phy_dq[16]));
 BUF_X1 _2144_ (.A(net42),
    .Z(phy_dq[17]));
 BUF_X1 _2145_ (.A(net43),
    .Z(phy_dq[18]));
 BUF_X1 _2146_ (.A(net44),
    .Z(phy_dq[19]));
 BUF_X1 _2147_ (.A(net46),
    .Z(phy_dq[20]));
 BUF_X1 _2148_ (.A(net47),
    .Z(phy_dq[21]));
 BUF_X1 _2149_ (.A(net48),
    .Z(phy_dq[22]));
 BUF_X1 _2150_ (.A(net49),
    .Z(phy_dq[23]));
 BUF_X1 _2151_ (.A(net50),
    .Z(phy_dq[24]));
 BUF_X1 _2152_ (.A(net51),
    .Z(phy_dq[25]));
 BUF_X1 _2153_ (.A(net52),
    .Z(phy_dq[26]));
 BUF_X1 _2154_ (.A(net53),
    .Z(phy_dq[27]));
 BUF_X1 _2155_ (.A(net54),
    .Z(phy_dq[28]));
 BUF_X1 _2156_ (.A(net55),
    .Z(phy_dq[29]));
 BUF_X1 _2157_ (.A(net57),
    .Z(phy_dq[30]));
 BUF_X1 _2158_ (.A(net58),
    .Z(phy_dq[31]));
 BUF_X1 _2159_ (.A(net59),
    .Z(phy_dq[32]));
 BUF_X1 _2160_ (.A(net60),
    .Z(phy_dq[33]));
 BUF_X1 _2161_ (.A(net61),
    .Z(phy_dq[34]));
 BUF_X1 _2162_ (.A(net62),
    .Z(phy_dq[35]));
 BUF_X1 _2163_ (.A(net63),
    .Z(phy_dq[36]));
 BUF_X1 _2164_ (.A(net64),
    .Z(phy_dq[37]));
 BUF_X1 _2165_ (.A(net65),
    .Z(phy_dq[38]));
 BUF_X1 _2166_ (.A(net66),
    .Z(phy_dq[39]));
 BUF_X1 _2167_ (.A(net68),
    .Z(phy_dq[40]));
 BUF_X1 _2168_ (.A(net69),
    .Z(phy_dq[41]));
 BUF_X1 _2169_ (.A(net70),
    .Z(phy_dq[42]));
 BUF_X1 _2170_ (.A(net71),
    .Z(phy_dq[43]));
 BUF_X1 _2171_ (.A(net72),
    .Z(phy_dq[44]));
 BUF_X1 _2172_ (.A(net73),
    .Z(phy_dq[45]));
 BUF_X1 _2173_ (.A(net74),
    .Z(phy_dq[46]));
 BUF_X1 _2174_ (.A(net75),
    .Z(phy_dq[47]));
 BUF_X1 _2175_ (.A(net76),
    .Z(phy_dq[48]));
 BUF_X1 _2176_ (.A(net77),
    .Z(phy_dq[49]));
 BUF_X1 _2177_ (.A(net79),
    .Z(phy_dq[50]));
 BUF_X1 _2178_ (.A(net80),
    .Z(phy_dq[51]));
 BUF_X1 _2179_ (.A(net81),
    .Z(phy_dq[52]));
 BUF_X1 _2180_ (.A(net82),
    .Z(phy_dq[53]));
 BUF_X1 _2181_ (.A(net83),
    .Z(phy_dq[54]));
 BUF_X1 _2182_ (.A(net84),
    .Z(phy_dq[55]));
 BUF_X1 _2183_ (.A(net85),
    .Z(phy_dq[56]));
 BUF_X1 _2184_ (.A(net86),
    .Z(phy_dq[57]));
 BUF_X1 _2185_ (.A(net87),
    .Z(phy_dq[58]));
 BUF_X1 _2186_ (.A(net88),
    .Z(phy_dq[59]));
 BUF_X1 _2187_ (.A(net90),
    .Z(phy_dq[60]));
 BUF_X1 _2188_ (.A(net91),
    .Z(phy_dq[61]));
 BUF_X1 _2189_ (.A(net92),
    .Z(phy_dq[62]));
 BUF_X1 _2190_ (.A(net93),
    .Z(phy_dq[63]));
 BUF_X1 _2191_ (.A(net201),
    .Z(phy_dqs_n[0]));
 BUF_X1 _2192_ (.A(net202),
    .Z(phy_dqs_n[1]));
 BUF_X1 _2193_ (.A(net203),
    .Z(phy_dqs_n[2]));
 BUF_X1 _2194_ (.A(net204),
    .Z(phy_dqs_n[3]));
 BUF_X1 _2195_ (.A(net205),
    .Z(phy_dqs_n[4]));
 BUF_X1 _2196_ (.A(net206),
    .Z(phy_dqs_n[5]));
 BUF_X1 _2197_ (.A(net207),
    .Z(phy_dqs_n[6]));
 BUF_X1 _2198_ (.A(net208),
    .Z(phy_dqs_n[7]));
 BUF_X1 _2199_ (.A(net210),
    .Z(phy_dqs_p[0]));
 BUF_X1 _2200_ (.A(net211),
    .Z(phy_dqs_p[1]));
 BUF_X1 _2201_ (.A(net212),
    .Z(phy_dqs_p[2]));
 BUF_X1 _2202_ (.A(net213),
    .Z(phy_dqs_p[3]));
 BUF_X1 _2203_ (.A(net214),
    .Z(phy_dqs_p[4]));
 BUF_X1 _2204_ (.A(net215),
    .Z(phy_dqs_p[5]));
 BUF_X1 _2205_ (.A(net216),
    .Z(phy_dqs_p[6]));
 BUF_X1 _2206_ (.A(net217),
    .Z(phy_dqs_p[7]));
 BUF_X1 _2207_ (.A(net218),
    .Z(phy_odt));
 DFF_X1 \active_row[0][0]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[0][0] ),
    .QN(_1135_));
 DFF_X1 \active_row[0][10]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[0][10] ),
    .QN(_1134_));
 DFF_X1 \active_row[0][11]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[0][11] ),
    .QN(_1133_));
 DFF_X1 \active_row[0][12]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[0][12] ),
    .QN(_1132_));
 DFF_X1 \active_row[0][13]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[0][13] ),
    .QN(_1131_));
 DFF_X1 \active_row[0][1]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[0][1] ),
    .QN(_1130_));
 DFF_X1 \active_row[0][2]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[0][2] ),
    .QN(_1129_));
 DFF_X1 \active_row[0][3]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[0][3] ),
    .QN(_1128_));
 DFF_X1 \active_row[0][4]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[0][4] ),
    .QN(_1127_));
 DFF_X1 \active_row[0][5]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[0][5] ),
    .QN(_1126_));
 DFF_X1 \active_row[0][6]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_4_3_0_clk),
    .Q(\active_row[0][6] ),
    .QN(_1125_));
 DFF_X1 \active_row[0][7]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[0][7] ),
    .QN(_1124_));
 DFF_X1 \active_row[0][8]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[0][8] ),
    .QN(_1123_));
 DFF_X1 \active_row[0][9]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[0][9] ),
    .QN(_1122_));
 DFF_X1 \active_row[1][0]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[1][0] ),
    .QN(_1121_));
 DFF_X1 \active_row[1][10]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[1][10] ),
    .QN(_1120_));
 DFF_X1 \active_row[1][11]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[1][11] ),
    .QN(_1119_));
 DFF_X1 \active_row[1][12]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[1][12] ),
    .QN(_1118_));
 DFF_X1 \active_row[1][13]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[1][13] ),
    .QN(_1117_));
 DFF_X1 \active_row[1][1]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[1][1] ),
    .QN(_1116_));
 DFF_X1 \active_row[1][2]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[1][2] ),
    .QN(_1115_));
 DFF_X1 \active_row[1][3]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[1][3] ),
    .QN(_1114_));
 DFF_X1 \active_row[1][4]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[1][4] ),
    .QN(_1113_));
 DFF_X1 \active_row[1][5]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[1][5] ),
    .QN(_1112_));
 DFF_X1 \active_row[1][6]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_4_3_0_clk),
    .Q(\active_row[1][6] ),
    .QN(_1111_));
 DFF_X1 \active_row[1][7]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[1][7] ),
    .QN(_1110_));
 DFF_X1 \active_row[1][8]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[1][8] ),
    .QN(_1109_));
 DFF_X1 \active_row[1][9]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[1][9] ),
    .QN(_1108_));
 DFF_X1 \active_row[2][0]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[2][0] ),
    .QN(_1107_));
 DFF_X1 \active_row[2][10]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[2][10] ),
    .QN(_1106_));
 DFF_X1 \active_row[2][11]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[2][11] ),
    .QN(_1105_));
 DFF_X1 \active_row[2][12]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[2][12] ),
    .QN(_1104_));
 DFF_X1 \active_row[2][13]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[2][13] ),
    .QN(_1103_));
 DFF_X1 \active_row[2][1]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[2][1] ),
    .QN(_1102_));
 DFF_X1 \active_row[2][2]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[2][2] ),
    .QN(_1101_));
 DFF_X1 \active_row[2][3]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[2][3] ),
    .QN(_1100_));
 DFF_X1 \active_row[2][4]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[2][4] ),
    .QN(_1099_));
 DFF_X1 \active_row[2][5]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[2][5] ),
    .QN(_1098_));
 DFF_X1 \active_row[2][6]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_4_3_0_clk),
    .Q(\active_row[2][6] ),
    .QN(_1097_));
 DFF_X1 \active_row[2][7]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[2][7] ),
    .QN(_1096_));
 DFF_X1 \active_row[2][8]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[2][8] ),
    .QN(_1095_));
 DFF_X1 \active_row[2][9]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[2][9] ),
    .QN(_1094_));
 DFF_X1 \active_row[3][0]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[3][0] ),
    .QN(_1093_));
 DFF_X1 \active_row[3][10]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[3][10] ),
    .QN(_1092_));
 DFF_X1 \active_row[3][11]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[3][11] ),
    .QN(_1091_));
 DFF_X1 \active_row[3][12]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[3][12] ),
    .QN(_1090_));
 DFF_X1 \active_row[3][13]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[3][13] ),
    .QN(_1089_));
 DFF_X1 \active_row[3][1]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[3][1] ),
    .QN(_1088_));
 DFF_X1 \active_row[3][2]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[3][2] ),
    .QN(_1087_));
 DFF_X1 \active_row[3][3]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[3][3] ),
    .QN(_1086_));
 DFF_X1 \active_row[3][4]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[3][4] ),
    .QN(_1085_));
 DFF_X1 \active_row[3][5]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[3][5] ),
    .QN(_1084_));
 DFF_X1 \active_row[3][6]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[3][6] ),
    .QN(_1083_));
 DFF_X1 \active_row[3][7]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[3][7] ),
    .QN(_1082_));
 DFF_X1 \active_row[3][8]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[3][8] ),
    .QN(_1081_));
 DFF_X1 \active_row[3][9]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[3][9] ),
    .QN(_1080_));
 DFF_X1 \active_row[4][0]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[4][0] ),
    .QN(_1079_));
 DFF_X1 \active_row[4][10]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[4][10] ),
    .QN(_1078_));
 DFF_X1 \active_row[4][11]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[4][11] ),
    .QN(_1077_));
 DFF_X1 \active_row[4][12]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[4][12] ),
    .QN(_1076_));
 DFF_X1 \active_row[4][13]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[4][13] ),
    .QN(_1075_));
 DFF_X1 \active_row[4][1]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[4][1] ),
    .QN(_1074_));
 DFF_X1 \active_row[4][2]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[4][2] ),
    .QN(_1073_));
 DFF_X1 \active_row[4][3]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[4][3] ),
    .QN(_1072_));
 DFF_X1 \active_row[4][4]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[4][4] ),
    .QN(_1071_));
 DFF_X1 \active_row[4][5]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[4][5] ),
    .QN(_1070_));
 DFF_X1 \active_row[4][6]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_4_3_0_clk),
    .Q(\active_row[4][6] ),
    .QN(_1069_));
 DFF_X1 \active_row[4][7]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[4][7] ),
    .QN(_1068_));
 DFF_X1 \active_row[4][8]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[4][8] ),
    .QN(_1067_));
 DFF_X1 \active_row[4][9]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[4][9] ),
    .QN(_1066_));
 DFF_X1 \active_row[5][0]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[5][0] ),
    .QN(_1065_));
 DFF_X1 \active_row[5][10]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[5][10] ),
    .QN(_1064_));
 DFF_X1 \active_row[5][11]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[5][11] ),
    .QN(_1063_));
 DFF_X1 \active_row[5][12]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[5][12] ),
    .QN(_1062_));
 DFF_X1 \active_row[5][13]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[5][13] ),
    .QN(_1061_));
 DFF_X1 \active_row[5][1]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[5][1] ),
    .QN(_1060_));
 DFF_X1 \active_row[5][2]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[5][2] ),
    .QN(_1059_));
 DFF_X1 \active_row[5][3]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_4_12_0_clk),
    .Q(\active_row[5][3] ),
    .QN(_1058_));
 DFF_X1 \active_row[5][4]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[5][4] ),
    .QN(_1057_));
 DFF_X1 \active_row[5][5]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[5][5] ),
    .QN(_1056_));
 DFF_X1 \active_row[5][6]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[5][6] ),
    .QN(_1055_));
 DFF_X1 \active_row[5][7]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[5][7] ),
    .QN(_1054_));
 DFF_X1 \active_row[5][8]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[5][8] ),
    .QN(_1053_));
 DFF_X1 \active_row[5][9]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[5][9] ),
    .QN(_1052_));
 DFF_X1 \active_row[6][0]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[6][0] ),
    .QN(_1051_));
 DFF_X1 \active_row[6][10]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[6][10] ),
    .QN(_1050_));
 DFF_X1 \active_row[6][11]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[6][11] ),
    .QN(_1049_));
 DFF_X1 \active_row[6][12]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[6][12] ),
    .QN(_1048_));
 DFF_X1 \active_row[6][13]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[6][13] ),
    .QN(_1047_));
 DFF_X1 \active_row[6][1]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[6][1] ),
    .QN(_1046_));
 DFF_X1 \active_row[6][2]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[6][2] ),
    .QN(_1045_));
 DFF_X1 \active_row[6][3]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[6][3] ),
    .QN(_1044_));
 DFF_X1 \active_row[6][4]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[6][4] ),
    .QN(_1043_));
 DFF_X1 \active_row[6][5]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[6][5] ),
    .QN(_1042_));
 DFF_X1 \active_row[6][6]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[6][6] ),
    .QN(_1041_));
 DFF_X1 \active_row[6][7]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[6][7] ),
    .QN(_1040_));
 DFF_X1 \active_row[6][8]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[6][8] ),
    .QN(_1039_));
 DFF_X1 \active_row[6][9]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[6][9] ),
    .QN(_1038_));
 DFF_X1 \active_row[7][0]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[7][0] ),
    .QN(_1037_));
 DFF_X1 \active_row[7][10]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_4_11_0_clk),
    .Q(\active_row[7][10] ),
    .QN(_1036_));
 DFF_X1 \active_row[7][11]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[7][11] ),
    .QN(_1035_));
 DFF_X1 \active_row[7][12]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[7][12] ),
    .QN(_1034_));
 DFF_X1 \active_row[7][13]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_4_15_0_clk),
    .Q(\active_row[7][13] ),
    .QN(_1033_));
 DFF_X1 \active_row[7][1]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_4_14_0_clk),
    .Q(\active_row[7][1] ),
    .QN(_1032_));
 DFF_X1 \active_row[7][2]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[7][2] ),
    .QN(_1031_));
 DFF_X1 \active_row[7][3]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[7][3] ),
    .QN(_1030_));
 DFF_X1 \active_row[7][4]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_4_10_0_clk),
    .Q(\active_row[7][4] ),
    .QN(_1029_));
 DFF_X1 \active_row[7][5]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_4_13_0_clk),
    .Q(\active_row[7][5] ),
    .QN(_1028_));
 DFF_X1 \active_row[7][6]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[7][6] ),
    .QN(_1027_));
 DFF_X1 \active_row[7][7]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_4_9_0_clk),
    .Q(\active_row[7][7] ),
    .QN(_1026_));
 DFF_X1 \active_row[7][8]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_4_8_0_clk),
    .Q(\active_row[7][8] ),
    .QN(_1025_));
 DFF_X1 \active_row[7][9]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_4_2_0_clk),
    .Q(\active_row[7][9] ),
    .QN(_1024_));
 DFF_X1 \addr_reg[0]$_SDFFE_PN0P_  (.D(_0158_),
    .CK(clknet_4_14_0_clk),
    .Q(net101),
    .QN(_1023_));
 DFF_X1 \addr_reg[10]$_SDFFE_PN0P_  (.D(_0159_),
    .CK(clknet_4_14_0_clk),
    .Q(net102),
    .QN(_1022_));
 DFF_X1 \addr_reg[11]$_SDFFE_PN0P_  (.D(_0160_),
    .CK(clknet_4_9_0_clk),
    .Q(net103),
    .QN(_1021_));
 DFF_X1 \addr_reg[12]$_SDFFE_PN0P_  (.D(_0161_),
    .CK(clknet_4_14_0_clk),
    .Q(net104),
    .QN(_1020_));
 DFF_X1 \addr_reg[13]$_SDFFE_PN0P_  (.D(_0162_),
    .CK(clknet_4_14_0_clk),
    .Q(net105),
    .QN(_1019_));
 DFF_X1 \addr_reg[1]$_SDFFE_PN0P_  (.D(_0163_),
    .CK(clknet_4_14_0_clk),
    .Q(net106),
    .QN(_1018_));
 DFF_X1 \addr_reg[2]$_SDFFE_PN0P_  (.D(_0164_),
    .CK(clknet_4_14_0_clk),
    .Q(net107),
    .QN(_1017_));
 DFF_X1 \addr_reg[3]$_SDFFE_PN0P_  (.D(_0165_),
    .CK(clknet_4_13_0_clk),
    .Q(net108),
    .QN(_1016_));
 DFF_X1 \addr_reg[4]$_SDFFE_PN0P_  (.D(_0166_),
    .CK(clknet_4_8_0_clk),
    .Q(net109),
    .QN(_1015_));
 DFF_X1 \addr_reg[5]$_SDFFE_PN0P_  (.D(_0167_),
    .CK(clknet_4_13_0_clk),
    .Q(net110),
    .QN(_1014_));
 DFF_X1 \addr_reg[6]$_SDFFE_PN0P_  (.D(_0168_),
    .CK(clknet_4_8_0_clk),
    .Q(net111),
    .QN(_1013_));
 DFF_X1 \addr_reg[7]$_SDFFE_PN0P_  (.D(_0169_),
    .CK(clknet_4_12_0_clk),
    .Q(net112),
    .QN(_1012_));
 DFF_X1 \addr_reg[8]$_SDFFE_PN0P_  (.D(_0170_),
    .CK(clknet_4_2_0_clk),
    .Q(net113),
    .QN(_1011_));
 DFF_X1 \addr_reg[9]$_SDFFE_PN0P_  (.D(_0171_),
    .CK(clknet_4_8_0_clk),
    .Q(net114),
    .QN(_1010_));
 DFF_X1 \bank_active[0]$_SDFFE_PN0P_  (.D(_0172_),
    .CK(clknet_4_6_0_clk),
    .Q(\bank_active[0] ),
    .QN(_0024_));
 DFF_X1 \bank_active[1]$_SDFFE_PN0P_  (.D(_0173_),
    .CK(clknet_4_7_0_clk),
    .Q(\bank_active[1] ),
    .QN(_0025_));
 DFF_X1 \bank_active[2]$_SDFFE_PN0P_  (.D(_0174_),
    .CK(clknet_4_6_0_clk),
    .Q(\bank_active[2] ),
    .QN(_0026_));
 DFF_X1 \bank_active[3]$_SDFFE_PN0P_  (.D(_0175_),
    .CK(clknet_4_13_0_clk),
    .Q(\bank_active[3] ),
    .QN(_0027_));
 DFF_X1 \bank_active[4]$_SDFFE_PN0P_  (.D(_0176_),
    .CK(clknet_4_6_0_clk),
    .Q(\bank_active[4] ),
    .QN(_0028_));
 DFF_X1 \bank_active[5]$_SDFFE_PN0P_  (.D(_0177_),
    .CK(clknet_4_7_0_clk),
    .Q(\bank_active[5] ),
    .QN(_0029_));
 DFF_X1 \bank_active[6]$_SDFFE_PN0P_  (.D(_0178_),
    .CK(clknet_4_6_0_clk),
    .Q(\bank_active[6] ),
    .QN(_0030_));
 DFF_X1 \bank_active[7]$_SDFFE_PN0P_  (.D(_0179_),
    .CK(clknet_4_7_0_clk),
    .Q(\bank_active[7] ),
    .QN(_0031_));
 DFF_X2 \bank_reg[0]$_SDFFE_PN0P_  (.D(_0180_),
    .CK(clknet_4_3_0_clk),
    .Q(net115),
    .QN(_1145_));
 DFF_X2 \bank_reg[1]$_SDFFE_PN0P_  (.D(_0181_),
    .CK(clknet_4_6_0_clk),
    .Q(net116),
    .QN(_1146_));
 DFF_X1 \bank_reg[2]$_SDFFE_PN0P_  (.D(_0182_),
    .CK(clknet_4_3_0_clk),
    .Q(net117),
    .QN(_1009_));
 DFF_X1 \burst_counter[0]$_SDFFE_PN0P_  (.D(_0183_),
    .CK(clknet_4_7_0_clk),
    .Q(\burst_counter[0] ),
    .QN(_1155_));
 DFF_X1 \burst_counter[1]$_SDFFE_PN0P_  (.D(_0184_),
    .CK(clknet_4_7_0_clk),
    .Q(\burst_counter[1] ),
    .QN(_1156_));
 DFF_X1 \burst_counter[2]$_SDFFE_PN0P_  (.D(_0185_),
    .CK(clknet_4_7_0_clk),
    .Q(\burst_counter[2] ),
    .QN(_1008_));
 DFF_X1 \burst_counter[3]$_SDFFE_PN0P_  (.D(_0186_),
    .CK(clknet_4_7_0_clk),
    .Q(\burst_counter[3] ),
    .QN(_1007_));
 DFF_X1 \cmd_reg[0]$_SDFF_PN1_  (.D(_0187_),
    .CK(clknet_4_4_0_clk),
    .Q(net130),
    .QN(_1006_));
 DFF_X1 \cmd_reg[1]$_SDFF_PN1_  (.D(_0188_),
    .CK(clknet_4_5_0_clk),
    .Q(net118),
    .QN(_1005_));
 DFF_X2 \cmd_reg[2]$_SDFF_PN1_  (.D(_0189_),
    .CK(clknet_4_5_0_clk),
    .Q(net128),
    .QN(_1136_));
 DFF_X1 \cmd_reg_valid$_DFF_P_  (.D(net33),
    .CK(clknet_4_1_0_clk),
    .Q(cmd_reg_valid),
    .QN(net119));
 DFF_X2 \curr_state[0]$_SDFFE_PN0P_  (.D(_0190_),
    .CK(clknet_4_1_0_clk),
    .Q(net196),
    .QN(_1180_));
 DFF_X2 \curr_state[1]$_SDFFE_PN0P_  (.D(_0191_),
    .CK(clknet_4_1_0_clk),
    .Q(net197),
    .QN(_1181_));
 DFF_X1 \init_done_reg$_SDFFE_PN0P_  (.D(_0192_),
    .CK(clknet_4_1_0_clk),
    .Q(net100),
    .QN(_1137_));
 DFF_X1 \init_state[0]$_DFF_P_  (.D(_0000_),
    .CK(clknet_4_1_0_clk),
    .Q(\init_state[0] ),
    .QN(_1138_));
 DFF_X1 \init_state[1]$_DFF_P_  (.D(_0001_),
    .CK(clknet_4_3_0_clk),
    .Q(\init_state[1] ),
    .QN(_1139_));
 DFF_X2 \init_state[2]$_DFF_P_  (.D(_0002_),
    .CK(clknet_4_3_0_clk),
    .Q(\init_state[2] ),
    .QN(_1140_));
 DFF_X1 \init_state[3]$_DFF_P_  (.D(_0003_),
    .CK(clknet_4_1_0_clk),
    .Q(\init_state[3] ),
    .QN(_1141_));
 DFF_X1 \init_state[4]$_DFF_P_  (.D(_0004_),
    .CK(clknet_4_1_0_clk),
    .Q(\init_state[4] ),
    .QN(_1142_));
 DFF_X1 \init_state[5]$_DFF_P_  (.D(_0005_),
    .CK(clknet_4_3_0_clk),
    .Q(\init_state[5] ),
    .QN(_1143_));
 DFF_X2 \init_state[6]$_DFF_P_  (.D(_0006_),
    .CK(clknet_4_3_0_clk),
    .Q(\init_state[6] ),
    .QN(_1144_));
 DFF_X1 \init_state[7]$_DFF_P_  (.D(_0007_),
    .CK(clknet_4_1_0_clk),
    .Q(\init_state[7] ),
    .QN(_0032_));
 DFF_X1 \rd_data_reg[0]$_DFFE_PP_  (.D(_0193_),
    .CK(net31),
    .Q(net131),
    .QN(_1004_));
 DFF_X1 \rd_data_reg[10]$_DFFE_PP_  (.D(_0194_),
    .CK(net31),
    .Q(net132),
    .QN(_1003_));
 DFF_X1 \rd_data_reg[11]$_DFFE_PP_  (.D(_0195_),
    .CK(net31),
    .Q(net133),
    .QN(_1002_));
 DFF_X1 \rd_data_reg[12]$_DFFE_PP_  (.D(_0196_),
    .CK(net31),
    .Q(net134),
    .QN(_1001_));
 DFF_X1 \rd_data_reg[13]$_DFFE_PP_  (.D(_0197_),
    .CK(net31),
    .Q(net135),
    .QN(_1000_));
 DFF_X1 \rd_data_reg[14]$_DFFE_PP_  (.D(_0198_),
    .CK(net31),
    .Q(net136),
    .QN(_0999_));
 DFF_X1 \rd_data_reg[15]$_DFFE_PP_  (.D(_0199_),
    .CK(net31),
    .Q(net137),
    .QN(_0998_));
 DFF_X1 \rd_data_reg[16]$_DFFE_PP_  (.D(_0200_),
    .CK(net31),
    .Q(net138),
    .QN(_0997_));
 DFF_X1 \rd_data_reg[17]$_DFFE_PP_  (.D(_0201_),
    .CK(net31),
    .Q(net139),
    .QN(_0996_));
 DFF_X1 \rd_data_reg[18]$_DFFE_PP_  (.D(_0202_),
    .CK(net31),
    .Q(net140),
    .QN(_0995_));
 DFF_X1 \rd_data_reg[19]$_DFFE_PP_  (.D(_0203_),
    .CK(net31),
    .Q(net141),
    .QN(_0994_));
 DFF_X1 \rd_data_reg[1]$_DFFE_PP_  (.D(_0204_),
    .CK(net31),
    .Q(net142),
    .QN(_0993_));
 DFF_X1 \rd_data_reg[20]$_DFFE_PP_  (.D(_0205_),
    .CK(net31),
    .Q(net143),
    .QN(_0992_));
 DFF_X1 \rd_data_reg[21]$_DFFE_PP_  (.D(_0206_),
    .CK(net31),
    .Q(net144),
    .QN(_0991_));
 DFF_X1 \rd_data_reg[22]$_DFFE_PP_  (.D(_0207_),
    .CK(net31),
    .Q(net145),
    .QN(_0990_));
 DFF_X1 \rd_data_reg[23]$_DFFE_PP_  (.D(_0208_),
    .CK(net31),
    .Q(net146),
    .QN(_0989_));
 DFF_X1 \rd_data_reg[24]$_DFFE_PP_  (.D(_0209_),
    .CK(net31),
    .Q(net147),
    .QN(_0988_));
 DFF_X1 \rd_data_reg[25]$_DFFE_PP_  (.D(_0210_),
    .CK(net31),
    .Q(net148),
    .QN(_0987_));
 DFF_X1 \rd_data_reg[26]$_DFFE_PP_  (.D(_0211_),
    .CK(net31),
    .Q(net149),
    .QN(_0986_));
 DFF_X1 \rd_data_reg[27]$_DFFE_PP_  (.D(_0212_),
    .CK(net31),
    .Q(net150),
    .QN(_0985_));
 DFF_X1 \rd_data_reg[28]$_DFFE_PP_  (.D(_0213_),
    .CK(net31),
    .Q(net151),
    .QN(_0984_));
 DFF_X1 \rd_data_reg[29]$_DFFE_PP_  (.D(_0214_),
    .CK(net31),
    .Q(net152),
    .QN(_0983_));
 DFF_X1 \rd_data_reg[2]$_DFFE_PP_  (.D(_0215_),
    .CK(net31),
    .Q(net153),
    .QN(_0982_));
 DFF_X1 \rd_data_reg[30]$_DFFE_PP_  (.D(_0216_),
    .CK(net31),
    .Q(net154),
    .QN(_0981_));
 DFF_X1 \rd_data_reg[31]$_DFFE_PP_  (.D(_0217_),
    .CK(net31),
    .Q(net155),
    .QN(_0980_));
 DFF_X1 \rd_data_reg[32]$_DFFE_PP_  (.D(_0218_),
    .CK(net31),
    .Q(net156),
    .QN(_0979_));
 DFF_X1 \rd_data_reg[33]$_DFFE_PP_  (.D(_0219_),
    .CK(net31),
    .Q(net157),
    .QN(_0978_));
 DFF_X1 \rd_data_reg[34]$_DFFE_PP_  (.D(_0220_),
    .CK(net31),
    .Q(net158),
    .QN(_0977_));
 DFF_X1 \rd_data_reg[35]$_DFFE_PP_  (.D(_0221_),
    .CK(net31),
    .Q(net159),
    .QN(_0976_));
 DFF_X1 \rd_data_reg[36]$_DFFE_PP_  (.D(_0222_),
    .CK(net31),
    .Q(net160),
    .QN(_0975_));
 DFF_X1 \rd_data_reg[37]$_DFFE_PP_  (.D(_0223_),
    .CK(net31),
    .Q(net161),
    .QN(_0974_));
 DFF_X1 \rd_data_reg[38]$_DFFE_PP_  (.D(_0224_),
    .CK(net31),
    .Q(net162),
    .QN(_0973_));
 DFF_X1 \rd_data_reg[39]$_DFFE_PP_  (.D(_0225_),
    .CK(net31),
    .Q(net163),
    .QN(_0972_));
 DFF_X1 \rd_data_reg[3]$_DFFE_PP_  (.D(_0226_),
    .CK(net31),
    .Q(net164),
    .QN(_0971_));
 DFF_X1 \rd_data_reg[40]$_DFFE_PP_  (.D(_0227_),
    .CK(net31),
    .Q(net165),
    .QN(_0970_));
 DFF_X1 \rd_data_reg[41]$_DFFE_PP_  (.D(_0228_),
    .CK(net31),
    .Q(net166),
    .QN(_0969_));
 DFF_X1 \rd_data_reg[42]$_DFFE_PP_  (.D(_0229_),
    .CK(net31),
    .Q(net167),
    .QN(_0968_));
 DFF_X1 \rd_data_reg[43]$_DFFE_PP_  (.D(_0230_),
    .CK(net31),
    .Q(net168),
    .QN(_0967_));
 DFF_X1 \rd_data_reg[44]$_DFFE_PP_  (.D(_0231_),
    .CK(net31),
    .Q(net169),
    .QN(_0966_));
 DFF_X1 \rd_data_reg[45]$_DFFE_PP_  (.D(_0232_),
    .CK(net31),
    .Q(net170),
    .QN(_0965_));
 DFF_X1 \rd_data_reg[46]$_DFFE_PP_  (.D(_0233_),
    .CK(net31),
    .Q(net171),
    .QN(_0964_));
 DFF_X1 \rd_data_reg[47]$_DFFE_PP_  (.D(_0234_),
    .CK(net31),
    .Q(net172),
    .QN(_0963_));
 DFF_X1 \rd_data_reg[48]$_DFFE_PP_  (.D(_0235_),
    .CK(net31),
    .Q(net173),
    .QN(_0962_));
 DFF_X1 \rd_data_reg[49]$_DFFE_PP_  (.D(_0236_),
    .CK(net31),
    .Q(net174),
    .QN(_0961_));
 DFF_X1 \rd_data_reg[4]$_DFFE_PP_  (.D(_0237_),
    .CK(net31),
    .Q(net175),
    .QN(_0960_));
 DFF_X1 \rd_data_reg[50]$_DFFE_PP_  (.D(_0238_),
    .CK(net31),
    .Q(net176),
    .QN(_0959_));
 DFF_X1 \rd_data_reg[51]$_DFFE_PP_  (.D(_0239_),
    .CK(net31),
    .Q(net177),
    .QN(_0958_));
 DFF_X1 \rd_data_reg[52]$_DFFE_PP_  (.D(_0240_),
    .CK(net31),
    .Q(net178),
    .QN(_0957_));
 DFF_X1 \rd_data_reg[53]$_DFFE_PP_  (.D(_0241_),
    .CK(net31),
    .Q(net179),
    .QN(_0956_));
 DFF_X1 \rd_data_reg[54]$_DFFE_PP_  (.D(_0242_),
    .CK(net31),
    .Q(net180),
    .QN(_0955_));
 DFF_X1 \rd_data_reg[55]$_DFFE_PP_  (.D(_0243_),
    .CK(net31),
    .Q(net181),
    .QN(_0954_));
 DFF_X1 \rd_data_reg[56]$_DFFE_PP_  (.D(_0244_),
    .CK(net31),
    .Q(net182),
    .QN(_0953_));
 DFF_X1 \rd_data_reg[57]$_DFFE_PP_  (.D(_0245_),
    .CK(net31),
    .Q(net183),
    .QN(_0952_));
 DFF_X1 \rd_data_reg[58]$_DFFE_PP_  (.D(_0246_),
    .CK(net31),
    .Q(net184),
    .QN(_0951_));
 DFF_X1 \rd_data_reg[59]$_DFFE_PP_  (.D(_0247_),
    .CK(net31),
    .Q(net185),
    .QN(_0950_));
 DFF_X1 \rd_data_reg[5]$_DFFE_PP_  (.D(_0248_),
    .CK(net31),
    .Q(net186),
    .QN(_0949_));
 DFF_X1 \rd_data_reg[60]$_DFFE_PP_  (.D(_0249_),
    .CK(net31),
    .Q(net187),
    .QN(_0948_));
 DFF_X1 \rd_data_reg[61]$_DFFE_PP_  (.D(_0250_),
    .CK(net31),
    .Q(net188),
    .QN(_0947_));
 DFF_X1 \rd_data_reg[62]$_DFFE_PP_  (.D(_0251_),
    .CK(net31),
    .Q(net189),
    .QN(_0946_));
 DFF_X1 \rd_data_reg[63]$_DFFE_PP_  (.D(_0252_),
    .CK(net31),
    .Q(net190),
    .QN(_0945_));
 DFF_X1 \rd_data_reg[6]$_DFFE_PP_  (.D(_0253_),
    .CK(net31),
    .Q(net191),
    .QN(_0944_));
 DFF_X1 \rd_data_reg[7]$_DFFE_PP_  (.D(_0254_),
    .CK(net31),
    .Q(net192),
    .QN(_0943_));
 DFF_X1 \rd_data_reg[8]$_DFFE_PP_  (.D(_0255_),
    .CK(net31),
    .Q(net193),
    .QN(_0942_));
 DFF_X1 \rd_data_reg[9]$_DFFE_PP_  (.D(_0256_),
    .CK(net31),
    .Q(net194),
    .QN(_0941_));
 DFF_X1 \rd_valid_reg$_SDFF_PN0_  (.D(_0257_),
    .CK(clknet_4_5_0_clk),
    .Q(net195),
    .QN(_0940_));
 DFF_X1 \refresh_counter[0]$_SDFF_PN0_  (.D(_0258_),
    .CK(clknet_4_1_0_clk),
    .Q(\refresh_counter[0] ),
    .QN(_1161_));
 DFF_X1 \refresh_counter[10]$_SDFF_PN0_  (.D(_0259_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[10] ),
    .QN(_0042_));
 DFF_X1 \refresh_counter[11]$_SDFF_PN0_  (.D(_0260_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[11] ),
    .QN(_0043_));
 DFF_X1 \refresh_counter[12]$_SDFF_PN0_  (.D(_0261_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[12] ),
    .QN(_0044_));
 DFF_X1 \refresh_counter[13]$_SDFF_PN0_  (.D(_0262_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[13] ),
    .QN(_0045_));
 DFF_X1 \refresh_counter[14]$_SDFF_PN0_  (.D(_0263_),
    .CK(clknet_4_1_0_clk),
    .Q(\refresh_counter[14] ),
    .QN(_0008_));
 DFF_X2 \refresh_counter[15]$_SDFF_PN0_  (.D(_0264_),
    .CK(clknet_4_1_0_clk),
    .Q(\refresh_counter[15] ),
    .QN(_0009_));
 DFF_X1 \refresh_counter[1]$_SDFF_PN0_  (.D(_0265_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[1] ),
    .QN(_0033_));
 DFF_X1 \refresh_counter[2]$_SDFF_PN0_  (.D(_0266_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[2] ),
    .QN(_0034_));
 DFF_X1 \refresh_counter[3]$_SDFF_PN0_  (.D(_0267_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[3] ),
    .QN(_0035_));
 DFF_X1 \refresh_counter[4]$_SDFF_PN0_  (.D(_0268_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[4] ),
    .QN(_0036_));
 DFF_X1 \refresh_counter[5]$_SDFF_PN0_  (.D(_0269_),
    .CK(clknet_4_2_0_clk),
    .Q(\refresh_counter[5] ),
    .QN(_0037_));
 DFF_X1 \refresh_counter[6]$_SDFF_PN0_  (.D(_0270_),
    .CK(clknet_4_2_0_clk),
    .Q(\refresh_counter[6] ),
    .QN(_0038_));
 DFF_X1 \refresh_counter[7]$_SDFF_PN0_  (.D(_0271_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[7] ),
    .QN(_0039_));
 DFF_X1 \refresh_counter[8]$_SDFF_PN0_  (.D(_0272_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[8] ),
    .QN(_0040_));
 DFF_X1 \refresh_counter[9]$_SDFF_PN0_  (.D(_0273_),
    .CK(clknet_4_0_0_clk),
    .Q(\refresh_counter[9] ),
    .QN(_0041_));
 DFF_X2 \timer[0]$_SDFF_PN0_  (.D(_0274_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[0] ),
    .QN(_1169_));
 DFF_X1 \timer[10]$_SDFF_PN0_  (.D(_0275_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[10] ),
    .QN(_0018_));
 DFF_X1 \timer[11]$_SDFF_PN0_  (.D(_0276_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[11] ),
    .QN(_0019_));
 DFF_X1 \timer[12]$_SDFF_PN0_  (.D(_0277_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[12] ),
    .QN(_0020_));
 DFF_X1 \timer[13]$_SDFF_PN0_  (.D(_0278_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[13] ),
    .QN(_0021_));
 DFF_X1 \timer[14]$_SDFF_PN0_  (.D(_0279_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[14] ),
    .QN(_0022_));
 DFF_X1 \timer[15]$_SDFF_PN0_  (.D(_0280_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[15] ),
    .QN(_0023_));
 DFF_X1 \timer[1]$_SDFF_PN0_  (.D(_0281_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[1] ),
    .QN(_1175_));
 DFF_X2 \timer[2]$_SDFF_PN0_  (.D(_0282_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[2] ),
    .QN(_0010_));
 DFF_X1 \timer[3]$_SDFF_PN0_  (.D(_0283_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[3] ),
    .QN(_0011_));
 DFF_X1 \timer[4]$_SDFF_PN0_  (.D(_0284_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[4] ),
    .QN(_0012_));
 DFF_X1 \timer[5]$_SDFF_PN0_  (.D(_0285_),
    .CK(clknet_4_4_0_clk),
    .Q(\timer[5] ),
    .QN(_0013_));
 DFF_X1 \timer[6]$_SDFF_PN0_  (.D(_0286_),
    .CK(clknet_4_6_0_clk),
    .Q(\timer[6] ),
    .QN(_0014_));
 DFF_X1 \timer[7]$_SDFF_PN0_  (.D(_0287_),
    .CK(clknet_4_7_0_clk),
    .Q(\timer[7] ),
    .QN(_0015_));
 DFF_X1 \timer[8]$_SDFF_PN0_  (.D(_0288_),
    .CK(clknet_4_7_0_clk),
    .Q(\timer[8] ),
    .QN(_0016_));
 DFF_X1 \timer[9]$_SDFF_PN0_  (.D(_0289_),
    .CK(clknet_4_5_0_clk),
    .Q(\timer[9] ),
    .QN(_0017_));
 DFF_X1 \wr_ready_reg$_SDFF_PN0_  (.D(_0290_),
    .CK(clknet_4_1_0_clk),
    .Q(net198),
    .QN(_0939_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_97 ();
 BUF_X1 input1 (.A(cmd_addr[0]),
    .Z(net1));
 BUF_X1 input2 (.A(cmd_addr[13]),
    .Z(net2));
 BUF_X1 input3 (.A(cmd_addr[14]),
    .Z(net3));
 BUF_X1 input4 (.A(cmd_addr[15]),
    .Z(net4));
 BUF_X1 input5 (.A(cmd_addr[16]),
    .Z(net5));
 BUF_X1 input6 (.A(cmd_addr[17]),
    .Z(net6));
 BUF_X1 input7 (.A(cmd_addr[18]),
    .Z(net7));
 BUF_X1 input8 (.A(cmd_addr[19]),
    .Z(net8));
 BUF_X1 input9 (.A(cmd_addr[1]),
    .Z(net9));
 BUF_X1 input10 (.A(cmd_addr[20]),
    .Z(net10));
 BUF_X1 input11 (.A(cmd_addr[21]),
    .Z(net11));
 BUF_X1 input12 (.A(cmd_addr[22]),
    .Z(net12));
 BUF_X1 input13 (.A(cmd_addr[23]),
    .Z(net13));
 BUF_X1 input14 (.A(cmd_addr[24]),
    .Z(net14));
 BUF_X1 input15 (.A(cmd_addr[25]),
    .Z(net15));
 BUF_X1 input16 (.A(cmd_addr[26]),
    .Z(net16));
 BUF_X1 input17 (.A(cmd_addr[27]),
    .Z(net17));
 BUF_X1 input18 (.A(cmd_addr[2]),
    .Z(net18));
 BUF_X1 input19 (.A(cmd_addr[3]),
    .Z(net19));
 BUF_X1 input20 (.A(cmd_addr[4]),
    .Z(net20));
 BUF_X1 input21 (.A(cmd_addr[5]),
    .Z(net21));
 BUF_X1 input22 (.A(cmd_addr[6]),
    .Z(net22));
 BUF_X1 input23 (.A(cmd_addr[7]),
    .Z(net23));
 BUF_X1 input24 (.A(cmd_addr[8]),
    .Z(net24));
 BUF_X1 input25 (.A(cmd_addr[9]),
    .Z(net25));
 BUF_X1 input26 (.A(cmd_burst_len[0]),
    .Z(net26));
 BUF_X1 input27 (.A(cmd_burst_len[1]),
    .Z(net27));
 BUF_X1 input28 (.A(cmd_burst_len[2]),
    .Z(net28));
 BUF_X1 input29 (.A(cmd_burst_len[3]),
    .Z(net29));
 BUF_X1 input30 (.A(cmd_write),
    .Z(net30));
 BUF_X8 input31 (.A(phy_clk),
    .Z(net31));
 BUF_X1 input32 (.A(rd_ready),
    .Z(net32));
 BUF_X1 input33 (.A(rst_n),
    .Z(net33));
 BUF_X1 input34 (.A(wr_data[0]),
    .Z(net34));
 BUF_X1 input35 (.A(wr_data[10]),
    .Z(net35));
 BUF_X1 input36 (.A(wr_data[11]),
    .Z(net36));
 BUF_X1 input37 (.A(wr_data[12]),
    .Z(net37));
 BUF_X1 input38 (.A(wr_data[13]),
    .Z(net38));
 BUF_X1 input39 (.A(wr_data[14]),
    .Z(net39));
 BUF_X1 input40 (.A(wr_data[15]),
    .Z(net40));
 BUF_X1 input41 (.A(wr_data[16]),
    .Z(net41));
 BUF_X1 input42 (.A(wr_data[17]),
    .Z(net42));
 BUF_X1 input43 (.A(wr_data[18]),
    .Z(net43));
 BUF_X1 input44 (.A(wr_data[19]),
    .Z(net44));
 BUF_X1 input45 (.A(wr_data[1]),
    .Z(net45));
 BUF_X1 input46 (.A(wr_data[20]),
    .Z(net46));
 BUF_X1 input47 (.A(wr_data[21]),
    .Z(net47));
 BUF_X1 input48 (.A(wr_data[22]),
    .Z(net48));
 BUF_X1 input49 (.A(wr_data[23]),
    .Z(net49));
 BUF_X1 input50 (.A(wr_data[24]),
    .Z(net50));
 BUF_X1 input51 (.A(wr_data[25]),
    .Z(net51));
 BUF_X1 input52 (.A(wr_data[26]),
    .Z(net52));
 BUF_X1 input53 (.A(wr_data[27]),
    .Z(net53));
 BUF_X1 input54 (.A(wr_data[28]),
    .Z(net54));
 BUF_X1 input55 (.A(wr_data[29]),
    .Z(net55));
 BUF_X1 input56 (.A(wr_data[2]),
    .Z(net56));
 BUF_X1 input57 (.A(wr_data[30]),
    .Z(net57));
 BUF_X1 input58 (.A(wr_data[31]),
    .Z(net58));
 BUF_X1 input59 (.A(wr_data[32]),
    .Z(net59));
 BUF_X1 input60 (.A(wr_data[33]),
    .Z(net60));
 BUF_X1 input61 (.A(wr_data[34]),
    .Z(net61));
 BUF_X1 input62 (.A(wr_data[35]),
    .Z(net62));
 BUF_X1 input63 (.A(wr_data[36]),
    .Z(net63));
 BUF_X1 input64 (.A(wr_data[37]),
    .Z(net64));
 BUF_X1 input65 (.A(wr_data[38]),
    .Z(net65));
 BUF_X1 input66 (.A(wr_data[39]),
    .Z(net66));
 BUF_X1 input67 (.A(wr_data[3]),
    .Z(net67));
 BUF_X1 input68 (.A(wr_data[40]),
    .Z(net68));
 BUF_X1 input69 (.A(wr_data[41]),
    .Z(net69));
 BUF_X1 input70 (.A(wr_data[42]),
    .Z(net70));
 BUF_X1 input71 (.A(wr_data[43]),
    .Z(net71));
 BUF_X1 input72 (.A(wr_data[44]),
    .Z(net72));
 BUF_X1 input73 (.A(wr_data[45]),
    .Z(net73));
 BUF_X1 input74 (.A(wr_data[46]),
    .Z(net74));
 BUF_X1 input75 (.A(wr_data[47]),
    .Z(net75));
 BUF_X1 input76 (.A(wr_data[48]),
    .Z(net76));
 BUF_X1 input77 (.A(wr_data[49]),
    .Z(net77));
 BUF_X1 input78 (.A(wr_data[4]),
    .Z(net78));
 BUF_X1 input79 (.A(wr_data[50]),
    .Z(net79));
 BUF_X1 input80 (.A(wr_data[51]),
    .Z(net80));
 BUF_X1 input81 (.A(wr_data[52]),
    .Z(net81));
 BUF_X1 input82 (.A(wr_data[53]),
    .Z(net82));
 BUF_X1 input83 (.A(wr_data[54]),
    .Z(net83));
 BUF_X1 input84 (.A(wr_data[55]),
    .Z(net84));
 BUF_X1 input85 (.A(wr_data[56]),
    .Z(net85));
 BUF_X1 input86 (.A(wr_data[57]),
    .Z(net86));
 BUF_X1 input87 (.A(wr_data[58]),
    .Z(net87));
 BUF_X1 input88 (.A(wr_data[59]),
    .Z(net88));
 BUF_X1 input89 (.A(wr_data[5]),
    .Z(net89));
 BUF_X1 input90 (.A(wr_data[60]),
    .Z(net90));
 BUF_X1 input91 (.A(wr_data[61]),
    .Z(net91));
 BUF_X1 input92 (.A(wr_data[62]),
    .Z(net92));
 BUF_X1 input93 (.A(wr_data[63]),
    .Z(net93));
 BUF_X1 input94 (.A(wr_data[6]),
    .Z(net94));
 BUF_X1 input95 (.A(wr_data[7]),
    .Z(net95));
 BUF_X1 input96 (.A(wr_data[8]),
    .Z(net96));
 BUF_X1 input97 (.A(wr_data[9]),
    .Z(net97));
 BUF_X1 input98 (.A(wr_valid),
    .Z(net98));
 BUF_X1 output99 (.A(net99),
    .Z(cmd_ready));
 BUF_X1 output100 (.A(net100),
    .Z(init_done));
 BUF_X1 output101 (.A(net101),
    .Z(phy_addr[0]));
 BUF_X1 output102 (.A(net102),
    .Z(phy_addr[10]));
 BUF_X1 output103 (.A(net103),
    .Z(phy_addr[11]));
 BUF_X1 output104 (.A(net104),
    .Z(phy_addr[12]));
 BUF_X1 output105 (.A(net105),
    .Z(phy_addr[13]));
 BUF_X1 output106 (.A(net106),
    .Z(phy_addr[1]));
 BUF_X1 output107 (.A(net107),
    .Z(phy_addr[2]));
 BUF_X1 output108 (.A(net108),
    .Z(phy_addr[3]));
 BUF_X1 output109 (.A(net109),
    .Z(phy_addr[4]));
 BUF_X1 output110 (.A(net110),
    .Z(phy_addr[5]));
 BUF_X1 output111 (.A(net111),
    .Z(phy_addr[6]));
 BUF_X1 output112 (.A(net112),
    .Z(phy_addr[7]));
 BUF_X1 output113 (.A(net113),
    .Z(phy_addr[8]));
 BUF_X1 output114 (.A(net114),
    .Z(phy_addr[9]));
 BUF_X1 output115 (.A(net115),
    .Z(phy_bank[0]));
 BUF_X1 output116 (.A(net116),
    .Z(phy_bank[1]));
 BUF_X1 output117 (.A(net117),
    .Z(phy_bank[2]));
 BUF_X1 output118 (.A(net118),
    .Z(phy_cas_n));
 BUF_X1 output119 (.A(net119),
    .Z(phy_cs_n));
 BUF_X1 output120 (.A(net120),
    .Z(phy_dm[0]));
 BUF_X1 output121 (.A(net121),
    .Z(phy_dm[1]));
 BUF_X1 output122 (.A(net122),
    .Z(phy_dm[2]));
 BUF_X1 output123 (.A(net123),
    .Z(phy_dm[3]));
 BUF_X1 output124 (.A(net124),
    .Z(phy_dm[4]));
 BUF_X1 output125 (.A(net125),
    .Z(phy_dm[5]));
 BUF_X1 output126 (.A(net126),
    .Z(phy_dm[6]));
 BUF_X1 output127 (.A(net127),
    .Z(phy_dm[7]));
 BUF_X1 output128 (.A(net128),
    .Z(phy_ras_n));
 BUF_X1 output129 (.A(net129),
    .Z(phy_reset_n));
 BUF_X1 output130 (.A(net130),
    .Z(phy_we_n));
 BUF_X1 output131 (.A(net131),
    .Z(rd_data[0]));
 BUF_X1 output132 (.A(net132),
    .Z(rd_data[10]));
 BUF_X1 output133 (.A(net133),
    .Z(rd_data[11]));
 BUF_X1 output134 (.A(net134),
    .Z(rd_data[12]));
 BUF_X1 output135 (.A(net135),
    .Z(rd_data[13]));
 BUF_X1 output136 (.A(net136),
    .Z(rd_data[14]));
 BUF_X1 output137 (.A(net137),
    .Z(rd_data[15]));
 BUF_X1 output138 (.A(net138),
    .Z(rd_data[16]));
 BUF_X1 output139 (.A(net139),
    .Z(rd_data[17]));
 BUF_X1 output140 (.A(net140),
    .Z(rd_data[18]));
 BUF_X1 output141 (.A(net141),
    .Z(rd_data[19]));
 BUF_X1 output142 (.A(net142),
    .Z(rd_data[1]));
 BUF_X1 output143 (.A(net143),
    .Z(rd_data[20]));
 BUF_X1 output144 (.A(net144),
    .Z(rd_data[21]));
 BUF_X1 output145 (.A(net145),
    .Z(rd_data[22]));
 BUF_X1 output146 (.A(net146),
    .Z(rd_data[23]));
 BUF_X1 output147 (.A(net147),
    .Z(rd_data[24]));
 BUF_X1 output148 (.A(net148),
    .Z(rd_data[25]));
 BUF_X1 output149 (.A(net149),
    .Z(rd_data[26]));
 BUF_X1 output150 (.A(net150),
    .Z(rd_data[27]));
 BUF_X1 output151 (.A(net151),
    .Z(rd_data[28]));
 BUF_X1 output152 (.A(net152),
    .Z(rd_data[29]));
 BUF_X1 output153 (.A(net153),
    .Z(rd_data[2]));
 BUF_X1 output154 (.A(net154),
    .Z(rd_data[30]));
 BUF_X1 output155 (.A(net155),
    .Z(rd_data[31]));
 BUF_X1 output156 (.A(net156),
    .Z(rd_data[32]));
 BUF_X1 output157 (.A(net157),
    .Z(rd_data[33]));
 BUF_X1 output158 (.A(net158),
    .Z(rd_data[34]));
 BUF_X1 output159 (.A(net159),
    .Z(rd_data[35]));
 BUF_X1 output160 (.A(net160),
    .Z(rd_data[36]));
 BUF_X1 output161 (.A(net161),
    .Z(rd_data[37]));
 BUF_X1 output162 (.A(net162),
    .Z(rd_data[38]));
 BUF_X1 output163 (.A(net163),
    .Z(rd_data[39]));
 BUF_X1 output164 (.A(net164),
    .Z(rd_data[3]));
 BUF_X1 output165 (.A(net165),
    .Z(rd_data[40]));
 BUF_X1 output166 (.A(net166),
    .Z(rd_data[41]));
 BUF_X1 output167 (.A(net167),
    .Z(rd_data[42]));
 BUF_X1 output168 (.A(net168),
    .Z(rd_data[43]));
 BUF_X1 output169 (.A(net169),
    .Z(rd_data[44]));
 BUF_X1 output170 (.A(net170),
    .Z(rd_data[45]));
 BUF_X1 output171 (.A(net171),
    .Z(rd_data[46]));
 BUF_X1 output172 (.A(net172),
    .Z(rd_data[47]));
 BUF_X1 output173 (.A(net173),
    .Z(rd_data[48]));
 BUF_X1 output174 (.A(net174),
    .Z(rd_data[49]));
 BUF_X1 output175 (.A(net175),
    .Z(rd_data[4]));
 BUF_X1 output176 (.A(net176),
    .Z(rd_data[50]));
 BUF_X1 output177 (.A(net177),
    .Z(rd_data[51]));
 BUF_X1 output178 (.A(net178),
    .Z(rd_data[52]));
 BUF_X1 output179 (.A(net179),
    .Z(rd_data[53]));
 BUF_X1 output180 (.A(net180),
    .Z(rd_data[54]));
 BUF_X1 output181 (.A(net181),
    .Z(rd_data[55]));
 BUF_X1 output182 (.A(net182),
    .Z(rd_data[56]));
 BUF_X1 output183 (.A(net183),
    .Z(rd_data[57]));
 BUF_X1 output184 (.A(net184),
    .Z(rd_data[58]));
 BUF_X1 output185 (.A(net185),
    .Z(rd_data[59]));
 BUF_X1 output186 (.A(net186),
    .Z(rd_data[5]));
 BUF_X1 output187 (.A(net187),
    .Z(rd_data[60]));
 BUF_X1 output188 (.A(net188),
    .Z(rd_data[61]));
 BUF_X1 output189 (.A(net189),
    .Z(rd_data[62]));
 BUF_X1 output190 (.A(net190),
    .Z(rd_data[63]));
 BUF_X1 output191 (.A(net191),
    .Z(rd_data[6]));
 BUF_X1 output192 (.A(net192),
    .Z(rd_data[7]));
 BUF_X1 output193 (.A(net193),
    .Z(rd_data[8]));
 BUF_X1 output194 (.A(net194),
    .Z(rd_data[9]));
 BUF_X1 output195 (.A(net195),
    .Z(rd_valid));
 BUF_X1 output196 (.A(net196),
    .Z(state[0]));
 BUF_X1 output197 (.A(net197),
    .Z(state[1]));
 BUF_X1 output198 (.A(net198),
    .Z(wr_ready));
 LOGIC0_X1 _2116__199 (.Z(net199));
 LOGIC0_X1 _2117__200 (.Z(net200));
 LOGIC0_X1 _2191__201 (.Z(net201));
 LOGIC0_X1 _2192__202 (.Z(net202));
 LOGIC0_X1 _2193__203 (.Z(net203));
 LOGIC0_X1 _2194__204 (.Z(net204));
 LOGIC0_X1 _2195__205 (.Z(net205));
 LOGIC0_X1 _2196__206 (.Z(net206));
 LOGIC0_X1 _2197__207 (.Z(net207));
 LOGIC0_X1 _2198__208 (.Z(net208));
 LOGIC1_X1 _2199__210 (.Z(net210));
 LOGIC1_X1 _2200__211 (.Z(net211));
 LOGIC1_X1 _2201__212 (.Z(net212));
 LOGIC1_X1 _2202__213 (.Z(net213));
 LOGIC1_X1 _2203__214 (.Z(net214));
 LOGIC1_X1 _2204__215 (.Z(net215));
 LOGIC1_X1 _2205__216 (.Z(net216));
 LOGIC1_X1 _2206__217 (.Z(net217));
 LOGIC1_X1 _2207__218 (.Z(net218));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 INV_X4 clkload0 (.A(clknet_4_0_0_clk));
 INV_X4 clkload1 (.A(clknet_4_1_0_clk));
 INV_X4 clkload2 (.A(clknet_4_2_0_clk));
 INV_X4 clkload3 (.A(clknet_4_3_0_clk));
 INV_X8 clkload4 (.A(clknet_4_4_0_clk));
 INV_X4 clkload5 (.A(clknet_4_5_0_clk));
 INV_X8 clkload6 (.A(clknet_4_6_0_clk));
 INV_X8 clkload7 (.A(clknet_4_7_0_clk));
 INV_X4 clkload8 (.A(clknet_4_8_0_clk));
 INV_X4 clkload9 (.A(clknet_4_9_0_clk));
 INV_X2 clkload10 (.A(clknet_4_11_0_clk));
 INV_X4 clkload11 (.A(clknet_4_12_0_clk));
 INV_X4 clkload12 (.A(clknet_4_13_0_clk));
 INV_X1 clkload13 (.A(clknet_4_14_0_clk));
 INV_X4 clkload14 (.A(clknet_4_15_0_clk));
 FILLCELL_X1 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_8 ();
 FILLCELL_X16 FILLER_0_40 ();
 FILLCELL_X2 FILLER_0_56 ();
 FILLCELL_X1 FILLER_0_58 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X4 FILLER_0_81 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X16 FILLER_0_92 ();
 FILLCELL_X4 FILLER_0_108 ();
 FILLCELL_X2 FILLER_0_112 ();
 FILLCELL_X1 FILLER_0_114 ();
 FILLCELL_X32 FILLER_0_118 ();
 FILLCELL_X1 FILLER_0_182 ();
 FILLCELL_X2 FILLER_0_208 ();
 FILLCELL_X4 FILLER_0_223 ();
 FILLCELL_X2 FILLER_0_227 ();
 FILLCELL_X16 FILLER_0_246 ();
 FILLCELL_X4 FILLER_0_262 ();
 FILLCELL_X1 FILLER_0_266 ();
 FILLCELL_X16 FILLER_0_284 ();
 FILLCELL_X4 FILLER_0_300 ();
 FILLCELL_X2 FILLER_0_304 ();
 FILLCELL_X1 FILLER_0_306 ();
 FILLCELL_X32 FILLER_0_313 ();
 FILLCELL_X16 FILLER_0_345 ();
 FILLCELL_X4 FILLER_0_361 ();
 FILLCELL_X2 FILLER_0_365 ();
 FILLCELL_X1 FILLER_0_367 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_97 ();
 FILLCELL_X4 FILLER_1_105 ();
 FILLCELL_X2 FILLER_1_109 ();
 FILLCELL_X32 FILLER_1_114 ();
 FILLCELL_X1 FILLER_1_146 ();
 FILLCELL_X4 FILLER_1_232 ();
 FILLCELL_X1 FILLER_1_243 ();
 FILLCELL_X1 FILLER_1_268 ();
 FILLCELL_X4 FILLER_1_276 ();
 FILLCELL_X2 FILLER_1_280 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X8 FILLER_1_353 ();
 FILLCELL_X4 FILLER_1_361 ();
 FILLCELL_X2 FILLER_1_365 ();
 FILLCELL_X1 FILLER_1_367 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X16 FILLER_2_97 ();
 FILLCELL_X8 FILLER_2_113 ();
 FILLCELL_X4 FILLER_2_121 ();
 FILLCELL_X2 FILLER_2_125 ();
 FILLCELL_X2 FILLER_2_151 ();
 FILLCELL_X8 FILLER_2_170 ();
 FILLCELL_X2 FILLER_2_178 ();
 FILLCELL_X8 FILLER_2_186 ();
 FILLCELL_X4 FILLER_2_194 ();
 FILLCELL_X16 FILLER_2_200 ();
 FILLCELL_X4 FILLER_2_216 ();
 FILLCELL_X2 FILLER_2_220 ();
 FILLCELL_X1 FILLER_2_222 ();
 FILLCELL_X4 FILLER_2_244 ();
 FILLCELL_X2 FILLER_2_248 ();
 FILLCELL_X16 FILLER_2_267 ();
 FILLCELL_X1 FILLER_2_300 ();
 FILLCELL_X32 FILLER_2_325 ();
 FILLCELL_X8 FILLER_2_357 ();
 FILLCELL_X2 FILLER_2_365 ();
 FILLCELL_X1 FILLER_2_367 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X4 FILLER_3_129 ();
 FILLCELL_X2 FILLER_3_133 ();
 FILLCELL_X1 FILLER_3_135 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X2 FILLER_3_157 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X4 FILLER_3_174 ();
 FILLCELL_X2 FILLER_3_178 ();
 FILLCELL_X1 FILLER_3_180 ();
 FILLCELL_X2 FILLER_3_188 ();
 FILLCELL_X4 FILLER_3_218 ();
 FILLCELL_X2 FILLER_3_229 ();
 FILLCELL_X4 FILLER_3_244 ();
 FILLCELL_X1 FILLER_3_248 ();
 FILLCELL_X8 FILLER_3_256 ();
 FILLCELL_X2 FILLER_3_264 ();
 FILLCELL_X1 FILLER_3_266 ();
 FILLCELL_X4 FILLER_3_274 ();
 FILLCELL_X2 FILLER_3_285 ();
 FILLCELL_X1 FILLER_3_287 ();
 FILLCELL_X8 FILLER_3_295 ();
 FILLCELL_X4 FILLER_3_303 ();
 FILLCELL_X2 FILLER_3_307 ();
 FILLCELL_X2 FILLER_3_316 ();
 FILLCELL_X4 FILLER_3_339 ();
 FILLCELL_X16 FILLER_3_350 ();
 FILLCELL_X2 FILLER_3_366 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X16 FILLER_4_33 ();
 FILLCELL_X8 FILLER_4_49 ();
 FILLCELL_X4 FILLER_4_57 ();
 FILLCELL_X1 FILLER_4_61 ();
 FILLCELL_X32 FILLER_4_71 ();
 FILLCELL_X32 FILLER_4_103 ();
 FILLCELL_X8 FILLER_4_135 ();
 FILLCELL_X16 FILLER_4_157 ();
 FILLCELL_X2 FILLER_4_173 ();
 FILLCELL_X1 FILLER_4_175 ();
 FILLCELL_X8 FILLER_4_193 ();
 FILLCELL_X4 FILLER_4_201 ();
 FILLCELL_X4 FILLER_4_236 ();
 FILLCELL_X2 FILLER_4_247 ();
 FILLCELL_X8 FILLER_4_256 ();
 FILLCELL_X2 FILLER_4_264 ();
 FILLCELL_X4 FILLER_4_283 ();
 FILLCELL_X2 FILLER_4_304 ();
 FILLCELL_X2 FILLER_4_323 ();
 FILLCELL_X4 FILLER_4_327 ();
 FILLCELL_X2 FILLER_4_331 ();
 FILLCELL_X2 FILLER_4_340 ();
 FILLCELL_X2 FILLER_4_359 ();
 FILLCELL_X1 FILLER_4_367 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_17 ();
 FILLCELL_X1 FILLER_5_21 ();
 FILLCELL_X1 FILLER_5_39 ();
 FILLCELL_X32 FILLER_5_75 ();
 FILLCELL_X32 FILLER_5_107 ();
 FILLCELL_X2 FILLER_5_139 ();
 FILLCELL_X1 FILLER_5_141 ();
 FILLCELL_X1 FILLER_5_149 ();
 FILLCELL_X4 FILLER_5_157 ();
 FILLCELL_X8 FILLER_5_185 ();
 FILLCELL_X2 FILLER_5_203 ();
 FILLCELL_X8 FILLER_5_212 ();
 FILLCELL_X2 FILLER_5_220 ();
 FILLCELL_X16 FILLER_5_260 ();
 FILLCELL_X8 FILLER_5_276 ();
 FILLCELL_X4 FILLER_5_288 ();
 FILLCELL_X16 FILLER_5_299 ();
 FILLCELL_X8 FILLER_5_315 ();
 FILLCELL_X1 FILLER_5_323 ();
 FILLCELL_X4 FILLER_5_346 ();
 FILLCELL_X2 FILLER_5_350 ();
 FILLCELL_X8 FILLER_5_359 ();
 FILLCELL_X1 FILLER_5_367 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_17 ();
 FILLCELL_X4 FILLER_6_25 ();
 FILLCELL_X2 FILLER_6_29 ();
 FILLCELL_X2 FILLER_6_36 ();
 FILLCELL_X1 FILLER_6_45 ();
 FILLCELL_X32 FILLER_6_86 ();
 FILLCELL_X8 FILLER_6_118 ();
 FILLCELL_X4 FILLER_6_126 ();
 FILLCELL_X1 FILLER_6_130 ();
 FILLCELL_X2 FILLER_6_148 ();
 FILLCELL_X1 FILLER_6_150 ();
 FILLCELL_X4 FILLER_6_168 ();
 FILLCELL_X1 FILLER_6_172 ();
 FILLCELL_X2 FILLER_6_180 ();
 FILLCELL_X4 FILLER_6_189 ();
 FILLCELL_X1 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_213 ();
 FILLCELL_X2 FILLER_6_245 ();
 FILLCELL_X2 FILLER_6_265 ();
 FILLCELL_X1 FILLER_6_267 ();
 FILLCELL_X4 FILLER_6_301 ();
 FILLCELL_X2 FILLER_6_305 ();
 FILLCELL_X1 FILLER_6_307 ();
 FILLCELL_X4 FILLER_6_325 ();
 FILLCELL_X2 FILLER_6_329 ();
 FILLCELL_X1 FILLER_6_331 ();
 FILLCELL_X8 FILLER_6_339 ();
 FILLCELL_X4 FILLER_6_347 ();
 FILLCELL_X16 FILLER_7_1 ();
 FILLCELL_X4 FILLER_7_17 ();
 FILLCELL_X2 FILLER_7_21 ();
 FILLCELL_X8 FILLER_7_46 ();
 FILLCELL_X4 FILLER_7_54 ();
 FILLCELL_X2 FILLER_7_58 ();
 FILLCELL_X1 FILLER_7_60 ();
 FILLCELL_X4 FILLER_7_72 ();
 FILLCELL_X32 FILLER_7_96 ();
 FILLCELL_X8 FILLER_7_128 ();
 FILLCELL_X4 FILLER_7_136 ();
 FILLCELL_X2 FILLER_7_140 ();
 FILLCELL_X1 FILLER_7_142 ();
 FILLCELL_X16 FILLER_7_150 ();
 FILLCELL_X8 FILLER_7_166 ();
 FILLCELL_X4 FILLER_7_181 ();
 FILLCELL_X2 FILLER_7_185 ();
 FILLCELL_X1 FILLER_7_194 ();
 FILLCELL_X2 FILLER_7_211 ();
 FILLCELL_X2 FILLER_7_230 ();
 FILLCELL_X4 FILLER_7_246 ();
 FILLCELL_X4 FILLER_7_268 ();
 FILLCELL_X2 FILLER_7_279 ();
 FILLCELL_X1 FILLER_7_281 ();
 FILLCELL_X8 FILLER_7_296 ();
 FILLCELL_X2 FILLER_7_304 ();
 FILLCELL_X8 FILLER_7_313 ();
 FILLCELL_X2 FILLER_7_321 ();
 FILLCELL_X8 FILLER_7_358 ();
 FILLCELL_X2 FILLER_7_366 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_17 ();
 FILLCELL_X4 FILLER_8_33 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X4 FILLER_8_73 ();
 FILLCELL_X1 FILLER_8_77 ();
 FILLCELL_X2 FILLER_8_82 ();
 FILLCELL_X32 FILLER_8_90 ();
 FILLCELL_X8 FILLER_8_122 ();
 FILLCELL_X2 FILLER_8_130 ();
 FILLCELL_X2 FILLER_8_173 ();
 FILLCELL_X1 FILLER_8_175 ();
 FILLCELL_X2 FILLER_8_179 ();
 FILLCELL_X1 FILLER_8_181 ();
 FILLCELL_X4 FILLER_8_187 ();
 FILLCELL_X8 FILLER_8_201 ();
 FILLCELL_X4 FILLER_8_209 ();
 FILLCELL_X2 FILLER_8_220 ();
 FILLCELL_X1 FILLER_8_222 ();
 FILLCELL_X8 FILLER_8_256 ();
 FILLCELL_X2 FILLER_8_264 ();
 FILLCELL_X1 FILLER_8_266 ();
 FILLCELL_X4 FILLER_8_274 ();
 FILLCELL_X2 FILLER_8_278 ();
 FILLCELL_X16 FILLER_8_297 ();
 FILLCELL_X8 FILLER_8_313 ();
 FILLCELL_X4 FILLER_8_338 ();
 FILLCELL_X2 FILLER_8_342 ();
 FILLCELL_X1 FILLER_8_344 ();
 FILLCELL_X4 FILLER_8_362 ();
 FILLCELL_X2 FILLER_8_366 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_9 ();
 FILLCELL_X1 FILLER_9_11 ();
 FILLCELL_X1 FILLER_9_32 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X4 FILLER_9_69 ();
 FILLCELL_X1 FILLER_9_77 ();
 FILLCELL_X32 FILLER_9_98 ();
 FILLCELL_X2 FILLER_9_130 ();
 FILLCELL_X1 FILLER_9_132 ();
 FILLCELL_X1 FILLER_9_150 ();
 FILLCELL_X2 FILLER_9_168 ();
 FILLCELL_X1 FILLER_9_170 ();
 FILLCELL_X1 FILLER_9_188 ();
 FILLCELL_X2 FILLER_9_196 ();
 FILLCELL_X8 FILLER_9_205 ();
 FILLCELL_X1 FILLER_9_213 ();
 FILLCELL_X2 FILLER_9_221 ();
 FILLCELL_X1 FILLER_9_223 ();
 FILLCELL_X8 FILLER_9_231 ();
 FILLCELL_X2 FILLER_9_239 ();
 FILLCELL_X16 FILLER_9_248 ();
 FILLCELL_X2 FILLER_9_281 ();
 FILLCELL_X1 FILLER_9_283 ();
 FILLCELL_X8 FILLER_9_291 ();
 FILLCELL_X4 FILLER_9_299 ();
 FILLCELL_X1 FILLER_9_303 ();
 FILLCELL_X4 FILLER_9_311 ();
 FILLCELL_X8 FILLER_9_329 ();
 FILLCELL_X2 FILLER_9_337 ();
 FILLCELL_X1 FILLER_9_339 ();
 FILLCELL_X4 FILLER_9_347 ();
 FILLCELL_X1 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_19 ();
 FILLCELL_X1 FILLER_10_23 ();
 FILLCELL_X1 FILLER_10_41 ();
 FILLCELL_X4 FILLER_10_55 ();
 FILLCELL_X1 FILLER_10_59 ();
 FILLCELL_X1 FILLER_10_67 ();
 FILLCELL_X32 FILLER_10_79 ();
 FILLCELL_X4 FILLER_10_111 ();
 FILLCELL_X4 FILLER_10_122 ();
 FILLCELL_X4 FILLER_10_150 ();
 FILLCELL_X1 FILLER_10_154 ();
 FILLCELL_X2 FILLER_10_162 ();
 FILLCELL_X4 FILLER_10_171 ();
 FILLCELL_X2 FILLER_10_175 ();
 FILLCELL_X2 FILLER_10_181 ();
 FILLCELL_X1 FILLER_10_194 ();
 FILLCELL_X2 FILLER_10_198 ();
 FILLCELL_X8 FILLER_10_203 ();
 FILLCELL_X4 FILLER_10_211 ();
 FILLCELL_X2 FILLER_10_215 ();
 FILLCELL_X1 FILLER_10_217 ();
 FILLCELL_X4 FILLER_10_225 ();
 FILLCELL_X8 FILLER_10_261 ();
 FILLCELL_X4 FILLER_10_269 ();
 FILLCELL_X2 FILLER_10_273 ();
 FILLCELL_X1 FILLER_10_275 ();
 FILLCELL_X8 FILLER_10_324 ();
 FILLCELL_X4 FILLER_10_332 ();
 FILLCELL_X2 FILLER_10_336 ();
 FILLCELL_X4 FILLER_10_362 ();
 FILLCELL_X2 FILLER_10_366 ();
 FILLCELL_X4 FILLER_11_22 ();
 FILLCELL_X2 FILLER_11_26 ();
 FILLCELL_X8 FILLER_11_31 ();
 FILLCELL_X4 FILLER_11_39 ();
 FILLCELL_X1 FILLER_11_60 ();
 FILLCELL_X16 FILLER_11_74 ();
 FILLCELL_X2 FILLER_11_90 ();
 FILLCELL_X4 FILLER_11_111 ();
 FILLCELL_X4 FILLER_11_132 ();
 FILLCELL_X2 FILLER_11_146 ();
 FILLCELL_X1 FILLER_11_148 ();
 FILLCELL_X8 FILLER_11_180 ();
 FILLCELL_X4 FILLER_11_188 ();
 FILLCELL_X1 FILLER_11_192 ();
 FILLCELL_X1 FILLER_11_257 ();
 FILLCELL_X4 FILLER_11_265 ();
 FILLCELL_X1 FILLER_11_269 ();
 FILLCELL_X8 FILLER_11_277 ();
 FILLCELL_X16 FILLER_11_288 ();
 FILLCELL_X4 FILLER_11_304 ();
 FILLCELL_X2 FILLER_11_308 ();
 FILLCELL_X4 FILLER_11_315 ();
 FILLCELL_X8 FILLER_11_336 ();
 FILLCELL_X1 FILLER_11_344 ();
 FILLCELL_X16 FILLER_11_352 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X4 FILLER_12_33 ();
 FILLCELL_X2 FILLER_12_37 ();
 FILLCELL_X2 FILLER_12_56 ();
 FILLCELL_X1 FILLER_12_58 ();
 FILLCELL_X2 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_68 ();
 FILLCELL_X16 FILLER_12_74 ();
 FILLCELL_X4 FILLER_12_90 ();
 FILLCELL_X1 FILLER_12_94 ();
 FILLCELL_X16 FILLER_12_99 ();
 FILLCELL_X2 FILLER_12_115 ();
 FILLCELL_X4 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_146 ();
 FILLCELL_X4 FILLER_12_155 ();
 FILLCELL_X2 FILLER_12_159 ();
 FILLCELL_X1 FILLER_12_161 ();
 FILLCELL_X1 FILLER_12_179 ();
 FILLCELL_X4 FILLER_12_189 ();
 FILLCELL_X2 FILLER_12_193 ();
 FILLCELL_X8 FILLER_12_213 ();
 FILLCELL_X4 FILLER_12_221 ();
 FILLCELL_X2 FILLER_12_262 ();
 FILLCELL_X4 FILLER_12_268 ();
 FILLCELL_X1 FILLER_12_272 ();
 FILLCELL_X8 FILLER_12_304 ();
 FILLCELL_X2 FILLER_12_323 ();
 FILLCELL_X2 FILLER_12_329 ();
 FILLCELL_X1 FILLER_12_331 ();
 FILLCELL_X2 FILLER_12_339 ();
 FILLCELL_X1 FILLER_12_341 ();
 FILLCELL_X2 FILLER_12_366 ();
 FILLCELL_X1 FILLER_13_1 ();
 FILLCELL_X16 FILLER_13_5 ();
 FILLCELL_X4 FILLER_13_21 ();
 FILLCELL_X1 FILLER_13_25 ();
 FILLCELL_X2 FILLER_13_56 ();
 FILLCELL_X1 FILLER_13_58 ();
 FILLCELL_X4 FILLER_13_69 ();
 FILLCELL_X2 FILLER_13_73 ();
 FILLCELL_X2 FILLER_13_96 ();
 FILLCELL_X2 FILLER_13_105 ();
 FILLCELL_X1 FILLER_13_107 ();
 FILLCELL_X8 FILLER_13_119 ();
 FILLCELL_X2 FILLER_13_127 ();
 FILLCELL_X2 FILLER_13_134 ();
 FILLCELL_X4 FILLER_13_162 ();
 FILLCELL_X1 FILLER_13_166 ();
 FILLCELL_X2 FILLER_13_198 ();
 FILLCELL_X1 FILLER_13_200 ();
 FILLCELL_X8 FILLER_13_205 ();
 FILLCELL_X4 FILLER_13_220 ();
 FILLCELL_X2 FILLER_13_224 ();
 FILLCELL_X1 FILLER_13_226 ();
 FILLCELL_X4 FILLER_13_234 ();
 FILLCELL_X2 FILLER_13_238 ();
 FILLCELL_X1 FILLER_13_240 ();
 FILLCELL_X8 FILLER_13_255 ();
 FILLCELL_X2 FILLER_13_263 ();
 FILLCELL_X16 FILLER_13_269 ();
 FILLCELL_X8 FILLER_13_285 ();
 FILLCELL_X2 FILLER_13_293 ();
 FILLCELL_X1 FILLER_13_295 ();
 FILLCELL_X1 FILLER_13_310 ();
 FILLCELL_X1 FILLER_13_314 ();
 FILLCELL_X1 FILLER_13_324 ();
 FILLCELL_X1 FILLER_13_329 ();
 FILLCELL_X8 FILLER_13_354 ();
 FILLCELL_X4 FILLER_13_362 ();
 FILLCELL_X2 FILLER_13_366 ();
 FILLCELL_X4 FILLER_14_18 ();
 FILLCELL_X16 FILLER_14_68 ();
 FILLCELL_X4 FILLER_14_84 ();
 FILLCELL_X2 FILLER_14_88 ();
 FILLCELL_X2 FILLER_14_93 ();
 FILLCELL_X1 FILLER_14_95 ();
 FILLCELL_X1 FILLER_14_114 ();
 FILLCELL_X4 FILLER_14_132 ();
 FILLCELL_X2 FILLER_14_163 ();
 FILLCELL_X1 FILLER_14_165 ();
 FILLCELL_X4 FILLER_14_180 ();
 FILLCELL_X1 FILLER_14_184 ();
 FILLCELL_X4 FILLER_14_202 ();
 FILLCELL_X1 FILLER_14_206 ();
 FILLCELL_X4 FILLER_14_224 ();
 FILLCELL_X4 FILLER_14_271 ();
 FILLCELL_X2 FILLER_14_292 ();
 FILLCELL_X1 FILLER_14_294 ();
 FILLCELL_X1 FILLER_14_302 ();
 FILLCELL_X1 FILLER_14_320 ();
 FILLCELL_X16 FILLER_14_338 ();
 FILLCELL_X8 FILLER_14_354 ();
 FILLCELL_X4 FILLER_14_362 ();
 FILLCELL_X2 FILLER_14_366 ();
 FILLCELL_X8 FILLER_15_4 ();
 FILLCELL_X4 FILLER_15_12 ();
 FILLCELL_X8 FILLER_15_19 ();
 FILLCELL_X2 FILLER_15_27 ();
 FILLCELL_X1 FILLER_15_29 ();
 FILLCELL_X1 FILLER_15_42 ();
 FILLCELL_X1 FILLER_15_58 ();
 FILLCELL_X1 FILLER_15_62 ();
 FILLCELL_X8 FILLER_15_73 ();
 FILLCELL_X4 FILLER_15_81 ();
 FILLCELL_X2 FILLER_15_85 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X2 FILLER_15_117 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X4 FILLER_15_125 ();
 FILLCELL_X1 FILLER_15_129 ();
 FILLCELL_X2 FILLER_15_151 ();
 FILLCELL_X2 FILLER_15_167 ();
 FILLCELL_X2 FILLER_15_172 ();
 FILLCELL_X1 FILLER_15_174 ();
 FILLCELL_X16 FILLER_15_189 ();
 FILLCELL_X4 FILLER_15_205 ();
 FILLCELL_X2 FILLER_15_209 ();
 FILLCELL_X8 FILLER_15_225 ();
 FILLCELL_X4 FILLER_15_233 ();
 FILLCELL_X2 FILLER_15_237 ();
 FILLCELL_X16 FILLER_15_242 ();
 FILLCELL_X8 FILLER_15_258 ();
 FILLCELL_X4 FILLER_15_266 ();
 FILLCELL_X1 FILLER_15_277 ();
 FILLCELL_X8 FILLER_15_285 ();
 FILLCELL_X2 FILLER_15_293 ();
 FILLCELL_X4 FILLER_15_302 ();
 FILLCELL_X2 FILLER_15_306 ();
 FILLCELL_X1 FILLER_15_308 ();
 FILLCELL_X4 FILLER_15_316 ();
 FILLCELL_X2 FILLER_15_320 ();
 FILLCELL_X4 FILLER_15_329 ();
 FILLCELL_X4 FILLER_15_340 ();
 FILLCELL_X1 FILLER_15_344 ();
 FILLCELL_X16 FILLER_15_352 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_9 ();
 FILLCELL_X1 FILLER_16_11 ();
 FILLCELL_X8 FILLER_16_29 ();
 FILLCELL_X4 FILLER_16_37 ();
 FILLCELL_X8 FILLER_16_44 ();
 FILLCELL_X2 FILLER_16_52 ();
 FILLCELL_X4 FILLER_16_65 ();
 FILLCELL_X2 FILLER_16_69 ();
 FILLCELL_X1 FILLER_16_71 ();
 FILLCELL_X4 FILLER_16_93 ();
 FILLCELL_X2 FILLER_16_97 ();
 FILLCELL_X1 FILLER_16_142 ();
 FILLCELL_X4 FILLER_16_159 ();
 FILLCELL_X1 FILLER_16_163 ();
 FILLCELL_X16 FILLER_16_182 ();
 FILLCELL_X4 FILLER_16_198 ();
 FILLCELL_X4 FILLER_16_219 ();
 FILLCELL_X1 FILLER_16_223 ();
 FILLCELL_X16 FILLER_16_241 ();
 FILLCELL_X4 FILLER_16_257 ();
 FILLCELL_X2 FILLER_16_261 ();
 FILLCELL_X1 FILLER_16_263 ();
 FILLCELL_X4 FILLER_16_288 ();
 FILLCELL_X1 FILLER_16_326 ();
 FILLCELL_X4 FILLER_16_331 ();
 FILLCELL_X16 FILLER_16_352 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X16 FILLER_17_9 ();
 FILLCELL_X1 FILLER_17_25 ();
 FILLCELL_X2 FILLER_17_56 ();
 FILLCELL_X4 FILLER_17_78 ();
 FILLCELL_X2 FILLER_17_82 ();
 FILLCELL_X1 FILLER_17_91 ();
 FILLCELL_X8 FILLER_17_96 ();
 FILLCELL_X4 FILLER_17_104 ();
 FILLCELL_X1 FILLER_17_108 ();
 FILLCELL_X8 FILLER_17_114 ();
 FILLCELL_X4 FILLER_17_122 ();
 FILLCELL_X1 FILLER_17_126 ();
 FILLCELL_X1 FILLER_17_146 ();
 FILLCELL_X1 FILLER_17_152 ();
 FILLCELL_X2 FILLER_17_156 ();
 FILLCELL_X8 FILLER_17_163 ();
 FILLCELL_X4 FILLER_17_171 ();
 FILLCELL_X2 FILLER_17_175 ();
 FILLCELL_X1 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_199 ();
 FILLCELL_X1 FILLER_17_201 ();
 FILLCELL_X4 FILLER_17_224 ();
 FILLCELL_X2 FILLER_17_228 ();
 FILLCELL_X2 FILLER_17_237 ();
 FILLCELL_X1 FILLER_17_239 ();
 FILLCELL_X4 FILLER_17_247 ();
 FILLCELL_X1 FILLER_17_251 ();
 FILLCELL_X16 FILLER_17_259 ();
 FILLCELL_X8 FILLER_17_275 ();
 FILLCELL_X2 FILLER_17_283 ();
 FILLCELL_X4 FILLER_17_292 ();
 FILLCELL_X2 FILLER_17_296 ();
 FILLCELL_X1 FILLER_17_298 ();
 FILLCELL_X8 FILLER_17_306 ();
 FILLCELL_X4 FILLER_17_314 ();
 FILLCELL_X2 FILLER_17_318 ();
 FILLCELL_X1 FILLER_17_320 ();
 FILLCELL_X1 FILLER_17_330 ();
 FILLCELL_X2 FILLER_17_338 ();
 FILLCELL_X1 FILLER_17_367 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X2 FILLER_18_24 ();
 FILLCELL_X1 FILLER_18_26 ();
 FILLCELL_X1 FILLER_18_37 ();
 FILLCELL_X4 FILLER_18_52 ();
 FILLCELL_X2 FILLER_18_56 ();
 FILLCELL_X8 FILLER_18_61 ();
 FILLCELL_X2 FILLER_18_69 ();
 FILLCELL_X1 FILLER_18_71 ();
 FILLCELL_X1 FILLER_18_83 ();
 FILLCELL_X1 FILLER_18_107 ();
 FILLCELL_X8 FILLER_18_112 ();
 FILLCELL_X4 FILLER_18_120 ();
 FILLCELL_X2 FILLER_18_124 ();
 FILLCELL_X4 FILLER_18_134 ();
 FILLCELL_X1 FILLER_18_138 ();
 FILLCELL_X2 FILLER_18_144 ();
 FILLCELL_X4 FILLER_18_168 ();
 FILLCELL_X2 FILLER_18_172 ();
 FILLCELL_X1 FILLER_18_174 ();
 FILLCELL_X2 FILLER_18_190 ();
 FILLCELL_X4 FILLER_18_197 ();
 FILLCELL_X1 FILLER_18_201 ();
 FILLCELL_X4 FILLER_18_223 ();
 FILLCELL_X1 FILLER_18_227 ();
 FILLCELL_X4 FILLER_18_235 ();
 FILLCELL_X2 FILLER_18_239 ();
 FILLCELL_X8 FILLER_18_262 ();
 FILLCELL_X1 FILLER_18_270 ();
 FILLCELL_X4 FILLER_18_278 ();
 FILLCELL_X1 FILLER_18_300 ();
 FILLCELL_X1 FILLER_18_304 ();
 FILLCELL_X1 FILLER_18_314 ();
 FILLCELL_X2 FILLER_18_324 ();
 FILLCELL_X2 FILLER_18_335 ();
 FILLCELL_X2 FILLER_18_354 ();
 FILLCELL_X4 FILLER_18_363 ();
 FILLCELL_X1 FILLER_18_367 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X2 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_18 ();
 FILLCELL_X1 FILLER_19_36 ();
 FILLCELL_X2 FILLER_19_41 ();
 FILLCELL_X4 FILLER_19_50 ();
 FILLCELL_X1 FILLER_19_58 ();
 FILLCELL_X2 FILLER_19_63 ();
 FILLCELL_X1 FILLER_19_65 ();
 FILLCELL_X8 FILLER_19_74 ();
 FILLCELL_X2 FILLER_19_82 ();
 FILLCELL_X16 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_114 ();
 FILLCELL_X2 FILLER_19_147 ();
 FILLCELL_X1 FILLER_19_149 ();
 FILLCELL_X4 FILLER_19_159 ();
 FILLCELL_X1 FILLER_19_191 ();
 FILLCELL_X4 FILLER_19_209 ();
 FILLCELL_X2 FILLER_19_213 ();
 FILLCELL_X1 FILLER_19_218 ();
 FILLCELL_X4 FILLER_19_261 ();
 FILLCELL_X2 FILLER_19_282 ();
 FILLCELL_X1 FILLER_19_284 ();
 FILLCELL_X2 FILLER_19_333 ();
 FILLCELL_X16 FILLER_19_351 ();
 FILLCELL_X1 FILLER_19_367 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_3 ();
 FILLCELL_X1 FILLER_20_23 ();
 FILLCELL_X1 FILLER_20_65 ();
 FILLCELL_X1 FILLER_20_71 ();
 FILLCELL_X2 FILLER_20_75 ();
 FILLCELL_X1 FILLER_20_83 ();
 FILLCELL_X1 FILLER_20_89 ();
 FILLCELL_X1 FILLER_20_93 ();
 FILLCELL_X1 FILLER_20_97 ();
 FILLCELL_X4 FILLER_20_100 ();
 FILLCELL_X1 FILLER_20_104 ();
 FILLCELL_X4 FILLER_20_110 ();
 FILLCELL_X2 FILLER_20_128 ();
 FILLCELL_X8 FILLER_20_141 ();
 FILLCELL_X1 FILLER_20_149 ();
 FILLCELL_X4 FILLER_20_172 ();
 FILLCELL_X4 FILLER_20_181 ();
 FILLCELL_X8 FILLER_20_199 ();
 FILLCELL_X4 FILLER_20_207 ();
 FILLCELL_X1 FILLER_20_228 ();
 FILLCELL_X4 FILLER_20_239 ();
 FILLCELL_X2 FILLER_20_243 ();
 FILLCELL_X4 FILLER_20_249 ();
 FILLCELL_X1 FILLER_20_253 ();
 FILLCELL_X4 FILLER_20_279 ();
 FILLCELL_X2 FILLER_20_283 ();
 FILLCELL_X1 FILLER_20_285 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X1 FILLER_20_347 ();
 FILLCELL_X4 FILLER_20_351 ();
 FILLCELL_X2 FILLER_20_355 ();
 FILLCELL_X1 FILLER_20_357 ();
 FILLCELL_X4 FILLER_20_361 ();
 FILLCELL_X2 FILLER_20_365 ();
 FILLCELL_X1 FILLER_20_367 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_9 ();
 FILLCELL_X8 FILLER_21_32 ();
 FILLCELL_X4 FILLER_21_40 ();
 FILLCELL_X1 FILLER_21_44 ();
 FILLCELL_X4 FILLER_21_47 ();
 FILLCELL_X1 FILLER_21_51 ();
 FILLCELL_X1 FILLER_21_60 ();
 FILLCELL_X4 FILLER_21_113 ();
 FILLCELL_X8 FILLER_21_162 ();
 FILLCELL_X4 FILLER_21_170 ();
 FILLCELL_X2 FILLER_21_174 ();
 FILLCELL_X1 FILLER_21_176 ();
 FILLCELL_X16 FILLER_21_196 ();
 FILLCELL_X8 FILLER_21_212 ();
 FILLCELL_X2 FILLER_21_220 ();
 FILLCELL_X4 FILLER_21_234 ();
 FILLCELL_X1 FILLER_21_238 ();
 FILLCELL_X4 FILLER_21_253 ();
 FILLCELL_X4 FILLER_21_266 ();
 FILLCELL_X1 FILLER_21_270 ();
 FILLCELL_X1 FILLER_21_278 ();
 FILLCELL_X4 FILLER_21_302 ();
 FILLCELL_X2 FILLER_21_313 ();
 FILLCELL_X1 FILLER_21_315 ();
 FILLCELL_X4 FILLER_21_329 ();
 FILLCELL_X4 FILLER_21_363 ();
 FILLCELL_X1 FILLER_21_367 ();
 FILLCELL_X4 FILLER_22_1 ();
 FILLCELL_X1 FILLER_22_5 ();
 FILLCELL_X4 FILLER_22_26 ();
 FILLCELL_X2 FILLER_22_30 ();
 FILLCELL_X1 FILLER_22_32 ();
 FILLCELL_X1 FILLER_22_48 ();
 FILLCELL_X1 FILLER_22_57 ();
 FILLCELL_X4 FILLER_22_66 ();
 FILLCELL_X1 FILLER_22_72 ();
 FILLCELL_X2 FILLER_22_77 ();
 FILLCELL_X2 FILLER_22_93 ();
 FILLCELL_X1 FILLER_22_95 ();
 FILLCELL_X2 FILLER_22_105 ();
 FILLCELL_X1 FILLER_22_107 ();
 FILLCELL_X4 FILLER_22_119 ();
 FILLCELL_X8 FILLER_22_126 ();
 FILLCELL_X1 FILLER_22_134 ();
 FILLCELL_X8 FILLER_22_139 ();
 FILLCELL_X1 FILLER_22_174 ();
 FILLCELL_X1 FILLER_22_179 ();
 FILLCELL_X2 FILLER_22_193 ();
 FILLCELL_X1 FILLER_22_195 ();
 FILLCELL_X16 FILLER_22_206 ();
 FILLCELL_X2 FILLER_22_263 ();
 FILLCELL_X1 FILLER_22_265 ();
 FILLCELL_X2 FILLER_22_283 ();
 FILLCELL_X2 FILLER_22_292 ();
 FILLCELL_X4 FILLER_22_300 ();
 FILLCELL_X2 FILLER_22_304 ();
 FILLCELL_X2 FILLER_22_326 ();
 FILLCELL_X1 FILLER_22_328 ();
 FILLCELL_X8 FILLER_22_332 ();
 FILLCELL_X2 FILLER_22_340 ();
 FILLCELL_X8 FILLER_22_359 ();
 FILLCELL_X1 FILLER_22_367 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_9 ();
 FILLCELL_X4 FILLER_23_17 ();
 FILLCELL_X1 FILLER_23_21 ();
 FILLCELL_X4 FILLER_23_26 ();
 FILLCELL_X2 FILLER_23_30 ();
 FILLCELL_X1 FILLER_23_32 ();
 FILLCELL_X4 FILLER_23_38 ();
 FILLCELL_X2 FILLER_23_46 ();
 FILLCELL_X1 FILLER_23_55 ();
 FILLCELL_X4 FILLER_23_65 ();
 FILLCELL_X2 FILLER_23_69 ();
 FILLCELL_X8 FILLER_23_81 ();
 FILLCELL_X4 FILLER_23_89 ();
 FILLCELL_X1 FILLER_23_93 ();
 FILLCELL_X4 FILLER_23_97 ();
 FILLCELL_X1 FILLER_23_101 ();
 FILLCELL_X4 FILLER_23_123 ();
 FILLCELL_X1 FILLER_23_127 ();
 FILLCELL_X2 FILLER_23_133 ();
 FILLCELL_X8 FILLER_23_139 ();
 FILLCELL_X2 FILLER_23_147 ();
 FILLCELL_X1 FILLER_23_149 ();
 FILLCELL_X16 FILLER_23_154 ();
 FILLCELL_X4 FILLER_23_170 ();
 FILLCELL_X2 FILLER_23_184 ();
 FILLCELL_X2 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_195 ();
 FILLCELL_X2 FILLER_23_200 ();
 FILLCELL_X1 FILLER_23_202 ();
 FILLCELL_X4 FILLER_23_206 ();
 FILLCELL_X2 FILLER_23_210 ();
 FILLCELL_X4 FILLER_23_229 ();
 FILLCELL_X2 FILLER_23_233 ();
 FILLCELL_X32 FILLER_23_239 ();
 FILLCELL_X16 FILLER_23_271 ();
 FILLCELL_X4 FILLER_23_287 ();
 FILLCELL_X1 FILLER_23_291 ();
 FILLCELL_X1 FILLER_23_307 ();
 FILLCELL_X4 FILLER_23_311 ();
 FILLCELL_X2 FILLER_23_315 ();
 FILLCELL_X4 FILLER_23_346 ();
 FILLCELL_X2 FILLER_23_350 ();
 FILLCELL_X1 FILLER_23_352 ();
 FILLCELL_X2 FILLER_23_356 ();
 FILLCELL_X1 FILLER_23_358 ();
 FILLCELL_X2 FILLER_23_362 ();
 FILLCELL_X1 FILLER_23_364 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_9 ();
 FILLCELL_X1 FILLER_24_11 ();
 FILLCELL_X2 FILLER_24_15 ();
 FILLCELL_X1 FILLER_24_20 ();
 FILLCELL_X1 FILLER_24_32 ();
 FILLCELL_X2 FILLER_24_41 ();
 FILLCELL_X1 FILLER_24_43 ();
 FILLCELL_X4 FILLER_24_52 ();
 FILLCELL_X2 FILLER_24_64 ();
 FILLCELL_X2 FILLER_24_88 ();
 FILLCELL_X2 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_99 ();
 FILLCELL_X2 FILLER_24_112 ();
 FILLCELL_X1 FILLER_24_124 ();
 FILLCELL_X2 FILLER_24_130 ();
 FILLCELL_X1 FILLER_24_132 ();
 FILLCELL_X2 FILLER_24_157 ();
 FILLCELL_X1 FILLER_24_159 ();
 FILLCELL_X4 FILLER_24_171 ();
 FILLCELL_X2 FILLER_24_175 ();
 FILLCELL_X1 FILLER_24_190 ();
 FILLCELL_X8 FILLER_24_199 ();
 FILLCELL_X4 FILLER_24_207 ();
 FILLCELL_X1 FILLER_24_211 ();
 FILLCELL_X8 FILLER_24_241 ();
 FILLCELL_X2 FILLER_24_249 ();
 FILLCELL_X8 FILLER_24_261 ();
 FILLCELL_X2 FILLER_24_269 ();
 FILLCELL_X4 FILLER_24_278 ();
 FILLCELL_X1 FILLER_24_282 ();
 FILLCELL_X1 FILLER_24_297 ();
 FILLCELL_X4 FILLER_24_305 ();
 FILLCELL_X2 FILLER_24_309 ();
 FILLCELL_X1 FILLER_24_315 ();
 FILLCELL_X1 FILLER_24_367 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_9 ();
 FILLCELL_X4 FILLER_25_17 ();
 FILLCELL_X1 FILLER_25_21 ();
 FILLCELL_X8 FILLER_25_25 ();
 FILLCELL_X1 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_38 ();
 FILLCELL_X1 FILLER_25_46 ();
 FILLCELL_X1 FILLER_25_50 ();
 FILLCELL_X1 FILLER_25_57 ();
 FILLCELL_X8 FILLER_25_62 ();
 FILLCELL_X4 FILLER_25_70 ();
 FILLCELL_X1 FILLER_25_78 ();
 FILLCELL_X4 FILLER_25_82 ();
 FILLCELL_X2 FILLER_25_98 ();
 FILLCELL_X1 FILLER_25_100 ();
 FILLCELL_X2 FILLER_25_114 ();
 FILLCELL_X1 FILLER_25_116 ();
 FILLCELL_X16 FILLER_25_130 ();
 FILLCELL_X2 FILLER_25_146 ();
 FILLCELL_X16 FILLER_25_169 ();
 FILLCELL_X4 FILLER_25_185 ();
 FILLCELL_X2 FILLER_25_196 ();
 FILLCELL_X16 FILLER_25_201 ();
 FILLCELL_X8 FILLER_25_217 ();
 FILLCELL_X1 FILLER_25_225 ();
 FILLCELL_X1 FILLER_25_233 ();
 FILLCELL_X4 FILLER_25_245 ();
 FILLCELL_X1 FILLER_25_256 ();
 FILLCELL_X2 FILLER_25_266 ();
 FILLCELL_X1 FILLER_25_320 ();
 FILLCELL_X4 FILLER_25_338 ();
 FILLCELL_X1 FILLER_25_342 ();
 FILLCELL_X8 FILLER_25_347 ();
 FILLCELL_X4 FILLER_25_355 ();
 FILLCELL_X2 FILLER_25_359 ();
 FILLCELL_X1 FILLER_25_361 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_17 ();
 FILLCELL_X1 FILLER_26_19 ();
 FILLCELL_X2 FILLER_26_70 ();
 FILLCELL_X1 FILLER_26_72 ();
 FILLCELL_X1 FILLER_26_95 ();
 FILLCELL_X2 FILLER_26_107 ();
 FILLCELL_X1 FILLER_26_109 ();
 FILLCELL_X2 FILLER_26_119 ();
 FILLCELL_X4 FILLER_26_125 ();
 FILLCELL_X8 FILLER_26_134 ();
 FILLCELL_X4 FILLER_26_142 ();
 FILLCELL_X2 FILLER_26_146 ();
 FILLCELL_X1 FILLER_26_148 ();
 FILLCELL_X4 FILLER_26_165 ();
 FILLCELL_X2 FILLER_26_169 ();
 FILLCELL_X1 FILLER_26_171 ();
 FILLCELL_X1 FILLER_26_181 ();
 FILLCELL_X2 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_195 ();
 FILLCELL_X16 FILLER_26_199 ();
 FILLCELL_X8 FILLER_26_215 ();
 FILLCELL_X4 FILLER_26_223 ();
 FILLCELL_X1 FILLER_26_227 ();
 FILLCELL_X8 FILLER_26_245 ();
 FILLCELL_X2 FILLER_26_253 ();
 FILLCELL_X8 FILLER_26_261 ();
 FILLCELL_X2 FILLER_26_269 ();
 FILLCELL_X4 FILLER_26_278 ();
 FILLCELL_X8 FILLER_26_289 ();
 FILLCELL_X1 FILLER_26_297 ();
 FILLCELL_X8 FILLER_26_307 ();
 FILLCELL_X2 FILLER_26_315 ();
 FILLCELL_X8 FILLER_26_328 ();
 FILLCELL_X2 FILLER_26_353 ();
 FILLCELL_X1 FILLER_26_361 ();
 FILLCELL_X2 FILLER_26_365 ();
 FILLCELL_X1 FILLER_26_367 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X1 FILLER_27_3 ();
 FILLCELL_X16 FILLER_27_7 ();
 FILLCELL_X4 FILLER_27_23 ();
 FILLCELL_X1 FILLER_27_27 ();
 FILLCELL_X8 FILLER_27_50 ();
 FILLCELL_X1 FILLER_27_62 ();
 FILLCELL_X1 FILLER_27_67 ();
 FILLCELL_X1 FILLER_27_72 ();
 FILLCELL_X1 FILLER_27_77 ();
 FILLCELL_X1 FILLER_27_98 ();
 FILLCELL_X8 FILLER_27_129 ();
 FILLCELL_X2 FILLER_27_137 ();
 FILLCELL_X2 FILLER_27_164 ();
 FILLCELL_X1 FILLER_27_166 ();
 FILLCELL_X32 FILLER_27_188 ();
 FILLCELL_X4 FILLER_27_220 ();
 FILLCELL_X1 FILLER_27_224 ();
 FILLCELL_X2 FILLER_27_237 ();
 FILLCELL_X4 FILLER_27_246 ();
 FILLCELL_X1 FILLER_27_250 ();
 FILLCELL_X1 FILLER_27_282 ();
 FILLCELL_X8 FILLER_27_300 ();
 FILLCELL_X4 FILLER_27_308 ();
 FILLCELL_X1 FILLER_27_312 ();
 FILLCELL_X8 FILLER_27_345 ();
 FILLCELL_X2 FILLER_27_360 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_5 ();
 FILLCELL_X1 FILLER_28_47 ();
 FILLCELL_X2 FILLER_28_73 ();
 FILLCELL_X1 FILLER_28_75 ();
 FILLCELL_X4 FILLER_28_80 ();
 FILLCELL_X2 FILLER_28_84 ();
 FILLCELL_X8 FILLER_28_96 ();
 FILLCELL_X4 FILLER_28_104 ();
 FILLCELL_X1 FILLER_28_108 ();
 FILLCELL_X8 FILLER_28_129 ();
 FILLCELL_X4 FILLER_28_137 ();
 FILLCELL_X2 FILLER_28_141 ();
 FILLCELL_X1 FILLER_28_143 ();
 FILLCELL_X1 FILLER_28_156 ();
 FILLCELL_X4 FILLER_28_163 ();
 FILLCELL_X2 FILLER_28_167 ();
 FILLCELL_X2 FILLER_28_176 ();
 FILLCELL_X1 FILLER_28_185 ();
 FILLCELL_X2 FILLER_28_200 ();
 FILLCELL_X1 FILLER_28_202 ();
 FILLCELL_X1 FILLER_28_234 ();
 FILLCELL_X8 FILLER_28_269 ();
 FILLCELL_X2 FILLER_28_277 ();
 FILLCELL_X1 FILLER_28_279 ();
 FILLCELL_X4 FILLER_28_287 ();
 FILLCELL_X1 FILLER_28_291 ();
 FILLCELL_X4 FILLER_28_301 ();
 FILLCELL_X2 FILLER_28_305 ();
 FILLCELL_X1 FILLER_28_307 ();
 FILLCELL_X4 FILLER_28_322 ();
 FILLCELL_X2 FILLER_28_326 ();
 FILLCELL_X8 FILLER_28_335 ();
 FILLCELL_X2 FILLER_28_343 ();
 FILLCELL_X2 FILLER_28_365 ();
 FILLCELL_X1 FILLER_28_367 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X2 FILLER_29_5 ();
 FILLCELL_X2 FILLER_29_10 ();
 FILLCELL_X1 FILLER_29_26 ();
 FILLCELL_X4 FILLER_29_43 ();
 FILLCELL_X2 FILLER_29_47 ();
 FILLCELL_X4 FILLER_29_54 ();
 FILLCELL_X2 FILLER_29_58 ();
 FILLCELL_X4 FILLER_29_74 ();
 FILLCELL_X4 FILLER_29_84 ();
 FILLCELL_X4 FILLER_29_94 ();
 FILLCELL_X4 FILLER_29_107 ();
 FILLCELL_X2 FILLER_29_111 ();
 FILLCELL_X2 FILLER_29_139 ();
 FILLCELL_X1 FILLER_29_141 ();
 FILLCELL_X1 FILLER_29_163 ();
 FILLCELL_X16 FILLER_29_171 ();
 FILLCELL_X8 FILLER_29_187 ();
 FILLCELL_X4 FILLER_29_195 ();
 FILLCELL_X4 FILLER_29_216 ();
 FILLCELL_X2 FILLER_29_220 ();
 FILLCELL_X2 FILLER_29_236 ();
 FILLCELL_X1 FILLER_29_238 ();
 FILLCELL_X4 FILLER_29_246 ();
 FILLCELL_X2 FILLER_29_250 ();
 FILLCELL_X1 FILLER_29_252 ();
 FILLCELL_X16 FILLER_29_260 ();
 FILLCELL_X8 FILLER_29_276 ();
 FILLCELL_X2 FILLER_29_284 ();
 FILLCELL_X1 FILLER_29_286 ();
 FILLCELL_X8 FILLER_29_291 ();
 FILLCELL_X1 FILLER_29_304 ();
 FILLCELL_X4 FILLER_29_322 ();
 FILLCELL_X1 FILLER_29_326 ();
 FILLCELL_X4 FILLER_29_344 ();
 FILLCELL_X1 FILLER_29_348 ();
 FILLCELL_X4 FILLER_29_356 ();
 FILLCELL_X2 FILLER_29_363 ();
 FILLCELL_X2 FILLER_30_4 ();
 FILLCELL_X1 FILLER_30_6 ();
 FILLCELL_X8 FILLER_30_10 ();
 FILLCELL_X2 FILLER_30_18 ();
 FILLCELL_X1 FILLER_30_20 ();
 FILLCELL_X1 FILLER_30_31 ();
 FILLCELL_X2 FILLER_30_37 ();
 FILLCELL_X2 FILLER_30_43 ();
 FILLCELL_X1 FILLER_30_58 ();
 FILLCELL_X2 FILLER_30_65 ();
 FILLCELL_X2 FILLER_30_71 ();
 FILLCELL_X2 FILLER_30_77 ();
 FILLCELL_X1 FILLER_30_106 ();
 FILLCELL_X2 FILLER_30_111 ();
 FILLCELL_X8 FILLER_30_136 ();
 FILLCELL_X2 FILLER_30_144 ();
 FILLCELL_X1 FILLER_30_146 ();
 FILLCELL_X2 FILLER_30_152 ();
 FILLCELL_X1 FILLER_30_154 ();
 FILLCELL_X1 FILLER_30_163 ();
 FILLCELL_X8 FILLER_30_166 ();
 FILLCELL_X1 FILLER_30_174 ();
 FILLCELL_X4 FILLER_30_192 ();
 FILLCELL_X1 FILLER_30_196 ();
 FILLCELL_X1 FILLER_30_221 ();
 FILLCELL_X2 FILLER_30_229 ();
 FILLCELL_X1 FILLER_30_231 ();
 FILLCELL_X8 FILLER_30_247 ();
 FILLCELL_X2 FILLER_30_255 ();
 FILLCELL_X1 FILLER_30_257 ();
 FILLCELL_X2 FILLER_30_266 ();
 FILLCELL_X4 FILLER_30_270 ();
 FILLCELL_X2 FILLER_30_284 ();
 FILLCELL_X1 FILLER_30_286 ();
 FILLCELL_X1 FILLER_30_291 ();
 FILLCELL_X1 FILLER_30_301 ();
 FILLCELL_X4 FILLER_30_323 ();
 FILLCELL_X2 FILLER_30_327 ();
 FILLCELL_X8 FILLER_30_336 ();
 FILLCELL_X2 FILLER_30_344 ();
 FILLCELL_X2 FILLER_30_366 ();
 FILLCELL_X2 FILLER_31_10 ();
 FILLCELL_X4 FILLER_31_36 ();
 FILLCELL_X2 FILLER_31_52 ();
 FILLCELL_X4 FILLER_31_92 ();
 FILLCELL_X1 FILLER_31_96 ();
 FILLCELL_X8 FILLER_31_101 ();
 FILLCELL_X1 FILLER_31_109 ();
 FILLCELL_X8 FILLER_31_119 ();
 FILLCELL_X1 FILLER_31_127 ();
 FILLCELL_X8 FILLER_31_133 ();
 FILLCELL_X4 FILLER_31_141 ();
 FILLCELL_X2 FILLER_31_145 ();
 FILLCELL_X1 FILLER_31_164 ();
 FILLCELL_X4 FILLER_31_199 ();
 FILLCELL_X2 FILLER_31_203 ();
 FILLCELL_X1 FILLER_31_256 ();
 FILLCELL_X1 FILLER_31_293 ();
 FILLCELL_X8 FILLER_31_318 ();
 FILLCELL_X2 FILLER_31_326 ();
 FILLCELL_X8 FILLER_31_335 ();
 FILLCELL_X8 FILLER_31_353 ();
 FILLCELL_X1 FILLER_31_361 ();
 FILLCELL_X2 FILLER_31_365 ();
 FILLCELL_X1 FILLER_31_367 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_3 ();
 FILLCELL_X16 FILLER_32_7 ();
 FILLCELL_X1 FILLER_32_23 ();
 FILLCELL_X2 FILLER_32_35 ();
 FILLCELL_X2 FILLER_32_43 ();
 FILLCELL_X1 FILLER_32_45 ();
 FILLCELL_X1 FILLER_32_49 ();
 FILLCELL_X2 FILLER_32_52 ();
 FILLCELL_X1 FILLER_32_54 ();
 FILLCELL_X2 FILLER_32_69 ();
 FILLCELL_X1 FILLER_32_71 ();
 FILLCELL_X8 FILLER_32_86 ();
 FILLCELL_X2 FILLER_32_94 ();
 FILLCELL_X1 FILLER_32_96 ();
 FILLCELL_X2 FILLER_32_102 ();
 FILLCELL_X2 FILLER_32_110 ();
 FILLCELL_X2 FILLER_32_121 ();
 FILLCELL_X1 FILLER_32_123 ();
 FILLCELL_X4 FILLER_32_141 ();
 FILLCELL_X32 FILLER_32_181 ();
 FILLCELL_X16 FILLER_32_213 ();
 FILLCELL_X2 FILLER_32_229 ();
 FILLCELL_X1 FILLER_32_231 ();
 FILLCELL_X8 FILLER_32_256 ();
 FILLCELL_X2 FILLER_32_264 ();
 FILLCELL_X1 FILLER_32_266 ();
 FILLCELL_X4 FILLER_32_271 ();
 FILLCELL_X1 FILLER_32_275 ();
 FILLCELL_X4 FILLER_32_283 ();
 FILLCELL_X1 FILLER_32_287 ();
 FILLCELL_X2 FILLER_32_291 ();
 FILLCELL_X4 FILLER_32_304 ();
 FILLCELL_X1 FILLER_32_308 ();
 FILLCELL_X2 FILLER_32_363 ();
 FILLCELL_X1 FILLER_33_4 ();
 FILLCELL_X1 FILLER_33_12 ();
 FILLCELL_X1 FILLER_33_16 ();
 FILLCELL_X4 FILLER_33_63 ();
 FILLCELL_X1 FILLER_33_67 ();
 FILLCELL_X16 FILLER_33_72 ();
 FILLCELL_X8 FILLER_33_88 ();
 FILLCELL_X1 FILLER_33_96 ();
 FILLCELL_X2 FILLER_33_102 ();
 FILLCELL_X1 FILLER_33_104 ();
 FILLCELL_X16 FILLER_33_114 ();
 FILLCELL_X8 FILLER_33_130 ();
 FILLCELL_X8 FILLER_33_151 ();
 FILLCELL_X4 FILLER_33_159 ();
 FILLCELL_X2 FILLER_33_163 ();
 FILLCELL_X1 FILLER_33_165 ();
 FILLCELL_X2 FILLER_33_183 ();
 FILLCELL_X1 FILLER_33_185 ();
 FILLCELL_X32 FILLER_33_203 ();
 FILLCELL_X4 FILLER_33_235 ();
 FILLCELL_X2 FILLER_33_239 ();
 FILLCELL_X4 FILLER_33_248 ();
 FILLCELL_X1 FILLER_33_252 ();
 FILLCELL_X2 FILLER_33_260 ();
 FILLCELL_X1 FILLER_33_262 ();
 FILLCELL_X2 FILLER_33_270 ();
 FILLCELL_X1 FILLER_33_272 ();
 FILLCELL_X2 FILLER_33_290 ();
 FILLCELL_X1 FILLER_33_292 ();
 FILLCELL_X8 FILLER_33_300 ();
 FILLCELL_X2 FILLER_33_308 ();
 FILLCELL_X32 FILLER_33_317 ();
 FILLCELL_X4 FILLER_33_349 ();
 FILLCELL_X2 FILLER_33_363 ();
 FILLCELL_X2 FILLER_34_4 ();
 FILLCELL_X2 FILLER_34_23 ();
 FILLCELL_X1 FILLER_34_25 ();
 FILLCELL_X8 FILLER_34_29 ();
 FILLCELL_X2 FILLER_34_37 ();
 FILLCELL_X2 FILLER_34_61 ();
 FILLCELL_X1 FILLER_34_63 ();
 FILLCELL_X8 FILLER_34_69 ();
 FILLCELL_X2 FILLER_34_77 ();
 FILLCELL_X16 FILLER_34_111 ();
 FILLCELL_X8 FILLER_34_127 ();
 FILLCELL_X4 FILLER_34_142 ();
 FILLCELL_X1 FILLER_34_146 ();
 FILLCELL_X4 FILLER_34_167 ();
 FILLCELL_X16 FILLER_34_178 ();
 FILLCELL_X2 FILLER_34_194 ();
 FILLCELL_X8 FILLER_34_200 ();
 FILLCELL_X4 FILLER_34_208 ();
 FILLCELL_X2 FILLER_34_212 ();
 FILLCELL_X2 FILLER_34_221 ();
 FILLCELL_X1 FILLER_34_223 ();
 FILLCELL_X16 FILLER_34_231 ();
 FILLCELL_X4 FILLER_34_247 ();
 FILLCELL_X2 FILLER_34_251 ();
 FILLCELL_X16 FILLER_34_270 ();
 FILLCELL_X2 FILLER_34_286 ();
 FILLCELL_X1 FILLER_34_288 ();
 FILLCELL_X4 FILLER_34_306 ();
 FILLCELL_X8 FILLER_34_317 ();
 FILLCELL_X4 FILLER_34_325 ();
 FILLCELL_X4 FILLER_34_343 ();
 FILLCELL_X2 FILLER_34_347 ();
 FILLCELL_X1 FILLER_34_352 ();
 FILLCELL_X2 FILLER_34_366 ();
 FILLCELL_X2 FILLER_35_1 ();
 FILLCELL_X4 FILLER_35_9 ();
 FILLCELL_X1 FILLER_35_13 ();
 FILLCELL_X4 FILLER_35_21 ();
 FILLCELL_X2 FILLER_35_25 ();
 FILLCELL_X1 FILLER_35_52 ();
 FILLCELL_X8 FILLER_35_56 ();
 FILLCELL_X2 FILLER_35_64 ();
 FILLCELL_X4 FILLER_35_69 ();
 FILLCELL_X2 FILLER_35_73 ();
 FILLCELL_X1 FILLER_35_75 ();
 FILLCELL_X4 FILLER_35_93 ();
 FILLCELL_X8 FILLER_35_120 ();
 FILLCELL_X4 FILLER_35_128 ();
 FILLCELL_X4 FILLER_35_149 ();
 FILLCELL_X1 FILLER_35_153 ();
 FILLCELL_X2 FILLER_35_159 ();
 FILLCELL_X1 FILLER_35_161 ();
 FILLCELL_X16 FILLER_35_171 ();
 FILLCELL_X8 FILLER_35_187 ();
 FILLCELL_X4 FILLER_35_195 ();
 FILLCELL_X2 FILLER_35_199 ();
 FILLCELL_X1 FILLER_35_201 ();
 FILLCELL_X8 FILLER_35_219 ();
 FILLCELL_X4 FILLER_35_234 ();
 FILLCELL_X2 FILLER_35_245 ();
 FILLCELL_X16 FILLER_35_254 ();
 FILLCELL_X2 FILLER_35_270 ();
 FILLCELL_X1 FILLER_35_272 ();
 FILLCELL_X1 FILLER_35_280 ();
 FILLCELL_X2 FILLER_35_288 ();
 FILLCELL_X8 FILLER_35_297 ();
 FILLCELL_X4 FILLER_35_305 ();
 FILLCELL_X2 FILLER_35_309 ();
 FILLCELL_X2 FILLER_35_345 ();
 FILLCELL_X1 FILLER_35_364 ();
 FILLCELL_X2 FILLER_36_4 ();
 FILLCELL_X16 FILLER_36_54 ();
 FILLCELL_X4 FILLER_36_70 ();
 FILLCELL_X2 FILLER_36_74 ();
 FILLCELL_X1 FILLER_36_76 ();
 FILLCELL_X1 FILLER_36_83 ();
 FILLCELL_X2 FILLER_36_89 ();
 FILLCELL_X4 FILLER_36_118 ();
 FILLCELL_X2 FILLER_36_122 ();
 FILLCELL_X1 FILLER_36_124 ();
 FILLCELL_X4 FILLER_36_129 ();
 FILLCELL_X2 FILLER_36_133 ();
 FILLCELL_X1 FILLER_36_135 ();
 FILLCELL_X4 FILLER_36_144 ();
 FILLCELL_X2 FILLER_36_148 ();
 FILLCELL_X1 FILLER_36_150 ();
 FILLCELL_X16 FILLER_36_189 ();
 FILLCELL_X8 FILLER_36_205 ();
 FILLCELL_X4 FILLER_36_213 ();
 FILLCELL_X4 FILLER_36_251 ();
 FILLCELL_X2 FILLER_36_255 ();
 FILLCELL_X1 FILLER_36_257 ();
 FILLCELL_X2 FILLER_36_265 ();
 FILLCELL_X1 FILLER_36_267 ();
 FILLCELL_X2 FILLER_36_285 ();
 FILLCELL_X1 FILLER_36_287 ();
 FILLCELL_X4 FILLER_36_305 ();
 FILLCELL_X1 FILLER_36_309 ();
 FILLCELL_X8 FILLER_36_317 ();
 FILLCELL_X4 FILLER_36_325 ();
 FILLCELL_X8 FILLER_36_336 ();
 FILLCELL_X2 FILLER_36_351 ();
 FILLCELL_X1 FILLER_36_353 ();
 FILLCELL_X2 FILLER_36_366 ();
 FILLCELL_X1 FILLER_37_7 ();
 FILLCELL_X32 FILLER_37_28 ();
 FILLCELL_X4 FILLER_37_60 ();
 FILLCELL_X1 FILLER_37_64 ();
 FILLCELL_X8 FILLER_37_85 ();
 FILLCELL_X2 FILLER_37_93 ();
 FILLCELL_X1 FILLER_37_95 ();
 FILLCELL_X1 FILLER_37_102 ();
 FILLCELL_X16 FILLER_37_110 ();
 FILLCELL_X4 FILLER_37_126 ();
 FILLCELL_X1 FILLER_37_130 ();
 FILLCELL_X4 FILLER_37_135 ();
 FILLCELL_X4 FILLER_37_149 ();
 FILLCELL_X2 FILLER_37_160 ();
 FILLCELL_X1 FILLER_37_162 ();
 FILLCELL_X32 FILLER_37_168 ();
 FILLCELL_X32 FILLER_37_200 ();
 FILLCELL_X4 FILLER_37_232 ();
 FILLCELL_X1 FILLER_37_236 ();
 FILLCELL_X8 FILLER_37_244 ();
 FILLCELL_X1 FILLER_37_252 ();
 FILLCELL_X4 FILLER_37_270 ();
 FILLCELL_X1 FILLER_37_274 ();
 FILLCELL_X8 FILLER_37_299 ();
 FILLCELL_X1 FILLER_37_307 ();
 FILLCELL_X1 FILLER_38_14 ();
 FILLCELL_X16 FILLER_38_25 ();
 FILLCELL_X8 FILLER_38_41 ();
 FILLCELL_X4 FILLER_38_49 ();
 FILLCELL_X8 FILLER_38_58 ();
 FILLCELL_X4 FILLER_38_66 ();
 FILLCELL_X2 FILLER_38_70 ();
 FILLCELL_X1 FILLER_38_72 ();
 FILLCELL_X8 FILLER_38_110 ();
 FILLCELL_X1 FILLER_38_118 ();
 FILLCELL_X1 FILLER_38_122 ();
 FILLCELL_X1 FILLER_38_142 ();
 FILLCELL_X2 FILLER_38_153 ();
 FILLCELL_X1 FILLER_38_155 ();
 FILLCELL_X32 FILLER_38_167 ();
 FILLCELL_X32 FILLER_38_199 ();
 FILLCELL_X2 FILLER_38_231 ();
 FILLCELL_X1 FILLER_38_233 ();
 FILLCELL_X32 FILLER_38_272 ();
 FILLCELL_X8 FILLER_38_304 ();
 FILLCELL_X4 FILLER_38_312 ();
 FILLCELL_X2 FILLER_38_323 ();
 FILLCELL_X2 FILLER_39_1 ();
 FILLCELL_X1 FILLER_39_3 ();
 FILLCELL_X8 FILLER_39_38 ();
 FILLCELL_X2 FILLER_39_46 ();
 FILLCELL_X1 FILLER_39_48 ();
 FILLCELL_X8 FILLER_39_52 ();
 FILLCELL_X1 FILLER_39_60 ();
 FILLCELL_X4 FILLER_39_84 ();
 FILLCELL_X4 FILLER_39_94 ();
 FILLCELL_X2 FILLER_39_98 ();
 FILLCELL_X1 FILLER_39_100 ();
 FILLCELL_X16 FILLER_39_116 ();
 FILLCELL_X2 FILLER_39_132 ();
 FILLCELL_X1 FILLER_39_141 ();
 FILLCELL_X4 FILLER_39_149 ();
 FILLCELL_X2 FILLER_39_160 ();
 FILLCELL_X16 FILLER_39_179 ();
 FILLCELL_X8 FILLER_39_195 ();
 FILLCELL_X1 FILLER_39_203 ();
 FILLCELL_X32 FILLER_39_207 ();
 FILLCELL_X32 FILLER_39_239 ();
 FILLCELL_X4 FILLER_39_271 ();
 FILLCELL_X1 FILLER_39_302 ();
 FILLCELL_X16 FILLER_39_310 ();
 FILLCELL_X4 FILLER_39_326 ();
 FILLCELL_X1 FILLER_39_330 ();
 FILLCELL_X4 FILLER_39_341 ();
 FILLCELL_X2 FILLER_39_345 ();
 FILLCELL_X2 FILLER_39_350 ();
 FILLCELL_X1 FILLER_39_352 ();
 FILLCELL_X4 FILLER_39_363 ();
 FILLCELL_X1 FILLER_39_367 ();
 FILLCELL_X2 FILLER_40_32 ();
 FILLCELL_X1 FILLER_40_34 ();
 FILLCELL_X2 FILLER_40_65 ();
 FILLCELL_X2 FILLER_40_84 ();
 FILLCELL_X32 FILLER_40_120 ();
 FILLCELL_X32 FILLER_40_152 ();
 FILLCELL_X32 FILLER_40_184 ();
 FILLCELL_X32 FILLER_40_216 ();
 FILLCELL_X32 FILLER_40_248 ();
 FILLCELL_X8 FILLER_40_280 ();
 FILLCELL_X4 FILLER_40_288 ();
 FILLCELL_X2 FILLER_40_297 ();
 FILLCELL_X8 FILLER_40_319 ();
 FILLCELL_X2 FILLER_40_327 ();
 FILLCELL_X2 FILLER_40_332 ();
 FILLCELL_X1 FILLER_40_361 ();
 FILLCELL_X2 FILLER_41_8 ();
 FILLCELL_X2 FILLER_41_13 ();
 FILLCELL_X1 FILLER_41_15 ();
 FILLCELL_X2 FILLER_41_19 ();
 FILLCELL_X1 FILLER_41_21 ();
 FILLCELL_X16 FILLER_41_53 ();
 FILLCELL_X4 FILLER_41_69 ();
 FILLCELL_X2 FILLER_41_73 ();
 FILLCELL_X1 FILLER_41_75 ();
 FILLCELL_X4 FILLER_41_82 ();
 FILLCELL_X2 FILLER_41_86 ();
 FILLCELL_X1 FILLER_41_88 ();
 FILLCELL_X8 FILLER_41_92 ();
 FILLCELL_X4 FILLER_41_100 ();
 FILLCELL_X2 FILLER_41_104 ();
 FILLCELL_X1 FILLER_41_106 ();
 FILLCELL_X32 FILLER_41_110 ();
 FILLCELL_X32 FILLER_41_142 ();
 FILLCELL_X32 FILLER_41_174 ();
 FILLCELL_X16 FILLER_41_206 ();
 FILLCELL_X8 FILLER_41_222 ();
 FILLCELL_X4 FILLER_41_230 ();
 FILLCELL_X2 FILLER_41_234 ();
 FILLCELL_X8 FILLER_41_243 ();
 FILLCELL_X1 FILLER_41_251 ();
 FILLCELL_X4 FILLER_41_259 ();
 FILLCELL_X16 FILLER_41_270 ();
 FILLCELL_X4 FILLER_41_286 ();
 FILLCELL_X1 FILLER_41_290 ();
 FILLCELL_X32 FILLER_41_298 ();
 FILLCELL_X2 FILLER_41_330 ();
 FILLCELL_X1 FILLER_41_332 ();
 FILLCELL_X8 FILLER_41_339 ();
 FILLCELL_X2 FILLER_41_347 ();
 FILLCELL_X1 FILLER_41_349 ();
 FILLCELL_X1 FILLER_41_367 ();
 FILLCELL_X2 FILLER_42_1 ();
 FILLCELL_X2 FILLER_42_20 ();
 FILLCELL_X2 FILLER_42_25 ();
 FILLCELL_X1 FILLER_42_27 ();
 FILLCELL_X4 FILLER_42_48 ();
 FILLCELL_X2 FILLER_42_52 ();
 FILLCELL_X16 FILLER_42_59 ();
 FILLCELL_X1 FILLER_42_75 ();
 FILLCELL_X4 FILLER_42_83 ();
 FILLCELL_X2 FILLER_42_87 ();
 FILLCELL_X1 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_101 ();
 FILLCELL_X16 FILLER_42_133 ();
 FILLCELL_X8 FILLER_42_149 ();
 FILLCELL_X32 FILLER_42_162 ();
 FILLCELL_X16 FILLER_42_194 ();
 FILLCELL_X2 FILLER_42_210 ();
 FILLCELL_X8 FILLER_42_217 ();
 FILLCELL_X4 FILLER_42_225 ();
 FILLCELL_X1 FILLER_42_229 ();
 FILLCELL_X4 FILLER_42_281 ();
 FILLCELL_X2 FILLER_42_288 ();
 FILLCELL_X1 FILLER_42_314 ();
 FILLCELL_X8 FILLER_42_337 ();
 FILLCELL_X4 FILLER_42_345 ();
 FILLCELL_X2 FILLER_42_356 ();
 FILLCELL_X1 FILLER_42_358 ();
 FILLCELL_X2 FILLER_42_362 ();
 FILLCELL_X1 FILLER_42_364 ();
 FILLCELL_X2 FILLER_43_7 ();
 FILLCELL_X1 FILLER_43_9 ();
 FILLCELL_X1 FILLER_43_16 ();
 FILLCELL_X32 FILLER_43_41 ();
 FILLCELL_X1 FILLER_43_73 ();
 FILLCELL_X32 FILLER_43_91 ();
 FILLCELL_X32 FILLER_43_123 ();
 FILLCELL_X32 FILLER_43_155 ();
 FILLCELL_X8 FILLER_43_187 ();
 FILLCELL_X2 FILLER_43_195 ();
 FILLCELL_X8 FILLER_43_204 ();
 FILLCELL_X8 FILLER_43_236 ();
 FILLCELL_X4 FILLER_43_244 ();
 FILLCELL_X2 FILLER_43_248 ();
 FILLCELL_X1 FILLER_43_250 ();
 FILLCELL_X4 FILLER_43_254 ();
 FILLCELL_X1 FILLER_43_258 ();
 FILLCELL_X8 FILLER_43_262 ();
 FILLCELL_X4 FILLER_43_270 ();
 FILLCELL_X1 FILLER_43_274 ();
 FILLCELL_X1 FILLER_43_299 ();
 FILLCELL_X1 FILLER_43_317 ();
 FILLCELL_X4 FILLER_43_325 ();
 FILLCELL_X1 FILLER_43_329 ();
 FILLCELL_X4 FILLER_43_340 ();
 FILLCELL_X1 FILLER_43_344 ();
 FILLCELL_X16 FILLER_44_53 ();
 FILLCELL_X8 FILLER_44_69 ();
 FILLCELL_X32 FILLER_44_84 ();
 FILLCELL_X32 FILLER_44_116 ();
 FILLCELL_X32 FILLER_44_148 ();
 FILLCELL_X8 FILLER_44_180 ();
 FILLCELL_X4 FILLER_44_188 ();
 FILLCELL_X4 FILLER_44_209 ();
 FILLCELL_X2 FILLER_44_213 ();
 FILLCELL_X1 FILLER_44_215 ();
 FILLCELL_X8 FILLER_44_223 ();
 FILLCELL_X2 FILLER_44_231 ();
 FILLCELL_X8 FILLER_44_240 ();
 FILLCELL_X8 FILLER_44_255 ();
 FILLCELL_X4 FILLER_44_263 ();
 FILLCELL_X8 FILLER_44_274 ();
 FILLCELL_X2 FILLER_44_282 ();
 FILLCELL_X16 FILLER_44_301 ();
 FILLCELL_X2 FILLER_44_317 ();
 FILLCELL_X2 FILLER_44_325 ();
 FILLCELL_X1 FILLER_44_327 ();
 FILLCELL_X2 FILLER_44_345 ();
 FILLCELL_X4 FILLER_44_356 ();
 FILLCELL_X2 FILLER_44_360 ();
 FILLCELL_X4 FILLER_45_38 ();
 FILLCELL_X1 FILLER_45_42 ();
 FILLCELL_X4 FILLER_45_94 ();
 FILLCELL_X2 FILLER_45_98 ();
 FILLCELL_X16 FILLER_45_103 ();
 FILLCELL_X8 FILLER_45_119 ();
 FILLCELL_X32 FILLER_45_130 ();
 FILLCELL_X8 FILLER_45_162 ();
 FILLCELL_X2 FILLER_45_170 ();
 FILLCELL_X8 FILLER_45_199 ();
 FILLCELL_X2 FILLER_45_207 ();
 FILLCELL_X1 FILLER_45_209 ();
 FILLCELL_X2 FILLER_45_227 ();
 FILLCELL_X2 FILLER_45_263 ();
 FILLCELL_X8 FILLER_45_282 ();
 FILLCELL_X1 FILLER_45_290 ();
 FILLCELL_X2 FILLER_45_298 ();
 FILLCELL_X1 FILLER_45_320 ();
 FILLCELL_X1 FILLER_45_324 ();
 FILLCELL_X1 FILLER_45_332 ();
 FILLCELL_X1 FILLER_45_336 ();
 FILLCELL_X2 FILLER_45_363 ();
 FILLCELL_X16 FILLER_46_63 ();
 FILLCELL_X4 FILLER_46_79 ();
 FILLCELL_X2 FILLER_46_83 ();
 FILLCELL_X8 FILLER_46_92 ();
 FILLCELL_X4 FILLER_46_100 ();
 FILLCELL_X8 FILLER_46_117 ();
 FILLCELL_X16 FILLER_46_132 ();
 FILLCELL_X2 FILLER_46_148 ();
 FILLCELL_X1 FILLER_46_150 ();
 FILLCELL_X4 FILLER_46_158 ();
 FILLCELL_X4 FILLER_46_165 ();
 FILLCELL_X1 FILLER_46_169 ();
 FILLCELL_X8 FILLER_46_177 ();
 FILLCELL_X4 FILLER_46_185 ();
 FILLCELL_X2 FILLER_46_189 ();
 FILLCELL_X1 FILLER_46_198 ();
 FILLCELL_X1 FILLER_46_205 ();
 FILLCELL_X2 FILLER_46_213 ();
 FILLCELL_X1 FILLER_46_215 ();
 FILLCELL_X8 FILLER_46_219 ();
 FILLCELL_X4 FILLER_46_240 ();
 FILLCELL_X1 FILLER_46_244 ();
 FILLCELL_X8 FILLER_46_251 ();
 FILLCELL_X1 FILLER_46_259 ();
 FILLCELL_X4 FILLER_46_270 ();
 FILLCELL_X2 FILLER_46_274 ();
 FILLCELL_X1 FILLER_46_276 ();
 FILLCELL_X2 FILLER_46_301 ();
 FILLCELL_X1 FILLER_46_303 ();
 FILLCELL_X4 FILLER_46_311 ();
 FILLCELL_X1 FILLER_46_315 ();
 FILLCELL_X4 FILLER_46_319 ();
 FILLCELL_X1 FILLER_46_323 ();
 FILLCELL_X1 FILLER_46_344 ();
 FILLCELL_X1 FILLER_46_367 ();
 FILLCELL_X1 FILLER_47_10 ();
 FILLCELL_X1 FILLER_47_26 ();
 FILLCELL_X1 FILLER_47_41 ();
 FILLCELL_X1 FILLER_47_49 ();
 FILLCELL_X1 FILLER_47_55 ();
 FILLCELL_X1 FILLER_47_59 ();
 FILLCELL_X4 FILLER_47_62 ();
 FILLCELL_X2 FILLER_47_71 ();
 FILLCELL_X2 FILLER_47_75 ();
 FILLCELL_X2 FILLER_47_100 ();
 FILLCELL_X1 FILLER_47_102 ();
 FILLCELL_X1 FILLER_47_146 ();
 FILLCELL_X2 FILLER_47_184 ();
 FILLCELL_X4 FILLER_47_220 ();
 FILLCELL_X1 FILLER_47_224 ();
 FILLCELL_X4 FILLER_47_242 ();
 FILLCELL_X1 FILLER_47_246 ();
 FILLCELL_X1 FILLER_47_290 ();
 FILLCELL_X2 FILLER_47_301 ();
 FILLCELL_X2 FILLER_47_306 ();
 FILLCELL_X2 FILLER_47_311 ();
 FILLCELL_X1 FILLER_47_313 ();
 FILLCELL_X1 FILLER_47_321 ();
 FILLCELL_X2 FILLER_47_363 ();
 FILLCELL_X1 FILLER_48_13 ();
 FILLCELL_X1 FILLER_48_17 ();
 FILLCELL_X2 FILLER_48_30 ();
 FILLCELL_X1 FILLER_48_32 ();
 FILLCELL_X1 FILLER_48_72 ();
 FILLCELL_X2 FILLER_48_76 ();
 FILLCELL_X1 FILLER_48_78 ();
 FILLCELL_X1 FILLER_48_82 ();
 FILLCELL_X4 FILLER_48_104 ();
 FILLCELL_X2 FILLER_48_108 ();
 FILLCELL_X2 FILLER_48_113 ();
 FILLCELL_X2 FILLER_48_118 ();
 FILLCELL_X1 FILLER_48_120 ();
 FILLCELL_X2 FILLER_48_127 ();
 FILLCELL_X1 FILLER_48_129 ();
 FILLCELL_X2 FILLER_48_142 ();
 FILLCELL_X1 FILLER_48_144 ();
 FILLCELL_X4 FILLER_48_148 ();
 FILLCELL_X4 FILLER_48_155 ();
 FILLCELL_X8 FILLER_48_162 ();
 FILLCELL_X1 FILLER_48_170 ();
 FILLCELL_X4 FILLER_48_183 ();
 FILLCELL_X8 FILLER_48_193 ();
 FILLCELL_X2 FILLER_48_207 ();
 FILLCELL_X1 FILLER_48_209 ();
 FILLCELL_X4 FILLER_48_216 ();
 FILLCELL_X1 FILLER_48_223 ();
 FILLCELL_X4 FILLER_48_233 ();
 FILLCELL_X8 FILLER_48_243 ();
 FILLCELL_X2 FILLER_48_254 ();
 FILLCELL_X4 FILLER_48_259 ();
 FILLCELL_X2 FILLER_48_263 ();
 FILLCELL_X1 FILLER_48_265 ();
 FILLCELL_X2 FILLER_48_269 ();
 FILLCELL_X4 FILLER_48_274 ();
 FILLCELL_X8 FILLER_48_281 ();
 FILLCELL_X2 FILLER_48_298 ();
 FILLCELL_X1 FILLER_48_300 ();
 FILLCELL_X2 FILLER_48_313 ();
 FILLCELL_X1 FILLER_48_324 ();
 FILLCELL_X2 FILLER_48_331 ();
 FILLCELL_X1 FILLER_48_333 ();
endmodule
