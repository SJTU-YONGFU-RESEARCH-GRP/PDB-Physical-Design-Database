module parameterized_pwm (clk,
    enable,
    pwm_out,
    rst_n,
    div,
    duty);
 input clk;
 input enable;
 output pwm_out;
 input rst_n;
 input [15:0] div;
 input [7:0] duty;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \div_counter[0] ;
 wire \div_counter[10] ;
 wire \div_counter[11] ;
 wire \div_counter[12] ;
 wire \div_counter[13] ;
 wire \div_counter[14] ;
 wire \div_counter[15] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_counter[5] ;
 wire \div_counter[6] ;
 wire \div_counter[7] ;
 wire \div_counter[8] ;
 wire \div_counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_1 _211_ (.A(net1),
    .Y(_138_));
 sky130_fd_sc_hd__inv_1 _212_ (.A(\div_counter[1] ),
    .Y(_141_));
 sky130_fd_sc_hd__inv_1 _213_ (.A(\div_counter[3] ),
    .Y(_144_));
 sky130_fd_sc_hd__inv_1 _214_ (.A(\div_counter[2] ),
    .Y(_147_));
 sky130_fd_sc_hd__inv_1 _215_ (.A(\div_counter[7] ),
    .Y(_150_));
 sky130_fd_sc_hd__inv_1 _216_ (.A(\div_counter[6] ),
    .Y(_153_));
 sky130_fd_sc_hd__inv_1 _217_ (.A(\div_counter[5] ),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _218_ (.A(\div_counter[4] ),
    .Y(_159_));
 sky130_fd_sc_hd__inv_1 _219_ (.A(\div_counter[15] ),
    .Y(_162_));
 sky130_fd_sc_hd__inv_1 _220_ (.A(\div_counter[14] ),
    .Y(_165_));
 sky130_fd_sc_hd__inv_1 _221_ (.A(\div_counter[13] ),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _222_ (.A(\div_counter[12] ),
    .Y(_171_));
 sky130_fd_sc_hd__inv_1 _223_ (.A(\div_counter[11] ),
    .Y(_174_));
 sky130_fd_sc_hd__inv_1 _224_ (.A(\div_counter[10] ),
    .Y(_177_));
 sky130_fd_sc_hd__inv_1 _225_ (.A(\div_counter[9] ),
    .Y(_180_));
 sky130_fd_sc_hd__inv_1 _226_ (.A(\div_counter[8] ),
    .Y(_183_));
 sky130_fd_sc_hd__inv_1 _227_ (.A(net24),
    .Y(_190_));
 sky130_fd_sc_hd__inv_1 _228_ (.A(net23),
    .Y(_193_));
 sky130_fd_sc_hd__inv_1 _229_ (.A(net22),
    .Y(_196_));
 sky130_fd_sc_hd__inv_1 _230_ (.A(net21),
    .Y(_199_));
 sky130_fd_sc_hd__inv_1 _231_ (.A(net20),
    .Y(_202_));
 sky130_fd_sc_hd__inv_1 _232_ (.A(net19),
    .Y(_205_));
 sky130_fd_sc_hd__inv_1 _233_ (.A(net18),
    .Y(_208_));
 sky130_fd_sc_hd__nand4_2 _234_ (.A(_164_),
    .B(_173_),
    .C(_170_),
    .D(_167_),
    .Y(_025_));
 sky130_fd_sc_hd__a21oi_1 _235_ (.A1(_182_),
    .A2(_184_),
    .B1(_181_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_1 _236_ (.A(_176_),
    .B(_179_),
    .Y(_027_));
 sky130_fd_sc_hd__a21oi_1 _237_ (.A1(_176_),
    .A2(_178_),
    .B1(_175_),
    .Y(_028_));
 sky130_fd_sc_hd__o21ai_0 _238_ (.A1(_026_),
    .A2(_027_),
    .B1(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__nand2b_2 _239_ (.A_N(_025_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__nor2b_1 _240_ (.A(_139_),
    .B_N(_143_),
    .Y(_031_));
 sky130_fd_sc_hd__o211ai_1 _241_ (.A1(_142_),
    .A2(_031_),
    .B1(_146_),
    .C1(_149_),
    .Y(_032_));
 sky130_fd_sc_hd__a21oi_1 _242_ (.A1(_146_),
    .A2(_148_),
    .B1(_145_),
    .Y(_033_));
 sky130_fd_sc_hd__nand4_2 _243_ (.A(_176_),
    .B(_185_),
    .C(_182_),
    .D(_179_),
    .Y(_034_));
 sky130_fd_sc_hd__nand4_1 _244_ (.A(_152_),
    .B(_161_),
    .C(_158_),
    .D(_155_),
    .Y(_035_));
 sky130_fd_sc_hd__a2111o_2 _245_ (.A1(_032_),
    .A2(_033_),
    .B1(_025_),
    .C1(_034_),
    .D1(_035_),
    .X(_036_));
 sky130_fd_sc_hd__nor2_1 _246_ (.A(_025_),
    .B(_034_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _247_ (.A(_152_),
    .B(_155_),
    .Y(_038_));
 sky130_fd_sc_hd__a21oi_1 _248_ (.A1(_158_),
    .A2(_160_),
    .B1(_157_),
    .Y(_039_));
 sky130_fd_sc_hd__a21oi_1 _249_ (.A1(_152_),
    .A2(_154_),
    .B1(_151_),
    .Y(_040_));
 sky130_fd_sc_hd__o21ai_1 _250_ (.A1(_038_),
    .A2(_039_),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand3_1 _251_ (.A(_170_),
    .B(_167_),
    .C(_172_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_1 _252_ (.A1(_167_),
    .A2(_169_),
    .B1(_166_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _253_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__a221oi_4 _254_ (.A1(_037_),
    .A2(_041_),
    .B1(_044_),
    .B2(_164_),
    .C1(_163_),
    .Y(_045_));
 sky130_fd_sc_hd__nor4_1 _255_ (.A(net16),
    .B(net15),
    .C(net3),
    .D(net6),
    .Y(_046_));
 sky130_fd_sc_hd__nor4_1 _256_ (.A(net2),
    .B(net5),
    .C(net4),
    .D(net7),
    .Y(_047_));
 sky130_fd_sc_hd__nand2_1 _257_ (.A(_046_),
    .B(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__nor4_1 _258_ (.A(net8),
    .B(net1),
    .C(net10),
    .D(net13),
    .Y(_049_));
 sky130_fd_sc_hd__nor4_1 _259_ (.A(net9),
    .B(net12),
    .C(net11),
    .D(net14),
    .Y(_050_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(_049_),
    .B(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__nand4_1 _261_ (.A(_143_),
    .B(_140_),
    .C(_146_),
    .D(_149_),
    .Y(_052_));
 sky130_fd_sc_hd__nor4_2 _262_ (.A(_025_),
    .B(_034_),
    .C(_035_),
    .D(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__o21bai_1 _263_ (.A1(_048_),
    .A2(_051_),
    .B1_N(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__a31oi_4 _264_ (.A1(_030_),
    .A2(_036_),
    .A3(_045_),
    .B1(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__nand2b_1 _265_ (.A_N(_055_),
    .B(net25),
    .Y(_056_));
 sky130_fd_sc_hd__and3_1 _266_ (.A(\counter[2] ),
    .B(\counter[3] ),
    .C(_186_),
    .X(_057_));
 sky130_fd_sc_hd__and3_1 _267_ (.A(\counter[4] ),
    .B(\counter[5] ),
    .C(_057_),
    .X(_058_));
 sky130_fd_sc_hd__and3_1 _268_ (.A(\counter[6] ),
    .B(\counter[7] ),
    .C(_058_),
    .X(_059_));
 sky130_fd_sc_hd__or3b_1 _269_ (.A(\counter[0] ),
    .B(_059_),
    .C_N(net26),
    .X(_060_));
 sky130_fd_sc_hd__clkinv_2 _270_ (.A(net25),
    .Y(_061_));
 sky130_fd_sc_hd__buf_6 _271_ (.A(_055_),
    .X(_062_));
 sky130_fd_sc_hd__buf_2 _272_ (.A(net26),
    .X(_063_));
 sky130_fd_sc_hd__o211ai_1 _273_ (.A1(_061_),
    .A2(_062_),
    .B1(\counter[0] ),
    .C1(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__o21ai_0 _274_ (.A1(_056_),
    .A2(_060_),
    .B1(_064_),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _275_ (.A(net26),
    .B(_187_),
    .Y(_065_));
 sky130_fd_sc_hd__o211ai_1 _276_ (.A1(_061_),
    .A2(_062_),
    .B1(\counter[1] ),
    .C1(_063_),
    .Y(_066_));
 sky130_fd_sc_hd__o21ai_0 _277_ (.A1(_056_),
    .A2(_065_),
    .B1(_066_),
    .Y(_001_));
 sky130_fd_sc_hd__buf_2 _278_ (.A(net25),
    .X(_067_));
 sky130_fd_sc_hd__nand2_1 _279_ (.A(_067_),
    .B(_186_),
    .Y(_068_));
 sky130_fd_sc_hd__o21ai_0 _280_ (.A1(_062_),
    .A2(_068_),
    .B1(\counter[2] ),
    .Y(_069_));
 sky130_fd_sc_hd__or3_1 _281_ (.A(\counter[2] ),
    .B(_062_),
    .C(_068_),
    .X(_070_));
 sky130_fd_sc_hd__a21boi_0 _282_ (.A1(_069_),
    .A2(_070_),
    .B1_N(_063_),
    .Y(_002_));
 sky130_fd_sc_hd__and3_1 _283_ (.A(\counter[2] ),
    .B(\counter[0] ),
    .C(\counter[1] ),
    .X(_071_));
 sky130_fd_sc_hd__or4b_1 _284_ (.A(_061_),
    .B(\counter[3] ),
    .C(_055_),
    .D_N(_071_),
    .X(_072_));
 sky130_fd_sc_hd__o21ai_0 _285_ (.A1(_059_),
    .A2(_071_),
    .B1(_067_),
    .Y(_073_));
 sky130_fd_sc_hd__o21ai_0 _286_ (.A1(_062_),
    .A2(_073_),
    .B1(\counter[3] ),
    .Y(_074_));
 sky130_fd_sc_hd__a21boi_0 _287_ (.A1(_072_),
    .A2(_074_),
    .B1_N(_063_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _288_ (.A(_067_),
    .B(_057_),
    .Y(_075_));
 sky130_fd_sc_hd__o21ai_0 _289_ (.A1(_062_),
    .A2(_075_),
    .B1(\counter[4] ),
    .Y(_076_));
 sky130_fd_sc_hd__or3_1 _290_ (.A(\counter[4] ),
    .B(_062_),
    .C(_075_),
    .X(_077_));
 sky130_fd_sc_hd__a21boi_0 _291_ (.A1(_076_),
    .A2(_077_),
    .B1_N(_063_),
    .Y(_004_));
 sky130_fd_sc_hd__and3_1 _292_ (.A(\counter[4] ),
    .B(\counter[3] ),
    .C(_071_),
    .X(_078_));
 sky130_fd_sc_hd__or4b_1 _293_ (.A(_061_),
    .B(\counter[5] ),
    .C(_055_),
    .D_N(_078_),
    .X(_079_));
 sky130_fd_sc_hd__o21ai_0 _294_ (.A1(_059_),
    .A2(_078_),
    .B1(_067_),
    .Y(_080_));
 sky130_fd_sc_hd__o21ai_0 _295_ (.A1(_062_),
    .A2(_080_),
    .B1(\counter[5] ),
    .Y(_081_));
 sky130_fd_sc_hd__a21boi_0 _296_ (.A1(_079_),
    .A2(_081_),
    .B1_N(_063_),
    .Y(_005_));
 sky130_fd_sc_hd__nand2_1 _297_ (.A(_067_),
    .B(_058_),
    .Y(_082_));
 sky130_fd_sc_hd__o21ai_0 _298_ (.A1(_062_),
    .A2(_082_),
    .B1(\counter[6] ),
    .Y(_083_));
 sky130_fd_sc_hd__or3_1 _299_ (.A(\counter[6] ),
    .B(_055_),
    .C(_082_),
    .X(_084_));
 sky130_fd_sc_hd__a21boi_0 _300_ (.A1(_083_),
    .A2(_084_),
    .B1_N(_063_),
    .Y(_006_));
 sky130_fd_sc_hd__nand2_1 _301_ (.A(net26),
    .B(\counter[6] ),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_1 _302_ (.A(\counter[5] ),
    .B(_078_),
    .Y(_086_));
 sky130_fd_sc_hd__a21oi_1 _303_ (.A1(\counter[5] ),
    .A2(_078_),
    .B1(_058_),
    .Y(_087_));
 sky130_fd_sc_hd__nand2_1 _304_ (.A(_067_),
    .B(\counter[6] ),
    .Y(_088_));
 sky130_fd_sc_hd__o311ai_0 _305_ (.A1(_062_),
    .A2(_087_),
    .A3(_088_),
    .B1(\counter[7] ),
    .C1(_063_),
    .Y(_089_));
 sky130_fd_sc_hd__o41ai_1 _306_ (.A1(\counter[7] ),
    .A2(_056_),
    .A3(_085_),
    .A4(_086_),
    .B1(_089_),
    .Y(_007_));
 sky130_fd_sc_hd__a31oi_4 _307_ (.A1(_030_),
    .A2(_036_),
    .A3(_045_),
    .B1(_053_),
    .Y(_090_));
 sky130_fd_sc_hd__nor3b_1 _308_ (.A(_061_),
    .B(\div_counter[0] ),
    .C_N(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__nor2b_1 _309_ (.A(_067_),
    .B_N(\div_counter[0] ),
    .Y(_092_));
 sky130_fd_sc_hd__o21a_1 _310_ (.A1(_091_),
    .A2(_092_),
    .B1(_063_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _311_ (.A(net25),
    .B(_188_),
    .Y(_093_));
 sky130_fd_sc_hd__nand3_2 _312_ (.A(\div_counter[2] ),
    .B(\div_counter[3] ),
    .C(\div_counter[4] ),
    .Y(_094_));
 sky130_fd_sc_hd__nand3_1 _313_ (.A(\div_counter[5] ),
    .B(\div_counter[6] ),
    .C(\div_counter[7] ),
    .Y(_095_));
 sky130_fd_sc_hd__nor3_2 _314_ (.A(_093_),
    .B(_094_),
    .C(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__nand3_1 _315_ (.A(\div_counter[8] ),
    .B(\div_counter[9] ),
    .C(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__xnor2_1 _316_ (.A(_177_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__o21ai_2 _317_ (.A1(_061_),
    .A2(_090_),
    .B1(net26),
    .Y(_099_));
 sky130_fd_sc_hd__buf_2 _318_ (.A(_099_),
    .X(_100_));
 sky130_fd_sc_hd__nor2_1 _319_ (.A(_098_),
    .B(_100_),
    .Y(_009_));
 sky130_fd_sc_hd__nor3_1 _320_ (.A(_183_),
    .B(_180_),
    .C(_177_),
    .Y(_101_));
 sky130_fd_sc_hd__nand3_1 _321_ (.A(net25),
    .B(\div_counter[0] ),
    .C(\div_counter[1] ),
    .Y(_102_));
 sky130_fd_sc_hd__nor2_1 _322_ (.A(_094_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__and3b_1 _323_ (.A_N(_095_),
    .B(_101_),
    .C(_103_),
    .X(_104_));
 sky130_fd_sc_hd__xnor2_1 _324_ (.A(\div_counter[11] ),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__nor2_1 _325_ (.A(_100_),
    .B(_105_),
    .Y(_010_));
 sky130_fd_sc_hd__nand3_1 _326_ (.A(\div_counter[11] ),
    .B(_096_),
    .C(_101_),
    .Y(_106_));
 sky130_fd_sc_hd__xnor2_1 _327_ (.A(_171_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__nor2_1 _328_ (.A(_100_),
    .B(_107_),
    .Y(_011_));
 sky130_fd_sc_hd__nand3_1 _329_ (.A(\div_counter[11] ),
    .B(\div_counter[12] ),
    .C(_104_),
    .Y(_108_));
 sky130_fd_sc_hd__xnor2_1 _330_ (.A(_168_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _331_ (.A(_100_),
    .B(_109_),
    .Y(_012_));
 sky130_fd_sc_hd__nor3_1 _332_ (.A(_174_),
    .B(_171_),
    .C(_168_),
    .Y(_110_));
 sky130_fd_sc_hd__nand3_1 _333_ (.A(_096_),
    .B(_101_),
    .C(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__xnor2_1 _334_ (.A(_165_),
    .B(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__nor2_1 _335_ (.A(_100_),
    .B(_112_),
    .Y(_013_));
 sky130_fd_sc_hd__nand3_1 _336_ (.A(\div_counter[14] ),
    .B(_104_),
    .C(_110_),
    .Y(_113_));
 sky130_fd_sc_hd__xnor2_1 _337_ (.A(_162_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _338_ (.A(_100_),
    .B(_114_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_061_),
    .B(\div_counter[1] ),
    .Y(_115_));
 sky130_fd_sc_hd__nand3_1 _340_ (.A(_067_),
    .B(_189_),
    .C(_090_),
    .Y(_116_));
 sky130_fd_sc_hd__a21boi_0 _341_ (.A1(_115_),
    .A2(_116_),
    .B1_N(net26),
    .Y(_015_));
 sky130_fd_sc_hd__xnor2_1 _342_ (.A(_147_),
    .B(_093_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _343_ (.A(_100_),
    .B(_117_),
    .Y(_016_));
 sky130_fd_sc_hd__nand4_1 _344_ (.A(_067_),
    .B(\div_counter[0] ),
    .C(\div_counter[2] ),
    .D(\div_counter[1] ),
    .Y(_118_));
 sky130_fd_sc_hd__xnor2_1 _345_ (.A(_144_),
    .B(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _346_ (.A(_100_),
    .B(_119_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_1 _347_ (.A(_093_),
    .B(_094_),
    .Y(_120_));
 sky130_fd_sc_hd__a41oi_1 _348_ (.A1(_067_),
    .A2(_188_),
    .A3(\div_counter[2] ),
    .A4(\div_counter[3] ),
    .B1(\div_counter[4] ),
    .Y(_121_));
 sky130_fd_sc_hd__nor3_1 _349_ (.A(_120_),
    .B(_099_),
    .C(_121_),
    .Y(_018_));
 sky130_fd_sc_hd__xnor2_1 _350_ (.A(\div_counter[5] ),
    .B(_103_),
    .Y(_122_));
 sky130_fd_sc_hd__nor2_1 _351_ (.A(_100_),
    .B(_122_),
    .Y(_019_));
 sky130_fd_sc_hd__nand2_1 _352_ (.A(\div_counter[5] ),
    .B(_120_),
    .Y(_123_));
 sky130_fd_sc_hd__xnor2_1 _353_ (.A(_153_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__nor2_1 _354_ (.A(_100_),
    .B(_124_),
    .Y(_020_));
 sky130_fd_sc_hd__nand3_1 _355_ (.A(\div_counter[5] ),
    .B(\div_counter[6] ),
    .C(_103_),
    .Y(_125_));
 sky130_fd_sc_hd__xnor2_1 _356_ (.A(_150_),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_099_),
    .B(_126_),
    .Y(_021_));
 sky130_fd_sc_hd__xnor2_1 _358_ (.A(\div_counter[8] ),
    .B(_096_),
    .Y(_127_));
 sky130_fd_sc_hd__nor2_1 _359_ (.A(_099_),
    .B(_127_),
    .Y(_022_));
 sky130_fd_sc_hd__nor4_1 _360_ (.A(_183_),
    .B(_094_),
    .C(_095_),
    .D(_102_),
    .Y(_128_));
 sky130_fd_sc_hd__xnor2_1 _361_ (.A(\div_counter[9] ),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _362_ (.A(_099_),
    .B(_129_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2b_1 _363_ (.A_N(\counter[0] ),
    .B(net17),
    .Y(_130_));
 sky130_fd_sc_hd__a21o_1 _364_ (.A1(_210_),
    .A2(_130_),
    .B1(_209_),
    .X(_131_));
 sky130_fd_sc_hd__a21o_1 _365_ (.A1(_207_),
    .A2(_131_),
    .B1(_206_),
    .X(_132_));
 sky130_fd_sc_hd__a211oi_1 _366_ (.A1(_204_),
    .A2(_132_),
    .B1(_203_),
    .C1(_200_),
    .Y(_133_));
 sky130_fd_sc_hd__o21ai_0 _367_ (.A1(_200_),
    .A2(_201_),
    .B1(_198_),
    .Y(_134_));
 sky130_fd_sc_hd__o21bai_1 _368_ (.A1(_133_),
    .A2(_134_),
    .B1_N(_197_),
    .Y(_135_));
 sky130_fd_sc_hd__a211oi_1 _369_ (.A1(_192_),
    .A2(_194_),
    .B1(_191_),
    .C1(_061_),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(_063_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__a31oi_1 _371_ (.A1(_192_),
    .A2(_195_),
    .A3(_135_),
    .B1(_137_),
    .Y(_024_));
 sky130_fd_sc_hd__ha_1 _372_ (.A(_138_),
    .B(\div_counter[0] ),
    .COUT(_139_),
    .SUM(_140_));
 sky130_fd_sc_hd__ha_1 _373_ (.A(net8),
    .B(_141_),
    .COUT(_142_),
    .SUM(_143_));
 sky130_fd_sc_hd__ha_1 _374_ (.A(net10),
    .B(_144_),
    .COUT(_145_),
    .SUM(_146_));
 sky130_fd_sc_hd__ha_1 _375_ (.A(net9),
    .B(_147_),
    .COUT(_148_),
    .SUM(_149_));
 sky130_fd_sc_hd__ha_1 _376_ (.A(net14),
    .B(_150_),
    .COUT(_151_),
    .SUM(_152_));
 sky130_fd_sc_hd__ha_1 _377_ (.A(net13),
    .B(_153_),
    .COUT(_154_),
    .SUM(_155_));
 sky130_fd_sc_hd__ha_1 _378_ (.A(net12),
    .B(_156_),
    .COUT(_157_),
    .SUM(_158_));
 sky130_fd_sc_hd__ha_1 _379_ (.A(net11),
    .B(_159_),
    .COUT(_160_),
    .SUM(_161_));
 sky130_fd_sc_hd__ha_1 _380_ (.A(net7),
    .B(_162_),
    .COUT(_163_),
    .SUM(_164_));
 sky130_fd_sc_hd__ha_1 _381_ (.A(net6),
    .B(_165_),
    .COUT(_166_),
    .SUM(_167_));
 sky130_fd_sc_hd__ha_1 _382_ (.A(net5),
    .B(_168_),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__ha_1 _383_ (.A(net4),
    .B(_171_),
    .COUT(_172_),
    .SUM(_173_));
 sky130_fd_sc_hd__ha_1 _384_ (.A(net3),
    .B(_174_),
    .COUT(_175_),
    .SUM(_176_));
 sky130_fd_sc_hd__ha_1 _385_ (.A(net2),
    .B(_177_),
    .COUT(_178_),
    .SUM(_179_));
 sky130_fd_sc_hd__ha_1 _386_ (.A(net16),
    .B(_180_),
    .COUT(_181_),
    .SUM(_182_));
 sky130_fd_sc_hd__ha_1 _387_ (.A(net15),
    .B(_183_),
    .COUT(_184_),
    .SUM(_185_));
 sky130_fd_sc_hd__ha_1 _388_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .COUT(_186_),
    .SUM(_187_));
 sky130_fd_sc_hd__ha_1 _389_ (.A(\div_counter[0] ),
    .B(\div_counter[1] ),
    .COUT(_188_),
    .SUM(_189_));
 sky130_fd_sc_hd__ha_1 _390_ (.A(\counter[7] ),
    .B(_190_),
    .COUT(_191_),
    .SUM(_192_));
 sky130_fd_sc_hd__ha_1 _391_ (.A(\counter[6] ),
    .B(_193_),
    .COUT(_194_),
    .SUM(_195_));
 sky130_fd_sc_hd__ha_1 _392_ (.A(\counter[5] ),
    .B(_196_),
    .COUT(_197_),
    .SUM(_198_));
 sky130_fd_sc_hd__ha_1 _393_ (.A(\counter[4] ),
    .B(_199_),
    .COUT(_200_),
    .SUM(_201_));
 sky130_fd_sc_hd__ha_1 _394_ (.A(\counter[3] ),
    .B(_202_),
    .COUT(_203_),
    .SUM(_204_));
 sky130_fd_sc_hd__ha_1 _395_ (.A(\counter[2] ),
    .B(_205_),
    .COUT(_206_),
    .SUM(_207_));
 sky130_fd_sc_hd__ha_1 _396_ (.A(\counter[1] ),
    .B(_208_),
    .COUT(_209_),
    .SUM(_210_));
 sky130_fd_sc_hd__dfxtp_1 \counter[0]$_SDFFE_PN0P_  (.D(_000_),
    .Q(\counter[0] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[1]$_SDFFE_PN0P_  (.D(_001_),
    .Q(\counter[1] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[2]$_SDFFE_PN0P_  (.D(_002_),
    .Q(\counter[2] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[3]$_SDFFE_PN0P_  (.D(_003_),
    .Q(\counter[3] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[4]$_SDFFE_PN0P_  (.D(_004_),
    .Q(\counter[4] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[5]$_SDFFE_PN0P_  (.D(_005_),
    .Q(\counter[5] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[6]$_SDFFE_PN0P_  (.D(_006_),
    .Q(\counter[6] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \counter[7]$_SDFFE_PN0P_  (.D(_007_),
    .Q(\counter[7] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[0]$_SDFFE_PN0P_  (.D(_008_),
    .Q(\div_counter[0] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[10]$_SDFFE_PN0P_  (.D(_009_),
    .Q(\div_counter[10] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[11]$_SDFFE_PN0P_  (.D(_010_),
    .Q(\div_counter[11] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[12]$_SDFFE_PN0P_  (.D(_011_),
    .Q(\div_counter[12] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[13]$_SDFFE_PN0P_  (.D(_012_),
    .Q(\div_counter[13] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[14]$_SDFFE_PN0P_  (.D(_013_),
    .Q(\div_counter[14] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[15]$_SDFFE_PN0P_  (.D(_014_),
    .Q(\div_counter[15] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[1]$_SDFFE_PN0P_  (.D(_015_),
    .Q(\div_counter[1] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[2]$_SDFFE_PN0P_  (.D(_016_),
    .Q(\div_counter[2] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[3]$_SDFFE_PN0P_  (.D(_017_),
    .Q(\div_counter[3] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[4]$_SDFFE_PN0P_  (.D(_018_),
    .Q(\div_counter[4] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[5]$_SDFFE_PN0P_  (.D(_019_),
    .Q(\div_counter[5] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[6]$_SDFFE_PN0P_  (.D(_020_),
    .Q(\div_counter[6] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[7]$_SDFFE_PN0P_  (.D(_021_),
    .Q(\div_counter[7] ),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[8]$_SDFFE_PN0P_  (.D(_022_),
    .Q(\div_counter[8] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \div_counter[9]$_SDFFE_PN0P_  (.D(_023_),
    .Q(\div_counter[9] ),
    .CLK(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__dfxtp_1 \pwm_reg$_SDFF_PN0_  (.D(_024_),
    .Q(net27),
    .CLK(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_43 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(div[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(div[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(div[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(div[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(div[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(div[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(div[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(div[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(div[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(div[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(div[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(div[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(div[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(div[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(div[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(div[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(duty[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(duty[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(duty[2]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(duty[3]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(duty[4]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(duty[5]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(duty[6]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(duty[7]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(enable),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(rst_n),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(pwm_out));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
endmodule
