module i2c_master_top (arst_i,
    scl_pad_i,
    scl_pad_o,
    scl_padoen_o,
    sda_pad_i,
    sda_pad_o,
    sda_padoen_o,
    wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_inta_o,
    wb_rst_i,
    wb_stb_i,
    wb_we_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o);
 input arst_i;
 input scl_pad_i;
 output scl_pad_o;
 output scl_padoen_o;
 input sda_pad_i;
 output sda_pad_o;
 output sda_padoen_o;
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 output wb_inta_o;
 input wb_rst_i;
 input wb_stb_i;
 input wb_we_i;
 input [2:0] wb_adr_i;
 input [7:0] wb_dat_i;
 output [7:0] wb_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire clknet_0_wb_clk_i;
 wire ack;
 wire al;
 wire \byte_controller.ack_out ;
 wire \byte_controller.bit_controller.al ;
 wire \byte_controller.bit_controller.busy ;
 wire \byte_controller.bit_controller.c_state[0] ;
 wire \byte_controller.bit_controller.c_state[10] ;
 wire \byte_controller.bit_controller.c_state[11] ;
 wire \byte_controller.bit_controller.c_state[12] ;
 wire \byte_controller.bit_controller.c_state[13] ;
 wire \byte_controller.bit_controller.c_state[14] ;
 wire \byte_controller.bit_controller.c_state[15] ;
 wire \byte_controller.bit_controller.c_state[16] ;
 wire \byte_controller.bit_controller.c_state[1] ;
 wire \byte_controller.bit_controller.c_state[2] ;
 wire \byte_controller.bit_controller.c_state[3] ;
 wire \byte_controller.bit_controller.c_state[4] ;
 wire \byte_controller.bit_controller.c_state[5] ;
 wire \byte_controller.bit_controller.c_state[6] ;
 wire \byte_controller.bit_controller.c_state[7] ;
 wire \byte_controller.bit_controller.c_state[8] ;
 wire \byte_controller.bit_controller.c_state[9] ;
 wire \byte_controller.bit_controller.clk_cnt[0] ;
 wire \byte_controller.bit_controller.clk_cnt[10] ;
 wire \byte_controller.bit_controller.clk_cnt[11] ;
 wire \byte_controller.bit_controller.clk_cnt[12] ;
 wire \byte_controller.bit_controller.clk_cnt[13] ;
 wire \byte_controller.bit_controller.clk_cnt[14] ;
 wire \byte_controller.bit_controller.clk_cnt[15] ;
 wire \byte_controller.bit_controller.clk_cnt[1] ;
 wire \byte_controller.bit_controller.clk_cnt[2] ;
 wire \byte_controller.bit_controller.clk_cnt[3] ;
 wire \byte_controller.bit_controller.clk_cnt[4] ;
 wire \byte_controller.bit_controller.clk_cnt[5] ;
 wire \byte_controller.bit_controller.clk_cnt[6] ;
 wire \byte_controller.bit_controller.clk_cnt[7] ;
 wire \byte_controller.bit_controller.clk_cnt[8] ;
 wire \byte_controller.bit_controller.clk_cnt[9] ;
 wire \byte_controller.bit_controller.clk_en ;
 wire \byte_controller.bit_controller.cmd_ack ;
 wire \byte_controller.bit_controller.cmd_stop ;
 wire \byte_controller.bit_controller.cnt[0] ;
 wire \byte_controller.bit_controller.cnt[10] ;
 wire \byte_controller.bit_controller.cnt[11] ;
 wire \byte_controller.bit_controller.cnt[12] ;
 wire \byte_controller.bit_controller.cnt[13] ;
 wire \byte_controller.bit_controller.cnt[14] ;
 wire \byte_controller.bit_controller.cnt[15] ;
 wire \byte_controller.bit_controller.cnt[1] ;
 wire \byte_controller.bit_controller.cnt[2] ;
 wire \byte_controller.bit_controller.cnt[3] ;
 wire \byte_controller.bit_controller.cnt[4] ;
 wire \byte_controller.bit_controller.cnt[5] ;
 wire \byte_controller.bit_controller.cnt[6] ;
 wire \byte_controller.bit_controller.cnt[7] ;
 wire \byte_controller.bit_controller.cnt[8] ;
 wire \byte_controller.bit_controller.cnt[9] ;
 wire \byte_controller.bit_controller.dSCL ;
 wire \byte_controller.bit_controller.dSDA ;
 wire \byte_controller.bit_controller.din ;
 wire \byte_controller.bit_controller.dout ;
 wire \byte_controller.bit_controller.dscl_oen ;
 wire \byte_controller.bit_controller.ena ;
 wire \byte_controller.bit_controller.sSCL ;
 wire \byte_controller.bit_controller.sSDA ;
 wire \byte_controller.bit_controller.sda_chk ;
 wire \byte_controller.bit_controller.sta_condition ;
 wire \byte_controller.bit_controller.sto_condition ;
 wire \byte_controller.c_state[0] ;
 wire \byte_controller.c_state[1] ;
 wire \byte_controller.c_state[2] ;
 wire \byte_controller.c_state[3] ;
 wire \byte_controller.c_state[4] ;
 wire \byte_controller.c_state[5] ;
 wire \byte_controller.cmd_ack ;
 wire \byte_controller.core_cmd[1] ;
 wire \byte_controller.core_cmd[2] ;
 wire \byte_controller.core_cmd[3] ;
 wire \byte_controller.core_cmd[4] ;
 wire \byte_controller.dcnt[0] ;
 wire \byte_controller.dcnt[1] ;
 wire \byte_controller.dcnt[2] ;
 wire \byte_controller.din[0] ;
 wire \byte_controller.din[1] ;
 wire \byte_controller.din[2] ;
 wire \byte_controller.din[3] ;
 wire \byte_controller.din[4] ;
 wire \byte_controller.din[5] ;
 wire \byte_controller.din[6] ;
 wire \byte_controller.din[7] ;
 wire \byte_controller.dout[0] ;
 wire \byte_controller.dout[1] ;
 wire \byte_controller.dout[2] ;
 wire \byte_controller.dout[3] ;
 wire \byte_controller.dout[4] ;
 wire \byte_controller.dout[5] ;
 wire \byte_controller.dout[6] ;
 wire \byte_controller.dout[7] ;
 wire \byte_controller.ld ;
 wire \byte_controller.read ;
 wire \byte_controller.shift ;
 wire \byte_controller.start ;
 wire \byte_controller.stop ;
 wire \byte_controller.write ;
 wire \cr[0] ;
 wire \cr[1] ;
 wire \cr[2] ;
 wire \ctr[0] ;
 wire \ctr[1] ;
 wire \ctr[2] ;
 wire \ctr[3] ;
 wire \ctr[4] ;
 wire \ctr[5] ;
 wire \ctr[6] ;
 wire irq_flag;
 wire rxack;
 wire tip;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire net23;

 BUF_X2 _0801_ (.A(\byte_controller.bit_controller.al ),
    .Z(_0127_));
 OR2_X1 _0802_ (.A1(net6),
    .A2(_0127_),
    .ZN(_0128_));
 CLKBUF_X3 _0803_ (.A(_0128_),
    .Z(_0129_));
 CLKBUF_X2 _0804_ (.A(\byte_controller.start ),
    .Z(_0130_));
 BUF_X2 _0805_ (.A(\byte_controller.read ),
    .Z(_0131_));
 NOR2_X2 _0806_ (.A1(_0131_),
    .A2(\byte_controller.write ),
    .ZN(_0132_));
 INV_X1 _0807_ (.A(\byte_controller.stop ),
    .ZN(_0133_));
 AOI21_X2 _0808_ (.A(\byte_controller.cmd_ack ),
    .B1(_0132_),
    .B2(_0133_),
    .ZN(_0134_));
 NAND3_X1 _0809_ (.A1(_0130_),
    .A2(\byte_controller.c_state[0] ),
    .A3(_0134_),
    .ZN(_0135_));
 BUF_X1 _0810_ (.A(_0033_),
    .Z(_0136_));
 NAND2_X1 _0811_ (.A1(_0136_),
    .A2(\byte_controller.c_state[5] ),
    .ZN(_0137_));
 AOI21_X1 _0812_ (.A(_0129_),
    .B1(_0135_),
    .B2(_0137_),
    .ZN(_0011_));
 CLKBUF_X2 _0813_ (.A(\byte_controller.c_state[2] ),
    .Z(_0138_));
 BUF_X2 _0814_ (.A(\byte_controller.bit_controller.cmd_ack ),
    .Z(_0139_));
 INV_X1 _0815_ (.A(_0139_),
    .ZN(_0140_));
 NOR2_X1 _0816_ (.A1(_0140_),
    .A2(_0128_),
    .ZN(_0141_));
 AND3_X1 _0817_ (.A1(_0138_),
    .A2(\byte_controller.stop ),
    .A3(_0141_),
    .ZN(_0142_));
 NAND2_X1 _0818_ (.A1(\byte_controller.c_state[0] ),
    .A2(_0134_),
    .ZN(_0143_));
 NOR3_X2 _0819_ (.A1(_0130_),
    .A2(_0129_),
    .A3(_0143_),
    .ZN(_0144_));
 AOI21_X1 _0820_ (.A(_0142_),
    .B1(_0144_),
    .B2(_0132_),
    .ZN(_0145_));
 BUF_X4 _0821_ (.A(net6),
    .Z(_0146_));
 NOR2_X4 _0822_ (.A1(_0146_),
    .A2(_0127_),
    .ZN(_0147_));
 NAND3_X1 _0823_ (.A1(_0136_),
    .A2(\byte_controller.c_state[1] ),
    .A3(_0147_),
    .ZN(_0148_));
 NAND2_X1 _0824_ (.A1(_0145_),
    .A2(_0148_),
    .ZN(_0007_));
 INV_X1 _0825_ (.A(\byte_controller.c_state[0] ),
    .ZN(_0149_));
 NOR2_X1 _0826_ (.A1(_0149_),
    .A2(_0134_),
    .ZN(_0150_));
 INV_X1 _0827_ (.A(\byte_controller.c_state[3] ),
    .ZN(_0151_));
 INV_X1 _0828_ (.A(\byte_controller.c_state[4] ),
    .ZN(_0152_));
 NAND2_X1 _0829_ (.A1(_0151_),
    .A2(_0152_),
    .ZN(_0153_));
 NOR4_X1 _0830_ (.A1(_0138_),
    .A2(\byte_controller.c_state[5] ),
    .A3(\byte_controller.c_state[1] ),
    .A4(_0153_),
    .ZN(_0154_));
 MUX2_X1 _0831_ (.A(_0140_),
    .B(_0149_),
    .S(_0154_),
    .Z(_0155_));
 OAI21_X2 _0832_ (.A(_0147_),
    .B1(_0150_),
    .B2(_0155_),
    .ZN(_0156_));
 INV_X1 _0833_ (.A(\byte_controller.core_cmd[4] ),
    .ZN(_0157_));
 OAI22_X1 _0834_ (.A1(_0129_),
    .A2(_0135_),
    .B1(_0156_),
    .B2(_0157_),
    .ZN(_0015_));
 AOI21_X1 _0835_ (.A(\byte_controller.c_state[1] ),
    .B1(_0133_),
    .B2(_0138_),
    .ZN(_0158_));
 OAI221_X1 _0836_ (.A(_0147_),
    .B1(_0134_),
    .B2(_0149_),
    .C1(_0158_),
    .C2(_0140_),
    .ZN(_0006_));
 INV_X1 _0837_ (.A(\byte_controller.core_cmd[3] ),
    .ZN(_0159_));
 OAI21_X1 _0838_ (.A(_0145_),
    .B1(_0156_),
    .B2(_0159_),
    .ZN(_0014_));
 INV_X1 _0839_ (.A(\byte_controller.dcnt[2] ),
    .ZN(_0160_));
 NAND2_X1 _0840_ (.A1(_0160_),
    .A2(_0796_),
    .ZN(_0161_));
 MUX2_X1 _0841_ (.A(\byte_controller.c_state[4] ),
    .B(\byte_controller.c_state[3] ),
    .S(_0161_),
    .Z(_0162_));
 NAND2_X1 _0842_ (.A1(_0141_),
    .A2(_0162_),
    .ZN(_0163_));
 INV_X1 _0843_ (.A(\byte_controller.core_cmd[2] ),
    .ZN(_0164_));
 AND2_X1 _0844_ (.A1(\byte_controller.c_state[5] ),
    .A2(_0141_),
    .ZN(_0165_));
 AOI21_X1 _0845_ (.A(_0165_),
    .B1(_0144_),
    .B2(\byte_controller.write ),
    .ZN(_0166_));
 OAI221_X1 _0846_ (.A(_0163_),
    .B1(_0156_),
    .B2(_0164_),
    .C1(_0131_),
    .C2(_0166_),
    .ZN(_0013_));
 OAI21_X1 _0847_ (.A(_0131_),
    .B1(_0144_),
    .B2(_0165_),
    .ZN(_0167_));
 MUX2_X1 _0848_ (.A(\byte_controller.c_state[3] ),
    .B(\byte_controller.c_state[4] ),
    .S(_0161_),
    .Z(_0168_));
 INV_X1 _0849_ (.A(_0168_),
    .ZN(_0169_));
 NAND2_X1 _0850_ (.A1(_0139_),
    .A2(_0147_),
    .ZN(_0170_));
 INV_X1 _0851_ (.A(\byte_controller.core_cmd[1] ),
    .ZN(_0171_));
 OAI221_X1 _0852_ (.A(_0167_),
    .B1(_0169_),
    .B2(_0170_),
    .C1(_0156_),
    .C2(_0171_),
    .ZN(_0012_));
 OAI21_X1 _0853_ (.A(_0147_),
    .B1(_0161_),
    .B2(_0136_),
    .ZN(_0172_));
 OAI21_X1 _0854_ (.A(_0167_),
    .B1(_0172_),
    .B2(_0152_),
    .ZN(_0010_));
 OAI22_X1 _0855_ (.A1(_0131_),
    .A2(_0166_),
    .B1(_0172_),
    .B2(_0151_),
    .ZN(_0009_));
 NAND2_X1 _0856_ (.A1(_0138_),
    .A2(_0136_),
    .ZN(_0173_));
 NAND4_X1 _0857_ (.A1(_0139_),
    .A2(_0160_),
    .A3(_0796_),
    .A4(_0153_),
    .ZN(_0174_));
 AOI21_X1 _0858_ (.A(_0129_),
    .B1(_0173_),
    .B2(_0174_),
    .ZN(_0008_));
 INV_X1 _0859_ (.A(_0146_),
    .ZN(_0175_));
 CLKBUF_X3 _0860_ (.A(_0175_),
    .Z(_0176_));
 AND3_X1 _0861_ (.A1(_0176_),
    .A2(\ctr[6] ),
    .A3(irq_flag),
    .ZN(_0005_));
 CLKBUF_X3 _0862_ (.A(_0146_),
    .Z(_0177_));
 CLKBUF_X3 _0863_ (.A(_0177_),
    .Z(_0178_));
 NOR3_X1 _0864_ (.A1(_0127_),
    .A2(\byte_controller.cmd_ack ),
    .A3(irq_flag),
    .ZN(_0179_));
 NOR3_X1 _0865_ (.A1(_0178_),
    .A2(\cr[0] ),
    .A3(_0179_),
    .ZN(_0001_));
 CLKBUF_X3 _0866_ (.A(_0177_),
    .Z(_0180_));
 NOR2_X1 _0867_ (.A1(_0180_),
    .A2(_0132_),
    .ZN(_0003_));
 AND2_X1 _0868_ (.A1(_0176_),
    .A2(\byte_controller.ack_out ),
    .ZN(_0002_));
 INV_X1 _0869_ (.A(_0130_),
    .ZN(_0181_));
 AOI21_X1 _0870_ (.A(_0127_),
    .B1(_0181_),
    .B2(al),
    .ZN(_0182_));
 NOR2_X1 _0871_ (.A1(_0180_),
    .A2(_0182_),
    .ZN(_0000_));
 NAND2_X1 _0872_ (.A1(\byte_controller.bit_controller.clk_en ),
    .A2(_0147_),
    .ZN(_0183_));
 BUF_X2 _0873_ (.A(\byte_controller.bit_controller.c_state[4] ),
    .Z(_0184_));
 BUF_X2 _0874_ (.A(\byte_controller.bit_controller.c_state[5] ),
    .Z(_0185_));
 INV_X1 _0875_ (.A(_0185_),
    .ZN(_0186_));
 CLKBUF_X3 _0876_ (.A(\byte_controller.bit_controller.c_state[9] ),
    .Z(_0187_));
 CLKBUF_X3 _0877_ (.A(\byte_controller.bit_controller.c_state[8] ),
    .Z(_0188_));
 BUF_X4 _0878_ (.A(\byte_controller.bit_controller.c_state[11] ),
    .Z(_0189_));
 BUF_X4 _0879_ (.A(\byte_controller.bit_controller.c_state[10] ),
    .Z(_0190_));
 OR4_X4 _0880_ (.A1(_0187_),
    .A2(_0188_),
    .A3(_0189_),
    .A4(_0190_),
    .ZN(_0191_));
 CLKBUF_X3 _0881_ (.A(_0032_),
    .Z(_0192_));
 BUF_X2 _0882_ (.A(\byte_controller.bit_controller.c_state[2] ),
    .Z(_0193_));
 BUF_X2 _0883_ (.A(\byte_controller.bit_controller.c_state[3] ),
    .Z(_0194_));
 NOR2_X4 _0884_ (.A1(_0193_),
    .A2(_0194_),
    .ZN(_0195_));
 NAND2_X1 _0885_ (.A1(_0192_),
    .A2(_0195_),
    .ZN(_0196_));
 BUF_X2 _0886_ (.A(\byte_controller.bit_controller.c_state[13] ),
    .Z(_0197_));
 CLKBUF_X3 _0887_ (.A(\byte_controller.bit_controller.c_state[12] ),
    .Z(_0198_));
 NOR2_X4 _0888_ (.A1(_0197_),
    .A2(_0198_),
    .ZN(_0199_));
 BUF_X2 _0889_ (.A(\byte_controller.bit_controller.c_state[1] ),
    .Z(_0200_));
 BUF_X2 _0890_ (.A(\byte_controller.bit_controller.c_state[0] ),
    .Z(_0201_));
 BUF_X2 _0891_ (.A(\byte_controller.bit_controller.c_state[15] ),
    .Z(_0202_));
 BUF_X4 _0892_ (.A(\byte_controller.bit_controller.c_state[14] ),
    .Z(_0203_));
 NOR4_X4 _0893_ (.A1(_0200_),
    .A2(_0201_),
    .A3(_0202_),
    .A4(_0203_),
    .ZN(_0204_));
 BUF_X2 _0894_ (.A(\byte_controller.bit_controller.c_state[7] ),
    .Z(_0205_));
 BUF_X2 _0895_ (.A(\byte_controller.bit_controller.c_state[6] ),
    .Z(_0206_));
 NOR2_X1 _0896_ (.A1(_0205_),
    .A2(_0206_),
    .ZN(_0207_));
 NAND3_X1 _0897_ (.A1(_0199_),
    .A2(_0204_),
    .A3(_0207_),
    .ZN(_0208_));
 NOR3_X1 _0898_ (.A1(_0191_),
    .A2(_0196_),
    .A3(_0208_),
    .ZN(_0209_));
 NAND3_X1 _0899_ (.A1(_0184_),
    .A2(_0186_),
    .A3(_0209_),
    .ZN(_0210_));
 NOR4_X4 _0900_ (.A1(_0187_),
    .A2(_0188_),
    .A3(_0189_),
    .A4(_0190_),
    .ZN(_0211_));
 NAND2_X2 _0901_ (.A1(_0199_),
    .A2(_0211_),
    .ZN(_0212_));
 NOR4_X4 _0902_ (.A1(_0184_),
    .A2(_0185_),
    .A3(_0205_),
    .A4(_0206_),
    .ZN(_0213_));
 NAND2_X1 _0903_ (.A1(_0204_),
    .A2(_0213_),
    .ZN(_0214_));
 NAND2_X1 _0904_ (.A1(\byte_controller.bit_controller.c_state[16] ),
    .A2(_0195_),
    .ZN(_0215_));
 NOR3_X2 _0905_ (.A1(_0212_),
    .A2(_0214_),
    .A3(_0215_),
    .ZN(_0216_));
 NAND4_X4 _0906_ (.A1(_0192_),
    .A2(_0204_),
    .A3(_0213_),
    .A4(_0195_),
    .ZN(_0217_));
 INV_X1 _0907_ (.A(_0197_),
    .ZN(_0218_));
 NAND2_X1 _0908_ (.A1(_0218_),
    .A2(_0198_),
    .ZN(_0219_));
 NOR3_X1 _0909_ (.A1(_0191_),
    .A2(_0217_),
    .A3(_0219_),
    .ZN(_0220_));
 NAND3_X1 _0910_ (.A1(_0192_),
    .A2(_0199_),
    .A3(_0195_),
    .ZN(_0221_));
 NOR2_X1 _0911_ (.A1(_0189_),
    .A2(_0190_),
    .ZN(_0222_));
 NAND2_X1 _0912_ (.A1(_0188_),
    .A2(_0222_),
    .ZN(_0223_));
 NOR4_X1 _0913_ (.A1(_0187_),
    .A2(_0214_),
    .A3(_0221_),
    .A4(_0223_),
    .ZN(_0224_));
 NOR3_X1 _0914_ (.A1(_0216_),
    .A2(_0220_),
    .A3(_0224_),
    .ZN(_0225_));
 AOI21_X1 _0915_ (.A(_0183_),
    .B1(_0210_),
    .B2(_0225_),
    .ZN(_0023_));
 NAND2_X1 _0916_ (.A1(_0176_),
    .A2(\byte_controller.bit_controller.sto_condition ),
    .ZN(_0226_));
 NOR2_X1 _0917_ (.A1(_0212_),
    .A2(_0217_),
    .ZN(_0227_));
 INV_X1 _0918_ (.A(\byte_controller.bit_controller.sSDA ),
    .ZN(_0228_));
 NAND2_X1 _0919_ (.A1(_0175_),
    .A2(_0228_),
    .ZN(_0025_));
 INV_X1 _0920_ (.A(\byte_controller.bit_controller.sda_chk ),
    .ZN(_0229_));
 INV_X1 _0921_ (.A(net10),
    .ZN(_0230_));
 OAI33_X1 _0922_ (.A1(\byte_controller.bit_controller.cmd_stop ),
    .A2(_0226_),
    .A3(_0227_),
    .B1(_0025_),
    .B2(_0229_),
    .B3(_0230_),
    .ZN(_0020_));
 NOR2_X1 _0923_ (.A1(\byte_controller.bit_controller.busy ),
    .A2(\byte_controller.bit_controller.sta_condition ),
    .ZN(_0231_));
 NOR3_X1 _0924_ (.A1(_0178_),
    .A2(\byte_controller.bit_controller.sto_condition ),
    .A3(_0231_),
    .ZN(_0021_));
 NOR4_X1 _0925_ (.A1(_0177_),
    .A2(_0228_),
    .A3(\byte_controller.bit_controller.dSDA ),
    .A4(_0034_),
    .ZN(_0029_));
 INV_X1 _0926_ (.A(\byte_controller.bit_controller.dSDA ),
    .ZN(_0232_));
 NOR3_X1 _0927_ (.A1(_0232_),
    .A2(_0034_),
    .A3(_0025_),
    .ZN(_0028_));
 CLKBUF_X2 _0928_ (.A(ack),
    .Z(_0233_));
 CLKBUF_X2 _0929_ (.A(\byte_controller.dout[7] ),
    .Z(_0234_));
 NOR3_X1 _0930_ (.A1(_0139_),
    .A2(_0233_),
    .A3(_0234_),
    .ZN(_0235_));
 OR2_X1 _0931_ (.A1(_0129_),
    .A2(_0235_),
    .ZN(_0236_));
 NOR2_X1 _0932_ (.A1(_0139_),
    .A2(_0233_),
    .ZN(_0237_));
 OAI21_X1 _0933_ (.A(_0138_),
    .B1(_0237_),
    .B2(_0030_),
    .ZN(_0238_));
 OAI21_X1 _0934_ (.A(_0238_),
    .B1(_0234_),
    .B2(_0138_),
    .ZN(_0239_));
 NAND2_X1 _0935_ (.A1(_0139_),
    .A2(\byte_controller.c_state[4] ),
    .ZN(_0240_));
 OAI22_X2 _0936_ (.A1(_0139_),
    .A2(_0234_),
    .B1(_0240_),
    .B2(_0233_),
    .ZN(_0241_));
 AOI221_X2 _0937_ (.A(_0236_),
    .B1(_0239_),
    .B2(_0152_),
    .C1(_0030_),
    .C2(_0241_),
    .ZN(_0017_));
 INV_X1 _0938_ (.A(_0136_),
    .ZN(_0242_));
 NAND3_X1 _0939_ (.A1(_0242_),
    .A2(\byte_controller.c_state[3] ),
    .A3(_0161_),
    .ZN(_0243_));
 AOI21_X1 _0940_ (.A(_0129_),
    .B1(_0240_),
    .B2(_0243_),
    .ZN(_0019_));
 NAND2_X1 _0941_ (.A1(_0139_),
    .A2(\byte_controller.c_state[5] ),
    .ZN(_0244_));
 AOI21_X1 _0942_ (.A(_0129_),
    .B1(_0143_),
    .B2(_0244_),
    .ZN(_0018_));
 NOR2_X1 _0943_ (.A1(_0170_),
    .A2(_0158_),
    .ZN(_0016_));
 BUF_X4 _0944_ (.A(net4),
    .Z(_0245_));
 CLKBUF_X3 _0945_ (.A(wb_adr_i[0]),
    .Z(_0246_));
 INV_X4 _0946_ (.A(_0246_),
    .ZN(_0247_));
 NOR2_X1 _0947_ (.A1(_0245_),
    .A2(_0247_),
    .ZN(_0248_));
 BUF_X4 _0948_ (.A(wb_adr_i[1]),
    .Z(_0249_));
 MUX2_X1 _0949_ (.A(\byte_controller.bit_controller.clk_cnt[8] ),
    .B(\byte_controller.dout[0] ),
    .S(_0249_),
    .Z(_0250_));
 NAND2_X1 _0950_ (.A1(_0248_),
    .A2(_0250_),
    .ZN(_0251_));
 INV_X1 _0951_ (.A(\ctr[0] ),
    .ZN(_0252_));
 AOI21_X1 _0952_ (.A(_0245_),
    .B1(_0249_),
    .B2(_0252_),
    .ZN(_0253_));
 INV_X4 _0953_ (.A(_0249_),
    .ZN(_0254_));
 AOI21_X1 _0954_ (.A(_0253_),
    .B1(irq_flag),
    .B2(_0254_),
    .ZN(_0255_));
 BUF_X4 _0955_ (.A(_0246_),
    .Z(_0256_));
 OAI21_X1 _0956_ (.A(_0251_),
    .B1(_0255_),
    .B2(_0256_),
    .ZN(_0257_));
 NOR2_X4 _0957_ (.A1(_0249_),
    .A2(_0247_),
    .ZN(_0258_));
 NOR2_X4 _0958_ (.A1(_0254_),
    .A2(_0246_),
    .ZN(_0259_));
 AOI221_X1 _0959_ (.A(_0257_),
    .B1(_0258_),
    .B2(\byte_controller.din[0] ),
    .C1(_0259_),
    .C2(\cr[0] ),
    .ZN(_0260_));
 NAND2_X4 _0960_ (.A1(_0254_),
    .A2(_0247_),
    .ZN(_0261_));
 OAI21_X1 _0961_ (.A(_0257_),
    .B1(_0261_),
    .B2(\byte_controller.bit_controller.clk_cnt[0] ),
    .ZN(_0262_));
 INV_X2 _0962_ (.A(_0245_),
    .ZN(_0263_));
 CLKBUF_X3 _0963_ (.A(_0263_),
    .Z(_0264_));
 AOI21_X1 _0964_ (.A(_0260_),
    .B1(_0262_),
    .B2(_0264_),
    .ZN(_0664_));
 BUF_X4 _0965_ (.A(_0249_),
    .Z(_0265_));
 MUX2_X1 _0966_ (.A(\byte_controller.bit_controller.clk_cnt[1] ),
    .B(\ctr[1] ),
    .S(_0265_),
    .Z(_0266_));
 MUX2_X1 _0967_ (.A(tip),
    .B(\cr[1] ),
    .S(_0265_),
    .Z(_0267_));
 MUX2_X1 _0968_ (.A(_0266_),
    .B(_0267_),
    .S(_0245_),
    .Z(_0268_));
 NAND2_X1 _0969_ (.A1(_0247_),
    .A2(_0268_),
    .ZN(_0269_));
 MUX2_X1 _0970_ (.A(\byte_controller.bit_controller.clk_cnt[9] ),
    .B(\byte_controller.dout[1] ),
    .S(_0265_),
    .Z(_0270_));
 NOR2_X1 _0971_ (.A1(_0263_),
    .A2(_0249_),
    .ZN(_0271_));
 AOI22_X1 _0972_ (.A1(_0263_),
    .A2(_0270_),
    .B1(_0271_),
    .B2(\byte_controller.din[1] ),
    .ZN(_0272_));
 OAI21_X1 _0973_ (.A(_0269_),
    .B1(_0272_),
    .B2(_0247_),
    .ZN(_0665_));
 MUX2_X1 _0974_ (.A(\byte_controller.bit_controller.clk_cnt[2] ),
    .B(\byte_controller.bit_controller.clk_cnt[10] ),
    .S(_0256_),
    .Z(_0273_));
 MUX2_X1 _0975_ (.A(\ctr[2] ),
    .B(\byte_controller.dout[2] ),
    .S(_0256_),
    .Z(_0274_));
 MUX2_X1 _0976_ (.A(_0273_),
    .B(_0274_),
    .S(_0265_),
    .Z(_0275_));
 NAND2_X1 _0977_ (.A1(_0264_),
    .A2(_0275_),
    .ZN(_0276_));
 AOI22_X1 _0978_ (.A1(\byte_controller.din[2] ),
    .A2(_0258_),
    .B1(_0259_),
    .B2(\cr[2] ),
    .ZN(_0277_));
 OAI21_X1 _0979_ (.A(_0276_),
    .B1(_0277_),
    .B2(_0264_),
    .ZN(_0666_));
 MUX2_X1 _0980_ (.A(\byte_controller.bit_controller.clk_cnt[3] ),
    .B(\byte_controller.bit_controller.clk_cnt[11] ),
    .S(_0256_),
    .Z(_0278_));
 MUX2_X1 _0981_ (.A(\ctr[3] ),
    .B(\byte_controller.dout[3] ),
    .S(_0256_),
    .Z(_0279_));
 MUX2_X1 _0982_ (.A(_0278_),
    .B(_0279_),
    .S(_0265_),
    .Z(_0280_));
 NAND2_X1 _0983_ (.A1(_0264_),
    .A2(_0280_),
    .ZN(_0281_));
 AOI22_X1 _0984_ (.A1(\byte_controller.din[3] ),
    .A2(_0258_),
    .B1(_0259_),
    .B2(_0233_),
    .ZN(_0282_));
 OAI21_X1 _0985_ (.A(_0281_),
    .B1(_0282_),
    .B2(_0264_),
    .ZN(_0667_));
 MUX2_X1 _0986_ (.A(\byte_controller.bit_controller.clk_cnt[4] ),
    .B(\byte_controller.bit_controller.clk_cnt[12] ),
    .S(_0246_),
    .Z(_0283_));
 MUX2_X1 _0987_ (.A(\ctr[4] ),
    .B(\byte_controller.dout[4] ),
    .S(_0256_),
    .Z(_0284_));
 MUX2_X1 _0988_ (.A(_0283_),
    .B(_0284_),
    .S(_0265_),
    .Z(_0285_));
 NAND2_X1 _0989_ (.A1(_0264_),
    .A2(_0285_),
    .ZN(_0286_));
 AOI22_X1 _0990_ (.A1(\byte_controller.din[4] ),
    .A2(_0258_),
    .B1(_0259_),
    .B2(\byte_controller.write ),
    .ZN(_0287_));
 OAI21_X1 _0991_ (.A(_0286_),
    .B1(_0287_),
    .B2(_0264_),
    .ZN(_0668_));
 MUX2_X1 _0992_ (.A(\byte_controller.bit_controller.clk_cnt[13] ),
    .B(\byte_controller.dout[5] ),
    .S(_0249_),
    .Z(_0288_));
 NAND2_X1 _0993_ (.A1(_0248_),
    .A2(_0288_),
    .ZN(_0289_));
 INV_X1 _0994_ (.A(\ctr[5] ),
    .ZN(_0290_));
 AOI21_X1 _0995_ (.A(net4),
    .B1(_0249_),
    .B2(_0290_),
    .ZN(_0291_));
 AOI21_X1 _0996_ (.A(_0291_),
    .B1(al),
    .B2(_0254_),
    .ZN(_0292_));
 OAI21_X1 _0997_ (.A(_0289_),
    .B1(_0292_),
    .B2(_0256_),
    .ZN(_0293_));
 AOI221_X1 _0998_ (.A(_0293_),
    .B1(_0258_),
    .B2(\byte_controller.din[5] ),
    .C1(_0131_),
    .C2(_0259_),
    .ZN(_0294_));
 OAI21_X1 _0999_ (.A(_0293_),
    .B1(_0261_),
    .B2(\byte_controller.bit_controller.clk_cnt[5] ),
    .ZN(_0295_));
 AOI21_X1 _1000_ (.A(_0294_),
    .B1(_0295_),
    .B2(_0264_),
    .ZN(_0669_));
 MUX2_X1 _1001_ (.A(\byte_controller.bit_controller.clk_cnt[6] ),
    .B(\byte_controller.bit_controller.clk_cnt[14] ),
    .S(_0246_),
    .Z(_0296_));
 MUX2_X1 _1002_ (.A(\ctr[6] ),
    .B(\byte_controller.dout[6] ),
    .S(_0256_),
    .Z(_0297_));
 MUX2_X1 _1003_ (.A(_0296_),
    .B(_0297_),
    .S(_0265_),
    .Z(_0298_));
 NAND2_X1 _1004_ (.A1(_0264_),
    .A2(_0298_),
    .ZN(_0299_));
 MUX2_X1 _1005_ (.A(\byte_controller.bit_controller.busy ),
    .B(\byte_controller.din[6] ),
    .S(_0256_),
    .Z(_0300_));
 AOI22_X1 _1006_ (.A1(\byte_controller.stop ),
    .A2(_0259_),
    .B1(_0300_),
    .B2(_0254_),
    .ZN(_0301_));
 OAI21_X1 _1007_ (.A(_0299_),
    .B1(_0301_),
    .B2(_0264_),
    .ZN(_0670_));
 MUX2_X1 _1008_ (.A(\byte_controller.bit_controller.clk_cnt[15] ),
    .B(_0234_),
    .S(_0249_),
    .Z(_0302_));
 AOI221_X1 _1009_ (.A(_0247_),
    .B1(\byte_controller.din[7] ),
    .B2(_0271_),
    .C1(_0302_),
    .C2(_0263_),
    .ZN(_0303_));
 NAND2_X1 _1010_ (.A1(_0265_),
    .A2(_0130_),
    .ZN(_0304_));
 NAND2_X1 _1011_ (.A1(_0254_),
    .A2(rxack),
    .ZN(_0305_));
 NAND3_X1 _1012_ (.A1(_0245_),
    .A2(_0304_),
    .A3(_0305_),
    .ZN(_0306_));
 BUF_X2 _1013_ (.A(\byte_controller.bit_controller.ena ),
    .Z(_0307_));
 MUX2_X1 _1014_ (.A(\byte_controller.bit_controller.clk_cnt[7] ),
    .B(_0307_),
    .S(_0265_),
    .Z(_0308_));
 OAI21_X1 _1015_ (.A(_0306_),
    .B1(_0308_),
    .B2(_0245_),
    .ZN(_0309_));
 AOI21_X1 _1016_ (.A(_0303_),
    .B1(_0309_),
    .B2(_0247_),
    .ZN(_0671_));
 NAND2_X1 _1017_ (.A1(net7),
    .A2(net5),
    .ZN(_0310_));
 NOR2_X1 _1018_ (.A1(net11),
    .A2(_0310_),
    .ZN(_0004_));
 NOR2_X2 _1019_ (.A1(_0146_),
    .A2(\byte_controller.bit_controller.sSCL ),
    .ZN(_0311_));
 INV_X1 _1020_ (.A(_0311_),
    .ZN(_0024_));
 BUF_X2 _1021_ (.A(_0146_),
    .Z(_0312_));
 OR2_X1 _1022_ (.A1(_0312_),
    .A2(net3),
    .ZN(_0027_));
 OR2_X1 _1023_ (.A1(_0312_),
    .A2(net2),
    .ZN(_0026_));
 INV_X1 _1024_ (.A(\byte_controller.bit_controller.cnt[15] ),
    .ZN(_0313_));
 INV_X1 _1025_ (.A(\byte_controller.bit_controller.cnt[14] ),
    .ZN(_0314_));
 BUF_X2 _1026_ (.A(\byte_controller.bit_controller.cnt[11] ),
    .Z(_0315_));
 NOR3_X4 _1027_ (.A1(_0315_),
    .A2(\byte_controller.bit_controller.cnt[13] ),
    .A3(\byte_controller.bit_controller.cnt[12] ),
    .ZN(_0316_));
 NAND3_X2 _1028_ (.A1(_0313_),
    .A2(_0314_),
    .A3(_0316_),
    .ZN(_0317_));
 INV_X1 _1029_ (.A(\byte_controller.bit_controller.cnt[4] ),
    .ZN(_0318_));
 CLKBUF_X2 _1030_ (.A(\byte_controller.bit_controller.cnt[2] ),
    .Z(_0319_));
 NOR2_X2 _1031_ (.A1(\byte_controller.bit_controller.cnt[3] ),
    .A2(_0319_),
    .ZN(_0320_));
 CLKBUF_X2 _1032_ (.A(\byte_controller.bit_controller.cnt[5] ),
    .Z(_0321_));
 NOR3_X2 _1033_ (.A1(_0321_),
    .A2(\byte_controller.bit_controller.cnt[7] ),
    .A3(\byte_controller.bit_controller.cnt[6] ),
    .ZN(_0322_));
 NAND4_X2 _1034_ (.A1(_0792_),
    .A2(_0318_),
    .A3(_0320_),
    .A4(_0322_),
    .ZN(_0323_));
 CLKBUF_X2 _1035_ (.A(\byte_controller.bit_controller.cnt[8] ),
    .Z(_0324_));
 NOR3_X1 _1036_ (.A1(\byte_controller.bit_controller.cnt[9] ),
    .A2(_0324_),
    .A3(\byte_controller.bit_controller.cnt[10] ),
    .ZN(_0325_));
 INV_X1 _1037_ (.A(_0325_),
    .ZN(_0326_));
 OR2_X2 _1038_ (.A1(_0323_),
    .A2(_0326_),
    .ZN(_0327_));
 OAI21_X4 _1039_ (.A(_0307_),
    .B1(_0317_),
    .B2(_0327_),
    .ZN(_0328_));
 NOR2_X1 _1040_ (.A1(_0146_),
    .A2(_0328_),
    .ZN(_0329_));
 CLKBUF_X3 _1041_ (.A(_0329_),
    .Z(_0330_));
 AOI21_X1 _1042_ (.A(_0330_),
    .B1(_0311_),
    .B2(\byte_controller.bit_controller.dscl_oen ),
    .ZN(_0022_));
 AOI21_X1 _1043_ (.A(_0030_),
    .B1(_0138_),
    .B2(_0140_),
    .ZN(_0331_));
 MUX2_X1 _1044_ (.A(\byte_controller.ack_out ),
    .B(\byte_controller.bit_controller.dout ),
    .S(_0331_),
    .Z(_0332_));
 AND2_X1 _1045_ (.A1(_0147_),
    .A2(_0332_),
    .ZN(_0037_));
 INV_X1 _1046_ (.A(_0031_),
    .ZN(_0333_));
 OR2_X1 _1047_ (.A1(_0197_),
    .A2(_0198_),
    .ZN(_0334_));
 INV_X1 _1048_ (.A(_0188_),
    .ZN(_0335_));
 NAND3_X1 _1049_ (.A1(_0187_),
    .A2(_0335_),
    .A3(_0222_),
    .ZN(_0336_));
 INV_X1 _1050_ (.A(_0187_),
    .ZN(_0337_));
 OAI21_X1 _1051_ (.A(_0188_),
    .B1(_0189_),
    .B2(_0190_),
    .ZN(_0338_));
 XOR2_X2 _1052_ (.A(_0189_),
    .B(_0190_),
    .Z(_0339_));
 OAI211_X2 _1053_ (.A(_0337_),
    .B(_0338_),
    .C1(_0339_),
    .C2(_0188_),
    .ZN(_0340_));
 AOI211_X2 _1054_ (.A(_0334_),
    .B(_0217_),
    .C1(_0336_),
    .C2(_0340_),
    .ZN(_0341_));
 OR2_X1 _1055_ (.A1(_0202_),
    .A2(_0203_),
    .ZN(_0342_));
 NAND3_X4 _1056_ (.A1(_0192_),
    .A2(_0213_),
    .A3(_0195_),
    .ZN(_0343_));
 XNOR2_X1 _1057_ (.A(_0200_),
    .B(_0201_),
    .ZN(_0344_));
 NOR4_X1 _1058_ (.A1(_0212_),
    .A2(_0342_),
    .A3(_0343_),
    .A4(_0344_),
    .ZN(_0345_));
 OR3_X1 _1059_ (.A1(_0128_),
    .A2(_0341_),
    .A3(_0345_),
    .ZN(_0346_));
 XNOR2_X1 _1060_ (.A(_0184_),
    .B(_0185_),
    .ZN(_0347_));
 NOR4_X1 _1061_ (.A1(_0191_),
    .A2(_0196_),
    .A3(_0208_),
    .A4(_0347_),
    .ZN(_0348_));
 INV_X1 _1062_ (.A(_0213_),
    .ZN(_0349_));
 NAND3_X1 _1063_ (.A1(_0199_),
    .A2(_0211_),
    .A3(_0204_),
    .ZN(_0350_));
 NOR3_X1 _1064_ (.A1(_0349_),
    .A2(_0215_),
    .A3(_0350_),
    .ZN(_0351_));
 XNOR2_X1 _1065_ (.A(_0197_),
    .B(_0198_),
    .ZN(_0352_));
 NAND2_X1 _1066_ (.A1(_0211_),
    .A2(_0204_),
    .ZN(_0353_));
 NOR3_X1 _1067_ (.A1(_0343_),
    .A2(_0352_),
    .A3(_0353_),
    .ZN(_0354_));
 OR3_X1 _1068_ (.A1(_0348_),
    .A2(_0351_),
    .A3(_0354_),
    .ZN(_0355_));
 XNOR2_X1 _1069_ (.A(_0202_),
    .B(_0203_),
    .ZN(_0356_));
 OR2_X1 _1070_ (.A1(_0200_),
    .A2(_0201_),
    .ZN(_0357_));
 OR3_X1 _1071_ (.A1(_0334_),
    .A2(_0191_),
    .A3(_0357_),
    .ZN(_0358_));
 OR3_X1 _1072_ (.A1(_0343_),
    .A2(_0356_),
    .A3(_0358_),
    .ZN(_0359_));
 OR4_X2 _1073_ (.A1(_0184_),
    .A2(_0185_),
    .A3(_0196_),
    .A4(_0350_),
    .ZN(_0360_));
 INV_X1 _1074_ (.A(_0205_),
    .ZN(_0361_));
 INV_X1 _1075_ (.A(_0206_),
    .ZN(_0362_));
 NOR2_X1 _1076_ (.A1(_0361_),
    .A2(_0362_),
    .ZN(_0363_));
 XNOR2_X1 _1077_ (.A(_0193_),
    .B(_0194_),
    .ZN(_0364_));
 AND2_X1 _1078_ (.A1(_0204_),
    .A2(_0213_),
    .ZN(_0365_));
 NAND4_X4 _1079_ (.A1(_0192_),
    .A2(_0199_),
    .A3(_0211_),
    .A4(_0365_),
    .ZN(_0366_));
 OAI221_X1 _1080_ (.A(_0359_),
    .B1(_0360_),
    .B2(_0363_),
    .C1(_0364_),
    .C2(_0366_),
    .ZN(_0367_));
 OAI33_X1 _1081_ (.A1(_0146_),
    .A2(_0127_),
    .A3(_0333_),
    .B1(_0346_),
    .B2(_0355_),
    .B3(_0367_),
    .ZN(_0368_));
 BUF_X4 _1082_ (.A(_0368_),
    .Z(_0369_));
 BUF_X8 _1083_ (.A(_0369_),
    .Z(_0370_));
 NAND2_X1 _1084_ (.A1(_0201_),
    .A2(_0370_),
    .ZN(_0371_));
 NAND2_X1 _1085_ (.A1(_0031_),
    .A2(_0147_),
    .ZN(_0372_));
 NAND2_X1 _1086_ (.A1(_0207_),
    .A2(_0372_),
    .ZN(_0373_));
 OR4_X2 _1087_ (.A1(_0346_),
    .A2(_0355_),
    .A3(_0360_),
    .A4(_0373_),
    .ZN(_0374_));
 OAI21_X1 _1088_ (.A(_0371_),
    .B1(_0374_),
    .B2(_0157_),
    .ZN(_0038_));
 NOR2_X2 _1089_ (.A1(_0031_),
    .A2(_0129_),
    .ZN(_0375_));
 CLKBUF_X3 _1090_ (.A(_0375_),
    .Z(_0376_));
 NAND2_X1 _1091_ (.A1(_0199_),
    .A2(_0204_),
    .ZN(_0377_));
 NOR3_X1 _1092_ (.A1(_0343_),
    .A2(_0377_),
    .A3(_0336_),
    .ZN(_0378_));
 AOI22_X1 _1093_ (.A1(_0190_),
    .A2(_0369_),
    .B1(_0376_),
    .B2(_0378_),
    .ZN(_0379_));
 INV_X1 _1094_ (.A(_0379_),
    .ZN(_0039_));
 NAND2_X1 _1095_ (.A1(_0189_),
    .A2(_0370_),
    .ZN(_0380_));
 OR3_X1 _1096_ (.A1(_0187_),
    .A2(_0343_),
    .A3(_0377_),
    .ZN(_0381_));
 INV_X1 _1097_ (.A(_0190_),
    .ZN(_0382_));
 NOR3_X1 _1098_ (.A1(_0188_),
    .A2(_0189_),
    .A3(_0382_),
    .ZN(_0383_));
 NAND2_X1 _1099_ (.A1(_0376_),
    .A2(_0383_),
    .ZN(_0384_));
 OAI21_X1 _1100_ (.A(_0380_),
    .B1(_0381_),
    .B2(_0384_),
    .ZN(_0040_));
 NAND2_X1 _1101_ (.A1(_0198_),
    .A2(_0370_),
    .ZN(_0385_));
 NAND4_X1 _1102_ (.A1(_0335_),
    .A2(_0189_),
    .A3(_0382_),
    .A4(_0375_),
    .ZN(_0386_));
 OAI21_X1 _1103_ (.A(_0385_),
    .B1(_0386_),
    .B2(_0381_),
    .ZN(_0041_));
 NAND2_X1 _1104_ (.A1(_0197_),
    .A2(_0370_),
    .ZN(_0387_));
 OAI21_X1 _1105_ (.A(_0387_),
    .B1(_0374_),
    .B2(_0164_),
    .ZN(_0042_));
 NOR4_X1 _1106_ (.A1(_0218_),
    .A2(_0198_),
    .A3(_0343_),
    .A4(_0353_),
    .ZN(_0388_));
 AOI22_X1 _1107_ (.A1(_0203_),
    .A2(_0369_),
    .B1(_0376_),
    .B2(_0388_),
    .ZN(_0389_));
 INV_X1 _1108_ (.A(_0389_),
    .ZN(_0043_));
 NAND2_X1 _1109_ (.A1(_0202_),
    .A2(_0370_),
    .ZN(_0390_));
 INV_X1 _1110_ (.A(_0202_),
    .ZN(_0391_));
 NOR2_X1 _1111_ (.A1(_0343_),
    .A2(_0358_),
    .ZN(_0392_));
 NAND4_X1 _1112_ (.A1(_0391_),
    .A2(_0203_),
    .A3(_0392_),
    .A4(_0376_),
    .ZN(_0393_));
 NAND2_X1 _1113_ (.A1(_0390_),
    .A2(_0393_),
    .ZN(_0044_));
 NAND2_X1 _1114_ (.A1(\byte_controller.bit_controller.c_state[16] ),
    .A2(_0370_),
    .ZN(_0394_));
 NOR2_X1 _1115_ (.A1(_0391_),
    .A2(_0203_),
    .ZN(_0395_));
 NAND3_X1 _1116_ (.A1(_0395_),
    .A2(_0392_),
    .A3(_0376_),
    .ZN(_0396_));
 NAND2_X1 _1117_ (.A1(_0394_),
    .A2(_0396_),
    .ZN(_0045_));
 NAND2_X1 _1118_ (.A1(_0200_),
    .A2(_0370_),
    .ZN(_0397_));
 INV_X1 _1119_ (.A(_0200_),
    .ZN(_0398_));
 NOR4_X2 _1120_ (.A1(_0334_),
    .A2(_0191_),
    .A3(_0342_),
    .A4(_0343_),
    .ZN(_0399_));
 NAND4_X1 _1121_ (.A1(_0398_),
    .A2(_0201_),
    .A3(_0399_),
    .A4(_0376_),
    .ZN(_0400_));
 NAND2_X1 _1122_ (.A1(_0397_),
    .A2(_0400_),
    .ZN(_0046_));
 NAND2_X1 _1123_ (.A1(_0193_),
    .A2(_0370_),
    .ZN(_0401_));
 NOR2_X1 _1124_ (.A1(_0398_),
    .A2(_0201_),
    .ZN(_0402_));
 NAND3_X1 _1125_ (.A1(_0402_),
    .A2(_0399_),
    .A3(_0376_),
    .ZN(_0403_));
 NAND2_X1 _1126_ (.A1(_0401_),
    .A2(_0403_),
    .ZN(_0047_));
 NAND2_X1 _1127_ (.A1(_0194_),
    .A2(_0370_),
    .ZN(_0404_));
 INV_X1 _1128_ (.A(_0194_),
    .ZN(_0405_));
 NAND3_X1 _1129_ (.A1(_0193_),
    .A2(_0405_),
    .A3(_0376_),
    .ZN(_0406_));
 OAI21_X1 _1130_ (.A(_0404_),
    .B1(_0406_),
    .B2(_0366_),
    .ZN(_0048_));
 NAND2_X1 _1131_ (.A1(_0184_),
    .A2(_0369_),
    .ZN(_0407_));
 INV_X1 _1132_ (.A(_0193_),
    .ZN(_0408_));
 NAND3_X1 _1133_ (.A1(_0408_),
    .A2(_0194_),
    .A3(_0376_),
    .ZN(_0409_));
 OAI21_X1 _1134_ (.A(_0407_),
    .B1(_0409_),
    .B2(_0366_),
    .ZN(_0049_));
 NAND2_X1 _1135_ (.A1(_0185_),
    .A2(_0369_),
    .ZN(_0410_));
 OAI21_X1 _1136_ (.A(_0410_),
    .B1(_0374_),
    .B2(_0159_),
    .ZN(_0050_));
 NAND2_X1 _1137_ (.A1(_0206_),
    .A2(_0370_),
    .ZN(_0411_));
 NOR2_X1 _1138_ (.A1(_0184_),
    .A2(_0186_),
    .ZN(_0412_));
 NAND3_X1 _1139_ (.A1(_0209_),
    .A2(_0412_),
    .A3(_0376_),
    .ZN(_0413_));
 NAND2_X1 _1140_ (.A1(_0411_),
    .A2(_0413_),
    .ZN(_0051_));
 NAND2_X1 _1141_ (.A1(_0205_),
    .A2(_0369_),
    .ZN(_0414_));
 NAND3_X1 _1142_ (.A1(_0361_),
    .A2(_0206_),
    .A3(_0375_),
    .ZN(_0415_));
 OAI21_X1 _1143_ (.A(_0414_),
    .B1(_0415_),
    .B2(_0360_),
    .ZN(_0052_));
 NAND2_X1 _1144_ (.A1(_0188_),
    .A2(_0369_),
    .ZN(_0416_));
 NAND3_X1 _1145_ (.A1(_0205_),
    .A2(_0362_),
    .A3(_0375_),
    .ZN(_0417_));
 OAI21_X1 _1146_ (.A(_0416_),
    .B1(_0417_),
    .B2(_0360_),
    .ZN(_0053_));
 NAND2_X1 _1147_ (.A1(_0187_),
    .A2(_0369_),
    .ZN(_0418_));
 OAI21_X1 _1148_ (.A(_0418_),
    .B1(_0374_),
    .B2(_0171_),
    .ZN(_0054_));
 MUX2_X1 _1149_ (.A(\byte_controller.bit_controller.cmd_stop ),
    .B(\byte_controller.core_cmd[3] ),
    .S(\byte_controller.bit_controller.clk_en ),
    .Z(_0419_));
 AND2_X1 _1150_ (.A1(_0176_),
    .A2(_0419_),
    .ZN(_0055_));
 INV_X1 _1151_ (.A(\byte_controller.bit_controller.cnt[0] ),
    .ZN(_0420_));
 INV_X1 _1152_ (.A(\byte_controller.bit_controller.sSCL ),
    .ZN(_0421_));
 NAND2_X1 _1153_ (.A1(\byte_controller.bit_controller.dscl_oen ),
    .A2(_0421_),
    .ZN(_0422_));
 MUX2_X1 _1154_ (.A(_0420_),
    .B(_0035_),
    .S(_0422_),
    .Z(_0423_));
 CLKBUF_X3 _1155_ (.A(_0328_),
    .Z(_0424_));
 MUX2_X1 _1156_ (.A(\byte_controller.bit_controller.cnt[0] ),
    .B(_0423_),
    .S(_0424_),
    .Z(_0425_));
 NOR2_X1 _1157_ (.A1(_0180_),
    .A2(_0425_),
    .ZN(_0056_));
 NOR3_X1 _1158_ (.A1(\byte_controller.bit_controller.cnt[9] ),
    .A2(_0324_),
    .A3(_0323_),
    .ZN(_0426_));
 NOR3_X1 _1159_ (.A1(_0177_),
    .A2(_0424_),
    .A3(_0426_),
    .ZN(_0427_));
 AND3_X2 _1160_ (.A1(\byte_controller.bit_controller.dscl_oen ),
    .A2(_0311_),
    .A3(_0328_),
    .ZN(_0428_));
 CLKBUF_X3 _1161_ (.A(_0428_),
    .Z(_0429_));
 OAI21_X1 _1162_ (.A(\byte_controller.bit_controller.cnt[10] ),
    .B1(_0427_),
    .B2(_0429_),
    .ZN(_0430_));
 AND2_X1 _1163_ (.A1(_0307_),
    .A2(_0327_),
    .ZN(_0431_));
 NAND2_X1 _1164_ (.A1(\byte_controller.bit_controller.dscl_oen ),
    .A2(_0311_),
    .ZN(_0432_));
 BUF_X2 _1165_ (.A(_0432_),
    .Z(_0433_));
 AOI22_X1 _1166_ (.A1(\byte_controller.bit_controller.clk_cnt[10] ),
    .A2(_0433_),
    .B1(_0317_),
    .B2(_0307_),
    .ZN(_0434_));
 OR2_X1 _1167_ (.A1(_0177_),
    .A2(_0434_),
    .ZN(_0435_));
 OAI21_X1 _1168_ (.A(_0430_),
    .B1(_0431_),
    .B2(_0435_),
    .ZN(_0057_));
 OR4_X1 _1169_ (.A1(\byte_controller.bit_controller.cnt[3] ),
    .A2(_0319_),
    .A3(\byte_controller.bit_controller.cnt[0] ),
    .A4(\byte_controller.bit_controller.cnt[1] ),
    .ZN(_0436_));
 NOR2_X1 _1170_ (.A1(\byte_controller.bit_controller.cnt[4] ),
    .A2(_0436_),
    .ZN(_0437_));
 NAND2_X2 _1171_ (.A1(_0322_),
    .A2(_0437_),
    .ZN(_0438_));
 NOR2_X2 _1172_ (.A1(_0326_),
    .A2(_0438_),
    .ZN(_0439_));
 NOR3_X1 _1173_ (.A1(_0177_),
    .A2(_0424_),
    .A3(_0439_),
    .ZN(_0440_));
 OAI21_X1 _1174_ (.A(_0315_),
    .B1(_0429_),
    .B2(_0440_),
    .ZN(_0441_));
 NOR4_X1 _1175_ (.A1(_0315_),
    .A2(_0326_),
    .A3(_0328_),
    .A4(_0438_),
    .ZN(_0442_));
 AND2_X1 _1176_ (.A1(_0432_),
    .A2(_0328_),
    .ZN(_0443_));
 AOI21_X1 _1177_ (.A(_0442_),
    .B1(_0443_),
    .B2(\byte_controller.bit_controller.clk_cnt[11] ),
    .ZN(_0444_));
 CLKBUF_X3 _1178_ (.A(_0177_),
    .Z(_0445_));
 OAI21_X1 _1179_ (.A(_0441_),
    .B1(_0444_),
    .B2(_0445_),
    .ZN(_0058_));
 BUF_X2 _1180_ (.A(_0328_),
    .Z(_0446_));
 NOR4_X1 _1181_ (.A1(_0315_),
    .A2(\byte_controller.bit_controller.cnt[12] ),
    .A3(_0327_),
    .A4(_0446_),
    .ZN(_0447_));
 AND3_X1 _1182_ (.A1(\byte_controller.bit_controller.clk_cnt[12] ),
    .A2(_0433_),
    .A3(_0446_),
    .ZN(_0448_));
 OAI21_X1 _1183_ (.A(_0176_),
    .B1(_0447_),
    .B2(_0448_),
    .ZN(_0449_));
 INV_X1 _1184_ (.A(_0315_),
    .ZN(_0450_));
 NOR2_X1 _1185_ (.A1(_0323_),
    .A2(_0326_),
    .ZN(_0451_));
 NAND2_X1 _1186_ (.A1(_0450_),
    .A2(_0451_),
    .ZN(_0452_));
 AOI21_X1 _1187_ (.A(_0429_),
    .B1(_0452_),
    .B2(_0330_),
    .ZN(_0453_));
 INV_X1 _1188_ (.A(\byte_controller.bit_controller.cnt[12] ),
    .ZN(_0454_));
 OAI21_X1 _1189_ (.A(_0449_),
    .B1(_0453_),
    .B2(_0454_),
    .ZN(_0059_));
 NAND2_X1 _1190_ (.A1(_0316_),
    .A2(_0439_),
    .ZN(_0455_));
 NAND2_X1 _1191_ (.A1(\byte_controller.bit_controller.clk_cnt[13] ),
    .A2(_0433_),
    .ZN(_0456_));
 MUX2_X1 _1192_ (.A(_0455_),
    .B(_0456_),
    .S(_0424_),
    .Z(_0457_));
 NAND3_X1 _1193_ (.A1(_0450_),
    .A2(_0454_),
    .A3(_0439_),
    .ZN(_0458_));
 AOI21_X1 _1194_ (.A(_0429_),
    .B1(_0458_),
    .B2(_0330_),
    .ZN(_0459_));
 INV_X1 _1195_ (.A(\byte_controller.bit_controller.cnt[13] ),
    .ZN(_0460_));
 OAI22_X1 _1196_ (.A1(_0180_),
    .A2(_0457_),
    .B1(_0459_),
    .B2(_0460_),
    .ZN(_0060_));
 NAND2_X1 _1197_ (.A1(_0314_),
    .A2(_0316_),
    .ZN(_0461_));
 NOR3_X1 _1198_ (.A1(_0461_),
    .A2(_0327_),
    .A3(_0424_),
    .ZN(_0462_));
 AND3_X1 _1199_ (.A1(\byte_controller.bit_controller.clk_cnt[14] ),
    .A2(_0433_),
    .A3(_0446_),
    .ZN(_0463_));
 OAI21_X1 _1200_ (.A(_0176_),
    .B1(_0462_),
    .B2(_0463_),
    .ZN(_0464_));
 NAND2_X1 _1201_ (.A1(_0316_),
    .A2(_0451_),
    .ZN(_0465_));
 AOI21_X1 _1202_ (.A(_0429_),
    .B1(_0465_),
    .B2(_0330_),
    .ZN(_0466_));
 OAI21_X1 _1203_ (.A(_0464_),
    .B1(_0466_),
    .B2(_0314_),
    .ZN(_0061_));
 OR3_X1 _1204_ (.A1(_0317_),
    .A2(_0326_),
    .A3(_0438_),
    .ZN(_0467_));
 NAND2_X1 _1205_ (.A1(\byte_controller.bit_controller.clk_cnt[15] ),
    .A2(_0433_),
    .ZN(_0468_));
 MUX2_X1 _1206_ (.A(_0467_),
    .B(_0468_),
    .S(_0424_),
    .Z(_0469_));
 NAND3_X1 _1207_ (.A1(_0314_),
    .A2(_0316_),
    .A3(_0439_),
    .ZN(_0470_));
 AOI21_X1 _1208_ (.A(_0428_),
    .B1(_0470_),
    .B2(_0330_),
    .ZN(_0471_));
 OAI22_X1 _1209_ (.A1(_0180_),
    .A2(_0469_),
    .B1(_0471_),
    .B2(_0313_),
    .ZN(_0062_));
 NAND2_X1 _1210_ (.A1(\byte_controller.bit_controller.cnt[1] ),
    .A2(_0429_),
    .ZN(_0472_));
 NOR2_X1 _1211_ (.A1(_0793_),
    .A2(_0424_),
    .ZN(_0473_));
 AOI21_X1 _1212_ (.A(_0473_),
    .B1(_0443_),
    .B2(\byte_controller.bit_controller.clk_cnt[1] ),
    .ZN(_0474_));
 OAI21_X1 _1213_ (.A(_0472_),
    .B1(_0474_),
    .B2(_0445_),
    .ZN(_0063_));
 INV_X1 _1214_ (.A(_0792_),
    .ZN(_0475_));
 NOR3_X1 _1215_ (.A1(_0319_),
    .A2(_0475_),
    .A3(_0446_),
    .ZN(_0476_));
 AOI21_X1 _1216_ (.A(_0476_),
    .B1(_0443_),
    .B2(\byte_controller.bit_controller.clk_cnt[2] ),
    .ZN(_0477_));
 AOI21_X1 _1217_ (.A(_0428_),
    .B1(_0330_),
    .B2(_0475_),
    .ZN(_0478_));
 INV_X1 _1218_ (.A(_0319_),
    .ZN(_0479_));
 OAI22_X1 _1219_ (.A1(_0180_),
    .A2(_0477_),
    .B1(_0478_),
    .B2(_0479_),
    .ZN(_0064_));
 NOR3_X1 _1220_ (.A1(_0319_),
    .A2(\byte_controller.bit_controller.cnt[0] ),
    .A3(\byte_controller.bit_controller.cnt[1] ),
    .ZN(_0480_));
 NOR3_X1 _1221_ (.A1(_0177_),
    .A2(_0424_),
    .A3(_0480_),
    .ZN(_0481_));
 OAI21_X1 _1222_ (.A(\byte_controller.bit_controller.cnt[3] ),
    .B1(_0429_),
    .B2(_0481_),
    .ZN(_0482_));
 NAND2_X1 _1223_ (.A1(\byte_controller.bit_controller.clk_cnt[3] ),
    .A2(_0433_),
    .ZN(_0483_));
 MUX2_X1 _1224_ (.A(_0436_),
    .B(_0483_),
    .S(_0424_),
    .Z(_0484_));
 OAI21_X1 _1225_ (.A(_0482_),
    .B1(_0484_),
    .B2(_0445_),
    .ZN(_0065_));
 NAND3_X1 _1226_ (.A1(_0792_),
    .A2(_0318_),
    .A3(_0320_),
    .ZN(_0485_));
 NAND2_X1 _1227_ (.A1(\byte_controller.bit_controller.clk_cnt[4] ),
    .A2(_0433_),
    .ZN(_0486_));
 MUX2_X1 _1228_ (.A(_0485_),
    .B(_0486_),
    .S(_0424_),
    .Z(_0487_));
 NAND2_X1 _1229_ (.A1(_0792_),
    .A2(_0320_),
    .ZN(_0488_));
 AOI21_X1 _1230_ (.A(_0428_),
    .B1(_0330_),
    .B2(_0488_),
    .ZN(_0489_));
 OAI22_X1 _1231_ (.A1(_0180_),
    .A2(_0487_),
    .B1(_0489_),
    .B2(_0318_),
    .ZN(_0066_));
 OR2_X1 _1232_ (.A1(\byte_controller.bit_controller.cnt[4] ),
    .A2(_0436_),
    .ZN(_0490_));
 NOR3_X1 _1233_ (.A1(_0321_),
    .A2(_0446_),
    .A3(_0490_),
    .ZN(_0491_));
 AOI21_X1 _1234_ (.A(_0491_),
    .B1(_0443_),
    .B2(\byte_controller.bit_controller.clk_cnt[5] ),
    .ZN(_0492_));
 AOI21_X1 _1235_ (.A(_0428_),
    .B1(_0490_),
    .B2(_0330_),
    .ZN(_0493_));
 INV_X1 _1236_ (.A(_0321_),
    .ZN(_0494_));
 OAI22_X1 _1237_ (.A1(_0180_),
    .A2(_0492_),
    .B1(_0493_),
    .B2(_0494_),
    .ZN(_0067_));
 NOR4_X1 _1238_ (.A1(_0321_),
    .A2(\byte_controller.bit_controller.cnt[6] ),
    .A3(_0485_),
    .A4(_0446_),
    .ZN(_0495_));
 AND3_X1 _1239_ (.A1(\byte_controller.bit_controller.clk_cnt[6] ),
    .A2(_0433_),
    .A3(_0446_),
    .ZN(_0496_));
 OAI21_X1 _1240_ (.A(_0176_),
    .B1(_0495_),
    .B2(_0496_),
    .ZN(_0497_));
 OR2_X1 _1241_ (.A1(_0321_),
    .A2(_0485_),
    .ZN(_0498_));
 AOI21_X1 _1242_ (.A(_0429_),
    .B1(_0498_),
    .B2(_0330_),
    .ZN(_0499_));
 INV_X1 _1243_ (.A(\byte_controller.bit_controller.cnt[6] ),
    .ZN(_0500_));
 OAI21_X1 _1244_ (.A(_0497_),
    .B1(_0499_),
    .B2(_0500_),
    .ZN(_0068_));
 NAND2_X1 _1245_ (.A1(\byte_controller.bit_controller.clk_cnt[7] ),
    .A2(_0433_),
    .ZN(_0501_));
 MUX2_X1 _1246_ (.A(_0438_),
    .B(_0501_),
    .S(_0446_),
    .Z(_0502_));
 NAND3_X1 _1247_ (.A1(_0494_),
    .A2(_0500_),
    .A3(_0437_),
    .ZN(_0503_));
 AOI21_X1 _1248_ (.A(_0428_),
    .B1(_0503_),
    .B2(_0329_),
    .ZN(_0504_));
 INV_X1 _1249_ (.A(\byte_controller.bit_controller.cnt[7] ),
    .ZN(_0505_));
 OAI22_X1 _1250_ (.A1(_0180_),
    .A2(_0502_),
    .B1(_0504_),
    .B2(_0505_),
    .ZN(_0069_));
 NAND2_X1 _1251_ (.A1(_0324_),
    .A2(_0429_),
    .ZN(_0506_));
 NOR3_X1 _1252_ (.A1(_0324_),
    .A2(_0323_),
    .A3(_0328_),
    .ZN(_0507_));
 AND2_X1 _1253_ (.A1(_0307_),
    .A2(_0323_),
    .ZN(_0508_));
 AOI221_X1 _1254_ (.A(_0507_),
    .B1(_0508_),
    .B2(_0324_),
    .C1(\byte_controller.bit_controller.clk_cnt[8] ),
    .C2(_0443_),
    .ZN(_0509_));
 OAI21_X1 _1255_ (.A(_0506_),
    .B1(_0509_),
    .B2(_0445_),
    .ZN(_0070_));
 NOR4_X1 _1256_ (.A1(\byte_controller.bit_controller.cnt[9] ),
    .A2(_0324_),
    .A3(_0446_),
    .A4(_0438_),
    .ZN(_0510_));
 AND3_X1 _1257_ (.A1(\byte_controller.bit_controller.clk_cnt[9] ),
    .A2(_0433_),
    .A3(_0446_),
    .ZN(_0511_));
 OAI21_X1 _1258_ (.A(_0176_),
    .B1(_0510_),
    .B2(_0511_),
    .ZN(_0512_));
 OR2_X1 _1259_ (.A1(_0324_),
    .A2(_0438_),
    .ZN(_0513_));
 AOI21_X1 _1260_ (.A(_0429_),
    .B1(_0513_),
    .B2(_0330_),
    .ZN(_0514_));
 INV_X1 _1261_ (.A(\byte_controller.bit_controller.cnt[9] ),
    .ZN(_0515_));
 OAI21_X1 _1262_ (.A(_0512_),
    .B1(_0514_),
    .B2(_0515_),
    .ZN(_0071_));
 NOR2_X1 _1263_ (.A1(_0421_),
    .A2(\byte_controller.bit_controller.dSCL ),
    .ZN(_0516_));
 MUX2_X1 _1264_ (.A(\byte_controller.bit_controller.dout ),
    .B(\byte_controller.bit_controller.sSDA ),
    .S(_0516_),
    .Z(_0072_));
 OAI21_X1 _1265_ (.A(_0333_),
    .B1(_0355_),
    .B2(_0378_),
    .ZN(_0517_));
 NOR2_X1 _1266_ (.A1(_0129_),
    .A2(_0517_),
    .ZN(_0518_));
 NOR2_X1 _1267_ (.A1(net9),
    .A2(_0129_),
    .ZN(_0519_));
 OAI21_X1 _1268_ (.A(_0338_),
    .B1(_0339_),
    .B2(_0188_),
    .ZN(_0520_));
 XNOR2_X1 _1269_ (.A(_0205_),
    .B(_0206_),
    .ZN(_0521_));
 OAI22_X1 _1270_ (.A1(_0520_),
    .A2(_0381_),
    .B1(_0521_),
    .B2(_0360_),
    .ZN(_0522_));
 OR2_X1 _1271_ (.A1(_0366_),
    .A2(_0364_),
    .ZN(_0523_));
 NAND2_X1 _1272_ (.A1(_0402_),
    .A2(_0399_),
    .ZN(_0524_));
 NAND3_X1 _1273_ (.A1(_0523_),
    .A2(_0359_),
    .A3(_0524_),
    .ZN(_0525_));
 OAI21_X1 _1274_ (.A(_0333_),
    .B1(_0522_),
    .B2(_0525_),
    .ZN(_0526_));
 AOI21_X1 _1275_ (.A(_0518_),
    .B1(_0519_),
    .B2(_0526_),
    .ZN(_0073_));
 NOR4_X2 _1276_ (.A1(_0212_),
    .A2(_0357_),
    .A3(_0343_),
    .A4(_0356_),
    .ZN(_0527_));
 AOI21_X1 _1277_ (.A(\byte_controller.bit_controller.sda_chk ),
    .B1(_0372_),
    .B2(_0527_),
    .ZN(_0528_));
 NOR2_X1 _1278_ (.A1(_0360_),
    .A2(_0521_),
    .ZN(_0529_));
 AOI21_X1 _1279_ (.A(_0366_),
    .B1(_0194_),
    .B2(_0193_),
    .ZN(_0530_));
 OR4_X1 _1280_ (.A1(_0346_),
    .A2(_0355_),
    .A3(_0529_),
    .A4(_0530_),
    .ZN(_0531_));
 AOI21_X1 _1281_ (.A(_0528_),
    .B1(_0531_),
    .B2(_0372_),
    .ZN(_0074_));
 OR2_X1 _1282_ (.A1(_0220_),
    .A2(_0346_),
    .ZN(_0532_));
 INV_X1 _1283_ (.A(\byte_controller.bit_controller.din ),
    .ZN(_0533_));
 NOR4_X2 _1284_ (.A1(_0218_),
    .A2(_0198_),
    .A3(_0191_),
    .A4(_0217_),
    .ZN(_0534_));
 NOR3_X1 _1285_ (.A1(_0216_),
    .A2(_0527_),
    .A3(_0534_),
    .ZN(_0535_));
 NOR2_X1 _1286_ (.A1(_0533_),
    .A2(_0535_),
    .ZN(_0536_));
 OAI21_X1 _1287_ (.A(_0372_),
    .B1(_0532_),
    .B2(_0536_),
    .ZN(_0537_));
 NOR2_X1 _1288_ (.A1(_0366_),
    .A2(_0364_),
    .ZN(_0538_));
 NOR3_X1 _1289_ (.A1(_0538_),
    .A2(_0527_),
    .A3(_0529_),
    .ZN(_0539_));
 NOR3_X1 _1290_ (.A1(_0216_),
    .A2(_0348_),
    .A3(_0534_),
    .ZN(_0540_));
 AOI21_X1 _1291_ (.A(_0031_),
    .B1(_0539_),
    .B2(_0540_),
    .ZN(_0541_));
 NOR2_X1 _1292_ (.A1(_0532_),
    .A2(_0536_),
    .ZN(_0542_));
 AOI22_X1 _1293_ (.A1(_0230_),
    .A2(_0537_),
    .B1(_0541_),
    .B2(_0542_),
    .ZN(_0075_));
 CLKBUF_X3 _1294_ (.A(\byte_controller.ld ),
    .Z(_0543_));
 INV_X2 _1295_ (.A(_0543_),
    .ZN(_0544_));
 CLKBUF_X3 _1296_ (.A(\byte_controller.shift ),
    .Z(_0545_));
 XNOR2_X1 _1297_ (.A(_0545_),
    .B(\byte_controller.dcnt[0] ),
    .ZN(_0546_));
 AOI21_X1 _1298_ (.A(_0445_),
    .B1(_0544_),
    .B2(_0546_),
    .ZN(_0076_));
 NOR2_X2 _1299_ (.A1(_0545_),
    .A2(_0543_),
    .ZN(_0547_));
 AOI21_X1 _1300_ (.A(_0547_),
    .B1(_0797_),
    .B2(_0036_),
    .ZN(_0548_));
 AOI21_X1 _1301_ (.A(_0548_),
    .B1(_0547_),
    .B2(\byte_controller.dcnt[1] ),
    .ZN(_0549_));
 NOR2_X1 _1302_ (.A1(_0180_),
    .A2(_0549_),
    .ZN(_0077_));
 INV_X1 _1303_ (.A(_0547_),
    .ZN(_0550_));
 NAND3_X1 _1304_ (.A1(\byte_controller.dcnt[2] ),
    .A2(_0798_),
    .A3(_0550_),
    .ZN(_0551_));
 OAI21_X1 _1305_ (.A(_0551_),
    .B1(_0798_),
    .B2(\byte_controller.dcnt[2] ),
    .ZN(_0552_));
 AOI221_X1 _1306_ (.A(_0146_),
    .B1(_0160_),
    .B2(_0547_),
    .C1(_0552_),
    .C2(_0036_),
    .ZN(_0078_));
 NOR2_X1 _1307_ (.A1(_0544_),
    .A2(\byte_controller.din[0] ),
    .ZN(_0553_));
 MUX2_X1 _1308_ (.A(\byte_controller.dout[0] ),
    .B(\byte_controller.bit_controller.dout ),
    .S(_0545_),
    .Z(_0554_));
 NOR2_X1 _1309_ (.A1(_0543_),
    .A2(_0554_),
    .ZN(_0555_));
 NOR3_X1 _1310_ (.A1(_0178_),
    .A2(_0553_),
    .A3(_0555_),
    .ZN(_0079_));
 NOR2_X1 _1311_ (.A1(_0544_),
    .A2(\byte_controller.din[1] ),
    .ZN(_0556_));
 MUX2_X1 _1312_ (.A(\byte_controller.dout[1] ),
    .B(\byte_controller.dout[0] ),
    .S(_0545_),
    .Z(_0557_));
 NOR2_X1 _1313_ (.A1(_0543_),
    .A2(_0557_),
    .ZN(_0558_));
 NOR3_X1 _1314_ (.A1(_0178_),
    .A2(_0556_),
    .A3(_0558_),
    .ZN(_0080_));
 NOR2_X1 _1315_ (.A1(_0544_),
    .A2(\byte_controller.din[2] ),
    .ZN(_0559_));
 MUX2_X1 _1316_ (.A(\byte_controller.dout[2] ),
    .B(\byte_controller.dout[1] ),
    .S(_0545_),
    .Z(_0560_));
 NOR2_X1 _1317_ (.A1(_0543_),
    .A2(_0560_),
    .ZN(_0561_));
 NOR3_X1 _1318_ (.A1(_0178_),
    .A2(_0559_),
    .A3(_0561_),
    .ZN(_0081_));
 NOR2_X1 _1319_ (.A1(_0544_),
    .A2(\byte_controller.din[3] ),
    .ZN(_0562_));
 MUX2_X1 _1320_ (.A(\byte_controller.dout[3] ),
    .B(\byte_controller.dout[2] ),
    .S(_0545_),
    .Z(_0563_));
 NOR2_X1 _1321_ (.A1(_0543_),
    .A2(_0563_),
    .ZN(_0564_));
 NOR3_X1 _1322_ (.A1(_0178_),
    .A2(_0562_),
    .A3(_0564_),
    .ZN(_0082_));
 NOR2_X1 _1323_ (.A1(_0544_),
    .A2(\byte_controller.din[4] ),
    .ZN(_0565_));
 MUX2_X1 _1324_ (.A(\byte_controller.dout[4] ),
    .B(\byte_controller.dout[3] ),
    .S(_0545_),
    .Z(_0566_));
 NOR2_X1 _1325_ (.A1(_0543_),
    .A2(_0566_),
    .ZN(_0567_));
 NOR3_X1 _1326_ (.A1(_0178_),
    .A2(_0565_),
    .A3(_0567_),
    .ZN(_0083_));
 NOR2_X1 _1327_ (.A1(_0544_),
    .A2(\byte_controller.din[5] ),
    .ZN(_0568_));
 MUX2_X1 _1328_ (.A(\byte_controller.dout[5] ),
    .B(\byte_controller.dout[4] ),
    .S(_0545_),
    .Z(_0569_));
 NOR2_X1 _1329_ (.A1(_0543_),
    .A2(_0569_),
    .ZN(_0570_));
 NOR3_X1 _1330_ (.A1(_0178_),
    .A2(_0568_),
    .A3(_0570_),
    .ZN(_0084_));
 NOR2_X1 _1331_ (.A1(_0544_),
    .A2(\byte_controller.din[6] ),
    .ZN(_0571_));
 MUX2_X1 _1332_ (.A(\byte_controller.dout[6] ),
    .B(\byte_controller.dout[5] ),
    .S(_0545_),
    .Z(_0572_));
 NOR2_X1 _1333_ (.A1(_0543_),
    .A2(_0572_),
    .ZN(_0573_));
 NOR3_X1 _1334_ (.A1(_0178_),
    .A2(_0571_),
    .A3(_0573_),
    .ZN(_0085_));
 NOR2_X1 _1335_ (.A1(_0544_),
    .A2(\byte_controller.din[7] ),
    .ZN(_0574_));
 MUX2_X1 _1336_ (.A(_0234_),
    .B(\byte_controller.dout[6] ),
    .S(_0545_),
    .Z(_0575_));
 NOR2_X1 _1337_ (.A1(_0543_),
    .A2(_0575_),
    .ZN(_0576_));
 NOR3_X1 _1338_ (.A1(_0178_),
    .A2(_0574_),
    .A3(_0576_),
    .ZN(_0086_));
 NAND3_X4 _1339_ (.A1(net7),
    .A2(net5),
    .A3(net8),
    .ZN(_0577_));
 NOR2_X4 _1340_ (.A1(_0146_),
    .A2(_0577_),
    .ZN(_0578_));
 BUF_X1 _1341_ (.A(wb_dat_i[0]),
    .Z(_0579_));
 NAND2_X1 _1342_ (.A1(_0245_),
    .A2(_0307_),
    .ZN(_0580_));
 NOR2_X1 _1343_ (.A1(_0261_),
    .A2(_0580_),
    .ZN(_0581_));
 MUX2_X1 _1344_ (.A(\cr[0] ),
    .B(_0579_),
    .S(_0581_),
    .Z(_0582_));
 AND2_X1 _1345_ (.A1(_0578_),
    .A2(_0582_),
    .ZN(_0087_));
 BUF_X1 _1346_ (.A(wb_dat_i[1]),
    .Z(_0583_));
 MUX2_X1 _1347_ (.A(\cr[1] ),
    .B(_0583_),
    .S(_0581_),
    .Z(_0584_));
 AND2_X1 _1348_ (.A1(_0578_),
    .A2(_0584_),
    .ZN(_0088_));
 BUF_X1 _1349_ (.A(wb_dat_i[2]),
    .Z(_0585_));
 MUX2_X1 _1350_ (.A(\cr[2] ),
    .B(_0585_),
    .S(_0581_),
    .Z(_0586_));
 AND2_X1 _1351_ (.A1(_0578_),
    .A2(_0586_),
    .ZN(_0089_));
 CLKBUF_X2 _1352_ (.A(wb_dat_i[3]),
    .Z(_0587_));
 NOR3_X4 _1353_ (.A1(_0261_),
    .A2(_0577_),
    .A3(_0580_),
    .ZN(_0588_));
 MUX2_X1 _1354_ (.A(_0233_),
    .B(_0587_),
    .S(_0588_),
    .Z(_0589_));
 AND2_X1 _1355_ (.A1(_0176_),
    .A2(_0589_),
    .ZN(_0090_));
 OAI21_X1 _1356_ (.A(_0577_),
    .B1(\byte_controller.cmd_ack ),
    .B2(_0127_),
    .ZN(_0590_));
 INV_X1 _1357_ (.A(_0590_),
    .ZN(_0591_));
 NOR3_X4 _1358_ (.A1(_0146_),
    .A2(_0588_),
    .A3(_0591_),
    .ZN(_0592_));
 NAND2_X1 _1359_ (.A1(\byte_controller.write ),
    .A2(_0592_),
    .ZN(_0593_));
 BUF_X2 _1360_ (.A(wb_dat_i[4]),
    .Z(_0594_));
 NAND2_X1 _1361_ (.A1(_0594_),
    .A2(_0578_),
    .ZN(_0595_));
 OAI21_X1 _1362_ (.A(_0593_),
    .B1(_0595_),
    .B2(_0592_),
    .ZN(_0091_));
 NAND2_X1 _1363_ (.A1(_0131_),
    .A2(_0592_),
    .ZN(_0596_));
 CLKBUF_X2 _1364_ (.A(wb_dat_i[5]),
    .Z(_0597_));
 NAND2_X1 _1365_ (.A1(_0597_),
    .A2(_0578_),
    .ZN(_0598_));
 OAI21_X1 _1366_ (.A(_0596_),
    .B1(_0598_),
    .B2(_0592_),
    .ZN(_0092_));
 NAND2_X1 _1367_ (.A1(\byte_controller.stop ),
    .A2(_0592_),
    .ZN(_0599_));
 CLKBUF_X2 _1368_ (.A(wb_dat_i[6]),
    .Z(_0600_));
 NAND2_X1 _1369_ (.A1(_0600_),
    .A2(_0578_),
    .ZN(_0601_));
 OAI21_X1 _1370_ (.A(_0599_),
    .B1(_0601_),
    .B2(_0592_),
    .ZN(_0093_));
 NAND2_X1 _1371_ (.A1(_0130_),
    .A2(_0592_),
    .ZN(_0602_));
 BUF_X1 _1372_ (.A(wb_dat_i[7]),
    .Z(_0603_));
 NAND2_X1 _1373_ (.A1(_0603_),
    .A2(_0578_),
    .ZN(_0604_));
 OAI21_X1 _1374_ (.A(_0602_),
    .B1(_0604_),
    .B2(_0592_),
    .ZN(_0094_));
 NOR2_X4 _1375_ (.A1(_0245_),
    .A2(_0577_),
    .ZN(_0605_));
 AND2_X1 _1376_ (.A1(_0259_),
    .A2(_0605_),
    .ZN(_0606_));
 BUF_X2 _1377_ (.A(_0606_),
    .Z(_0607_));
 NAND2_X1 _1378_ (.A1(_0579_),
    .A2(_0607_),
    .ZN(_0608_));
 NAND2_X2 _1379_ (.A1(_0259_),
    .A2(_0605_),
    .ZN(_0609_));
 NAND2_X1 _1380_ (.A1(\ctr[0] ),
    .A2(_0609_),
    .ZN(_0610_));
 AOI21_X1 _1381_ (.A(_0445_),
    .B1(_0608_),
    .B2(_0610_),
    .ZN(_0095_));
 NAND2_X1 _1382_ (.A1(_0583_),
    .A2(_0607_),
    .ZN(_0611_));
 NAND2_X1 _1383_ (.A1(\ctr[1] ),
    .A2(_0609_),
    .ZN(_0612_));
 AOI21_X1 _1384_ (.A(_0445_),
    .B1(_0611_),
    .B2(_0612_),
    .ZN(_0096_));
 NAND2_X1 _1385_ (.A1(_0585_),
    .A2(_0607_),
    .ZN(_0613_));
 NAND2_X1 _1386_ (.A1(\ctr[2] ),
    .A2(_0609_),
    .ZN(_0614_));
 AOI21_X1 _1387_ (.A(_0445_),
    .B1(_0613_),
    .B2(_0614_),
    .ZN(_0097_));
 NAND2_X1 _1388_ (.A1(_0587_),
    .A2(_0607_),
    .ZN(_0615_));
 NAND2_X1 _1389_ (.A1(\ctr[3] ),
    .A2(_0609_),
    .ZN(_0616_));
 AOI21_X1 _1390_ (.A(_0445_),
    .B1(_0615_),
    .B2(_0616_),
    .ZN(_0098_));
 NAND2_X1 _1391_ (.A1(_0594_),
    .A2(_0607_),
    .ZN(_0617_));
 NAND2_X1 _1392_ (.A1(\ctr[4] ),
    .A2(_0609_),
    .ZN(_0618_));
 AOI21_X1 _1393_ (.A(_0445_),
    .B1(_0617_),
    .B2(_0618_),
    .ZN(_0099_));
 CLKBUF_X3 _1394_ (.A(_0177_),
    .Z(_0619_));
 NAND2_X1 _1395_ (.A1(_0597_),
    .A2(_0607_),
    .ZN(_0620_));
 NAND2_X1 _1396_ (.A1(\ctr[5] ),
    .A2(_0609_),
    .ZN(_0621_));
 AOI21_X1 _1397_ (.A(_0619_),
    .B1(_0620_),
    .B2(_0621_),
    .ZN(_0100_));
 NAND2_X1 _1398_ (.A1(_0600_),
    .A2(_0607_),
    .ZN(_0622_));
 NAND2_X1 _1399_ (.A1(\ctr[6] ),
    .A2(_0609_),
    .ZN(_0623_));
 AOI21_X1 _1400_ (.A(_0619_),
    .B1(_0622_),
    .B2(_0623_),
    .ZN(_0101_));
 NAND2_X1 _1401_ (.A1(_0603_),
    .A2(_0607_),
    .ZN(_0624_));
 NAND2_X1 _1402_ (.A1(_0307_),
    .A2(_0609_),
    .ZN(_0625_));
 AOI21_X1 _1403_ (.A(_0619_),
    .B1(_0624_),
    .B2(_0625_),
    .ZN(_0102_));
 NOR3_X4 _1404_ (.A1(_0245_),
    .A2(_0261_),
    .A3(_0577_),
    .ZN(_0626_));
 MUX2_X1 _1405_ (.A(\byte_controller.bit_controller.clk_cnt[0] ),
    .B(_0579_),
    .S(_0626_),
    .Z(_0627_));
 OR2_X1 _1406_ (.A1(_0312_),
    .A2(_0627_),
    .ZN(_0103_));
 NAND2_X1 _1407_ (.A1(_0258_),
    .A2(_0605_),
    .ZN(_0628_));
 NAND2_X2 _1408_ (.A1(_0176_),
    .A2(_0628_),
    .ZN(_0629_));
 NAND3_X4 _1409_ (.A1(_0263_),
    .A2(_0258_),
    .A3(_0578_),
    .ZN(_0630_));
 OAI22_X1 _1410_ (.A1(\byte_controller.bit_controller.clk_cnt[10] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0585_),
    .ZN(_0631_));
 INV_X1 _1411_ (.A(_0631_),
    .ZN(_0104_));
 OAI22_X1 _1412_ (.A1(\byte_controller.bit_controller.clk_cnt[11] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0587_),
    .ZN(_0632_));
 INV_X1 _1413_ (.A(_0632_),
    .ZN(_0105_));
 OAI22_X1 _1414_ (.A1(\byte_controller.bit_controller.clk_cnt[12] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0594_),
    .ZN(_0633_));
 INV_X1 _1415_ (.A(_0633_),
    .ZN(_0106_));
 OAI22_X1 _1416_ (.A1(\byte_controller.bit_controller.clk_cnt[13] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0597_),
    .ZN(_0634_));
 INV_X1 _1417_ (.A(_0634_),
    .ZN(_0107_));
 OAI22_X1 _1418_ (.A1(\byte_controller.bit_controller.clk_cnt[14] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0600_),
    .ZN(_0635_));
 INV_X1 _1419_ (.A(_0635_),
    .ZN(_0108_));
 OAI22_X1 _1420_ (.A1(\byte_controller.bit_controller.clk_cnt[15] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0603_),
    .ZN(_0636_));
 INV_X1 _1421_ (.A(_0636_),
    .ZN(_0109_));
 MUX2_X1 _1422_ (.A(\byte_controller.bit_controller.clk_cnt[1] ),
    .B(_0583_),
    .S(_0626_),
    .Z(_0637_));
 OR2_X1 _1423_ (.A1(_0312_),
    .A2(_0637_),
    .ZN(_0110_));
 MUX2_X1 _1424_ (.A(\byte_controller.bit_controller.clk_cnt[2] ),
    .B(_0585_),
    .S(_0626_),
    .Z(_0638_));
 OR2_X1 _1425_ (.A1(_0312_),
    .A2(_0638_),
    .ZN(_0111_));
 MUX2_X1 _1426_ (.A(\byte_controller.bit_controller.clk_cnt[3] ),
    .B(_0587_),
    .S(_0626_),
    .Z(_0639_));
 OR2_X1 _1427_ (.A1(_0312_),
    .A2(_0639_),
    .ZN(_0112_));
 MUX2_X1 _1428_ (.A(\byte_controller.bit_controller.clk_cnt[4] ),
    .B(_0594_),
    .S(_0626_),
    .Z(_0640_));
 OR2_X1 _1429_ (.A1(_0312_),
    .A2(_0640_),
    .ZN(_0113_));
 MUX2_X1 _1430_ (.A(\byte_controller.bit_controller.clk_cnt[5] ),
    .B(_0597_),
    .S(_0626_),
    .Z(_0641_));
 OR2_X1 _1431_ (.A1(_0312_),
    .A2(_0641_),
    .ZN(_0114_));
 MUX2_X1 _1432_ (.A(\byte_controller.bit_controller.clk_cnt[6] ),
    .B(_0600_),
    .S(_0626_),
    .Z(_0642_));
 OR2_X1 _1433_ (.A1(_0312_),
    .A2(_0642_),
    .ZN(_0115_));
 MUX2_X1 _1434_ (.A(\byte_controller.bit_controller.clk_cnt[7] ),
    .B(_0603_),
    .S(_0626_),
    .Z(_0643_));
 OR2_X1 _1435_ (.A1(_0177_),
    .A2(_0643_),
    .ZN(_0116_));
 OAI22_X1 _1436_ (.A1(\byte_controller.bit_controller.clk_cnt[8] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0579_),
    .ZN(_0644_));
 INV_X1 _1437_ (.A(_0644_),
    .ZN(_0117_));
 OAI22_X1 _1438_ (.A1(\byte_controller.bit_controller.clk_cnt[9] ),
    .A2(_0629_),
    .B1(_0630_),
    .B2(_0583_),
    .ZN(_0645_));
 INV_X1 _1439_ (.A(_0645_),
    .ZN(_0118_));
 NOR4_X4 _1440_ (.A1(_0245_),
    .A2(_0254_),
    .A3(_0247_),
    .A4(_0577_),
    .ZN(_0646_));
 NAND2_X1 _1441_ (.A1(_0579_),
    .A2(_0646_),
    .ZN(_0647_));
 NAND3_X4 _1442_ (.A1(_0265_),
    .A2(_0256_),
    .A3(_0605_),
    .ZN(_0648_));
 NAND2_X1 _1443_ (.A1(\byte_controller.din[0] ),
    .A2(_0648_),
    .ZN(_0649_));
 AOI21_X1 _1444_ (.A(_0619_),
    .B1(_0647_),
    .B2(_0649_),
    .ZN(_0119_));
 NAND2_X1 _1445_ (.A1(_0583_),
    .A2(_0646_),
    .ZN(_0650_));
 NAND2_X1 _1446_ (.A1(\byte_controller.din[1] ),
    .A2(_0648_),
    .ZN(_0651_));
 AOI21_X1 _1447_ (.A(_0619_),
    .B1(_0650_),
    .B2(_0651_),
    .ZN(_0120_));
 NAND2_X1 _1448_ (.A1(_0585_),
    .A2(_0646_),
    .ZN(_0652_));
 NAND2_X1 _1449_ (.A1(\byte_controller.din[2] ),
    .A2(_0648_),
    .ZN(_0653_));
 AOI21_X1 _1450_ (.A(_0619_),
    .B1(_0652_),
    .B2(_0653_),
    .ZN(_0121_));
 NAND2_X1 _1451_ (.A1(_0587_),
    .A2(_0646_),
    .ZN(_0654_));
 NAND2_X1 _1452_ (.A1(\byte_controller.din[3] ),
    .A2(_0648_),
    .ZN(_0655_));
 AOI21_X1 _1453_ (.A(_0619_),
    .B1(_0654_),
    .B2(_0655_),
    .ZN(_0122_));
 NAND2_X1 _1454_ (.A1(_0594_),
    .A2(_0646_),
    .ZN(_0656_));
 NAND2_X1 _1455_ (.A1(\byte_controller.din[4] ),
    .A2(_0648_),
    .ZN(_0657_));
 AOI21_X1 _1456_ (.A(_0619_),
    .B1(_0656_),
    .B2(_0657_),
    .ZN(_0123_));
 NAND2_X1 _1457_ (.A1(_0597_),
    .A2(_0646_),
    .ZN(_0658_));
 NAND2_X1 _1458_ (.A1(\byte_controller.din[5] ),
    .A2(_0648_),
    .ZN(_0659_));
 AOI21_X1 _1459_ (.A(_0619_),
    .B1(_0658_),
    .B2(_0659_),
    .ZN(_0124_));
 NAND2_X1 _1460_ (.A1(_0600_),
    .A2(_0646_),
    .ZN(_0660_));
 NAND2_X1 _1461_ (.A1(\byte_controller.din[6] ),
    .A2(_0648_),
    .ZN(_0661_));
 AOI21_X1 _1462_ (.A(_0619_),
    .B1(_0660_),
    .B2(_0661_),
    .ZN(_0125_));
 NAND2_X1 _1463_ (.A1(_0603_),
    .A2(_0646_),
    .ZN(_0662_));
 NAND2_X1 _1464_ (.A1(\byte_controller.din[7] ),
    .A2(_0648_),
    .ZN(_0663_));
 AOI21_X1 _1465_ (.A(_0312_),
    .B1(_0662_),
    .B2(_0663_),
    .ZN(_0126_));
 HA_X1 _1466_ (.A(_0790_),
    .B(_0791_),
    .CO(_0792_),
    .S(_0793_));
 HA_X1 _1467_ (.A(_0794_),
    .B(_0795_),
    .CO(_0796_),
    .S(_0797_));
 HA_X1 _1468_ (.A(_0794_),
    .B(_0795_),
    .CO(_0798_),
    .S(_0799_));
 CLKBUF_X3 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 BUF_X1 _1470_ (.A(net21),
    .Z(scl_pad_o));
 BUF_X1 _1471_ (.A(net22),
    .Z(sda_pad_o));
 DFFR_X1 \al$_DFF_PN0_  (.D(_0000_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(al),
    .QN(_0755_));
 DFFR_X1 \byte_controller.ack_out$_DFFE_PN0P_  (.D(_0037_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.ack_out ),
    .QN(_0756_));
 DFFR_X1 \byte_controller.bit_controller.al$_DFF_PN0_  (.D(_0020_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.al ),
    .QN(_0757_));
 DFFR_X1 \byte_controller.bit_controller.busy$_DFF_PN0_  (.D(_0021_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.busy ),
    .QN(_0754_));
 DFFR_X1 \byte_controller.bit_controller.c_state[0]$_DFFE_PN0P_  (.D(_0038_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[0] ),
    .QN(_0753_));
 DFFR_X1 \byte_controller.bit_controller.c_state[10]$_DFFE_PN0P_  (.D(_0039_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[10] ),
    .QN(_0752_));
 DFFR_X1 \byte_controller.bit_controller.c_state[11]$_DFFE_PN0P_  (.D(_0040_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[11] ),
    .QN(_0751_));
 DFFR_X1 \byte_controller.bit_controller.c_state[12]$_DFFE_PN0P_  (.D(_0041_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[12] ),
    .QN(_0750_));
 DFFR_X1 \byte_controller.bit_controller.c_state[13]$_DFFE_PN0P_  (.D(_0042_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[13] ),
    .QN(_0749_));
 DFFR_X1 \byte_controller.bit_controller.c_state[14]$_DFFE_PN0P_  (.D(_0043_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[14] ),
    .QN(_0748_));
 DFFR_X1 \byte_controller.bit_controller.c_state[15]$_DFFE_PN0P_  (.D(_0044_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[15] ),
    .QN(_0747_));
 DFFR_X1 \byte_controller.bit_controller.c_state[16]$_DFFE_PN0P_  (.D(_0045_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[16] ),
    .QN(_0032_));
 DFFR_X1 \byte_controller.bit_controller.c_state[1]$_DFFE_PN0P_  (.D(_0046_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[1] ),
    .QN(_0746_));
 DFFR_X1 \byte_controller.bit_controller.c_state[2]$_DFFE_PN0P_  (.D(_0047_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[2] ),
    .QN(_0745_));
 DFFR_X1 \byte_controller.bit_controller.c_state[3]$_DFFE_PN0P_  (.D(_0048_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[3] ),
    .QN(_0744_));
 DFFR_X1 \byte_controller.bit_controller.c_state[4]$_DFFE_PN0P_  (.D(_0049_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[4] ),
    .QN(_0743_));
 DFFR_X1 \byte_controller.bit_controller.c_state[5]$_DFFE_PN0P_  (.D(_0050_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[5] ),
    .QN(_0742_));
 DFFR_X1 \byte_controller.bit_controller.c_state[6]$_DFFE_PN0P_  (.D(_0051_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[6] ),
    .QN(_0741_));
 DFFR_X1 \byte_controller.bit_controller.c_state[7]$_DFFE_PN0P_  (.D(_0052_),
    .RN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[7] ),
    .QN(_0740_));
 DFFR_X1 \byte_controller.bit_controller.c_state[8]$_DFFE_PN0P_  (.D(_0053_),
    .RN(net1),
    .CK(clknet_4_15_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[8] ),
    .QN(_0739_));
 DFFR_X1 \byte_controller.bit_controller.c_state[9]$_DFFE_PN0P_  (.D(_0054_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.c_state[9] ),
    .QN(_0758_));
 DFFS_X2 \byte_controller.bit_controller.clk_en$_DFF_PN1_  (.D(_0022_),
    .SN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_en ),
    .QN(_0031_));
 DFFR_X1 \byte_controller.bit_controller.cmd_ack$_DFF_PN0_  (.D(_0023_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cmd_ack ),
    .QN(_0033_));
 DFFR_X1 \byte_controller.bit_controller.cmd_stop$_DFFE_PN0P_  (.D(_0055_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cmd_stop ),
    .QN(_0738_));
 DFFR_X1 \byte_controller.bit_controller.cnt[0]$_DFFE_PN0P_  (.D(_0056_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[0] ),
    .QN(_0790_));
 DFFR_X1 \byte_controller.bit_controller.cnt[10]$_DFFE_PN0P_  (.D(_0057_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[10] ),
    .QN(_0737_));
 DFFR_X1 \byte_controller.bit_controller.cnt[11]$_DFFE_PN0P_  (.D(_0058_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[11] ),
    .QN(_0736_));
 DFFR_X2 \byte_controller.bit_controller.cnt[12]$_DFFE_PN0P_  (.D(_0059_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[12] ),
    .QN(_0735_));
 DFFR_X1 \byte_controller.bit_controller.cnt[13]$_DFFE_PN0P_  (.D(_0060_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[13] ),
    .QN(_0734_));
 DFFR_X1 \byte_controller.bit_controller.cnt[14]$_DFFE_PN0P_  (.D(_0061_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[14] ),
    .QN(_0733_));
 DFFR_X1 \byte_controller.bit_controller.cnt[15]$_DFFE_PN0P_  (.D(_0062_),
    .RN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[15] ),
    .QN(_0732_));
 DFFR_X1 \byte_controller.bit_controller.cnt[1]$_DFFE_PN0P_  (.D(_0063_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[1] ),
    .QN(_0791_));
 DFFR_X1 \byte_controller.bit_controller.cnt[2]$_DFFE_PN0P_  (.D(_0064_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[2] ),
    .QN(_0731_));
 DFFR_X1 \byte_controller.bit_controller.cnt[3]$_DFFE_PN0P_  (.D(_0065_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[3] ),
    .QN(_0730_));
 DFFR_X1 \byte_controller.bit_controller.cnt[4]$_DFFE_PN0P_  (.D(_0066_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[4] ),
    .QN(_0729_));
 DFFR_X1 \byte_controller.bit_controller.cnt[5]$_DFFE_PN0P_  (.D(_0067_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[5] ),
    .QN(_0728_));
 DFFR_X1 \byte_controller.bit_controller.cnt[6]$_DFFE_PN0P_  (.D(_0068_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[6] ),
    .QN(_0727_));
 DFFR_X1 \byte_controller.bit_controller.cnt[7]$_DFFE_PN0P_  (.D(_0069_),
    .RN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[7] ),
    .QN(_0726_));
 DFFR_X1 \byte_controller.bit_controller.cnt[8]$_DFFE_PN0P_  (.D(_0070_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[8] ),
    .QN(_0725_));
 DFFR_X1 \byte_controller.bit_controller.cnt[9]$_DFFE_PN0P_  (.D(_0071_),
    .RN(net1),
    .CK(clknet_4_7_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.cnt[9] ),
    .QN(_0759_));
 DFFS_X1 \byte_controller.bit_controller.dSCL$_DFF_PN1_  (.D(_0024_),
    .SN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.dSCL ),
    .QN(_0760_));
 DFFS_X1 \byte_controller.bit_controller.dSDA$_DFF_PN1_  (.D(_0025_),
    .SN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.dSDA ),
    .QN(_0724_));
 DFF_X1 \byte_controller.bit_controller.dout$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.dout ),
    .QN(_0761_));
 DFF_X1 \byte_controller.bit_controller.dscl_oen$_DFF_P_  (.D(net9),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.dscl_oen ),
    .QN(_0762_));
 DFFS_X1 \byte_controller.bit_controller.sSCL$_DFF_PN1_  (.D(_0026_),
    .SN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.sSCL ),
    .QN(_0034_));
 DFFS_X1 \byte_controller.bit_controller.sSDA$_DFF_PN1_  (.D(_0027_),
    .SN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.sSDA ),
    .QN(_0723_));
 DFFS_X1 \byte_controller.bit_controller.scl_oen$_DFFE_PN1P_  (.D(_0073_),
    .SN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(net9),
    .QN(_0722_));
 DFFR_X1 \byte_controller.bit_controller.sda_chk$_DFFE_PN0P_  (.D(_0074_),
    .RN(net1),
    .CK(clknet_4_13_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.sda_chk ),
    .QN(_0721_));
 DFFS_X1 \byte_controller.bit_controller.sda_oen$_DFFE_PN1P_  (.D(_0075_),
    .SN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(net10),
    .QN(_0763_));
 DFFR_X1 \byte_controller.bit_controller.sta_condition$_DFF_PN0_  (.D(_0028_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.sta_condition ),
    .QN(_0764_));
 DFFR_X1 \byte_controller.bit_controller.sto_condition$_DFF_PN0_  (.D(_0029_),
    .RN(net1),
    .CK(clknet_4_12_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.sto_condition ),
    .QN(_0765_));
 DFFS_X1 \byte_controller.c_state[0]$_DFF_PN1_  (.D(_0006_),
    .SN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.c_state[0] ),
    .QN(_0766_));
 DFFR_X1 \byte_controller.c_state[1]$_DFF_PN0_  (.D(_0007_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.c_state[1] ),
    .QN(_0767_));
 DFFR_X1 \byte_controller.c_state[2]$_DFF_PN0_  (.D(_0008_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.c_state[2] ),
    .QN(_0030_));
 DFFR_X1 \byte_controller.c_state[3]$_DFF_PN0_  (.D(_0009_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.c_state[3] ),
    .QN(_0768_));
 DFFR_X1 \byte_controller.c_state[4]$_DFF_PN0_  (.D(_0010_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.c_state[4] ),
    .QN(_0769_));
 DFFR_X1 \byte_controller.c_state[5]$_DFF_PN0_  (.D(_0011_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.c_state[5] ),
    .QN(_0770_));
 DFFR_X1 \byte_controller.cmd_ack$_DFF_PN0_  (.D(_0016_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.cmd_ack ),
    .QN(_0771_));
 DFFR_X1 \byte_controller.core_cmd[1]$_DFF_PN0_  (.D(_0012_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.core_cmd[1] ),
    .QN(_0772_));
 DFFR_X1 \byte_controller.core_cmd[2]$_DFF_PN0_  (.D(_0013_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.core_cmd[2] ),
    .QN(_0773_));
 DFFR_X1 \byte_controller.core_cmd[3]$_DFF_PN0_  (.D(_0014_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.core_cmd[3] ),
    .QN(_0774_));
 DFFR_X1 \byte_controller.core_cmd[4]$_DFF_PN0_  (.D(_0015_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(\byte_controller.core_cmd[4] ),
    .QN(_0775_));
 DFFR_X1 \byte_controller.core_txd$_DFF_PN0_  (.D(_0017_),
    .RN(net1),
    .CK(clknet_4_14_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.din ),
    .QN(_0720_));
 DFFR_X1 \byte_controller.dcnt[0]$_DFFE_PN0P_  (.D(_0076_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.dcnt[0] ),
    .QN(_0794_));
 DFFR_X1 \byte_controller.dcnt[1]$_DFFE_PN0P_  (.D(_0077_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.dcnt[1] ),
    .QN(_0795_));
 DFFR_X1 \byte_controller.dcnt[2]$_DFFE_PN0P_  (.D(_0078_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.dcnt[2] ),
    .QN(_0776_));
 DFFR_X1 \byte_controller.ld$_DFF_PN0_  (.D(_0018_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.ld ),
    .QN(_0036_));
 DFFR_X1 \byte_controller.shift$_DFF_PN0_  (.D(_0019_),
    .RN(net1),
    .CK(clknet_4_10_0_wb_clk_i),
    .Q(\byte_controller.shift ),
    .QN(_0719_));
 DFFR_X1 \byte_controller.sr[0]$_DFFE_PN0P_  (.D(_0079_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.dout[0] ),
    .QN(_0718_));
 DFFR_X1 \byte_controller.sr[1]$_DFFE_PN0P_  (.D(_0080_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\byte_controller.dout[1] ),
    .QN(_0717_));
 DFFR_X1 \byte_controller.sr[2]$_DFFE_PN0P_  (.D(_0081_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\byte_controller.dout[2] ),
    .QN(_0716_));
 DFFR_X1 \byte_controller.sr[3]$_DFFE_PN0P_  (.D(_0082_),
    .RN(net1),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(\byte_controller.dout[3] ),
    .QN(_0715_));
 DFFR_X1 \byte_controller.sr[4]$_DFFE_PN0P_  (.D(_0083_),
    .RN(net1),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(\byte_controller.dout[4] ),
    .QN(_0714_));
 DFFR_X1 \byte_controller.sr[5]$_DFFE_PN0P_  (.D(_0084_),
    .RN(net1),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(\byte_controller.dout[5] ),
    .QN(_0713_));
 DFFR_X1 \byte_controller.sr[6]$_DFFE_PN0P_  (.D(_0085_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.dout[6] ),
    .QN(_0712_));
 DFFR_X1 \byte_controller.sr[7]$_DFFE_PN0P_  (.D(_0086_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(\byte_controller.dout[7] ),
    .QN(_0711_));
 DFFR_X1 \cr[0]$_DFFE_PN0P_  (.D(_0087_),
    .RN(net1),
    .CK(clknet_4_3_0_wb_clk_i),
    .Q(\cr[0] ),
    .QN(_0710_));
 DFFR_X1 \cr[1]$_DFFE_PN0P_  (.D(_0088_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\cr[1] ),
    .QN(_0709_));
 DFFR_X1 \cr[2]$_DFFE_PN0P_  (.D(_0089_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\cr[2] ),
    .QN(_0708_));
 DFFR_X1 \cr[3]$_DFFE_PN0P_  (.D(_0090_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(ack),
    .QN(_0707_));
 DFFR_X2 \cr[4]$_DFFE_PN0P_  (.D(_0091_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(\byte_controller.write ),
    .QN(_0706_));
 DFFR_X1 \cr[5]$_DFFE_PN0P_  (.D(_0092_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(\byte_controller.read ),
    .QN(_0705_));
 DFFR_X1 \cr[6]$_DFFE_PN0P_  (.D(_0093_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(\byte_controller.stop ),
    .QN(_0704_));
 DFFR_X1 \cr[7]$_DFFE_PN0P_  (.D(_0094_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(\byte_controller.start ),
    .QN(_0703_));
 DFFR_X1 \ctr[0]$_DFFE_PN0P_  (.D(_0095_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\ctr[0] ),
    .QN(_0702_));
 DFFR_X1 \ctr[1]$_DFFE_PN0P_  (.D(_0096_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\ctr[1] ),
    .QN(_0701_));
 DFFR_X1 \ctr[2]$_DFFE_PN0P_  (.D(_0097_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\ctr[2] ),
    .QN(_0700_));
 DFFR_X1 \ctr[3]$_DFFE_PN0P_  (.D(_0098_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\ctr[3] ),
    .QN(_0699_));
 DFFR_X1 \ctr[4]$_DFFE_PN0P_  (.D(_0099_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\ctr[4] ),
    .QN(_0698_));
 DFFR_X1 \ctr[5]$_DFFE_PN0P_  (.D(_0100_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\ctr[5] ),
    .QN(_0697_));
 DFFR_X1 \ctr[6]$_DFFE_PN0P_  (.D(_0101_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\ctr[6] ),
    .QN(_0696_));
 DFFR_X1 \ctr[7]$_DFFE_PN0P_  (.D(_0102_),
    .RN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.ena ),
    .QN(_0777_));
 DFFR_X1 \irq_flag$_DFF_PN0_  (.D(_0001_),
    .RN(net1),
    .CK(clknet_4_9_0_wb_clk_i),
    .Q(irq_flag),
    .QN(_0695_));
 DFFS_X1 \prer[0]$_DFFE_PN1P_  (.D(_0103_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[0] ),
    .QN(_0035_));
 DFFS_X1 \prer[10]$_DFFE_PN1P_  (.D(_0104_),
    .SN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[10] ),
    .QN(_0694_));
 DFFS_X1 \prer[11]$_DFFE_PN1P_  (.D(_0105_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[11] ),
    .QN(_0693_));
 DFFS_X1 \prer[12]$_DFFE_PN1P_  (.D(_0106_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[12] ),
    .QN(_0692_));
 DFFS_X1 \prer[13]$_DFFE_PN1P_  (.D(_0107_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[13] ),
    .QN(_0691_));
 DFFS_X1 \prer[14]$_DFFE_PN1P_  (.D(_0108_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[14] ),
    .QN(_0690_));
 DFFS_X1 \prer[15]$_DFFE_PN1P_  (.D(_0109_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[15] ),
    .QN(_0689_));
 DFFS_X1 \prer[1]$_DFFE_PN1P_  (.D(_0110_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[1] ),
    .QN(_0688_));
 DFFS_X1 \prer[2]$_DFFE_PN1P_  (.D(_0111_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[2] ),
    .QN(_0687_));
 DFFS_X1 \prer[3]$_DFFE_PN1P_  (.D(_0112_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[3] ),
    .QN(_0686_));
 DFFS_X1 \prer[4]$_DFFE_PN1P_  (.D(_0113_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[4] ),
    .QN(_0685_));
 DFFS_X2 \prer[5]$_DFFE_PN1P_  (.D(_0114_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[5] ),
    .QN(_0684_));
 DFFS_X1 \prer[6]$_DFFE_PN1P_  (.D(_0115_),
    .SN(net1),
    .CK(clknet_4_5_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[6] ),
    .QN(_0683_));
 DFFS_X1 \prer[7]$_DFFE_PN1P_  (.D(_0116_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[7] ),
    .QN(_0682_));
 DFFS_X1 \prer[8]$_DFFE_PN1P_  (.D(_0117_),
    .SN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[8] ),
    .QN(_0681_));
 DFFS_X1 \prer[9]$_DFFE_PN1P_  (.D(_0118_),
    .SN(net1),
    .CK(clknet_4_4_0_wb_clk_i),
    .Q(\byte_controller.bit_controller.clk_cnt[9] ),
    .QN(_0778_));
 DFFR_X1 \rxack$_DFF_PN0_  (.D(_0002_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(rxack),
    .QN(_0779_));
 DFFR_X1 \tip$_DFF_PN0_  (.D(_0003_),
    .RN(net1),
    .CK(clknet_4_11_0_wb_clk_i),
    .Q(tip),
    .QN(_0680_));
 DFFR_X1 \txr[0]$_DFFE_PN0P_  (.D(_0119_),
    .RN(net1),
    .CK(clknet_4_3_0_wb_clk_i),
    .Q(\byte_controller.din[0] ),
    .QN(_0679_));
 DFFR_X1 \txr[1]$_DFFE_PN0P_  (.D(_0120_),
    .RN(net1),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(\byte_controller.din[1] ),
    .QN(_0678_));
 DFFR_X1 \txr[2]$_DFFE_PN0P_  (.D(_0121_),
    .RN(net1),
    .CK(clknet_4_3_0_wb_clk_i),
    .Q(\byte_controller.din[2] ),
    .QN(_0677_));
 DFFR_X1 \txr[3]$_DFFE_PN0P_  (.D(_0122_),
    .RN(net1),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(\byte_controller.din[3] ),
    .QN(_0676_));
 DFFR_X1 \txr[4]$_DFFE_PN0P_  (.D(_0123_),
    .RN(net1),
    .CK(clknet_4_3_0_wb_clk_i),
    .Q(\byte_controller.din[4] ),
    .QN(_0675_));
 DFFR_X1 \txr[5]$_DFFE_PN0P_  (.D(_0124_),
    .RN(net1),
    .CK(clknet_4_3_0_wb_clk_i),
    .Q(\byte_controller.din[5] ),
    .QN(_0674_));
 DFFR_X1 \txr[6]$_DFFE_PN0P_  (.D(_0125_),
    .RN(net1),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(\byte_controller.din[6] ),
    .QN(_0673_));
 DFFR_X1 \txr[7]$_DFFE_PN0P_  (.D(_0126_),
    .RN(net1),
    .CK(clknet_4_6_0_wb_clk_i),
    .Q(\byte_controller.din[7] ),
    .QN(_0780_));
 DFF_X1 \wb_ack_o$_DFF_P_  (.D(_0004_),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(net11),
    .QN(_0781_));
 DFF_X1 \wb_dat_o[0]$_DFF_P_  (.D(_0664_),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(net12),
    .QN(_0782_));
 DFF_X1 \wb_dat_o[1]$_DFF_P_  (.D(_0665_),
    .CK(clknet_4_1_0_wb_clk_i),
    .Q(net13),
    .QN(_0783_));
 DFF_X1 \wb_dat_o[2]$_DFF_P_  (.D(_0666_),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(net14),
    .QN(_0784_));
 DFF_X1 \wb_dat_o[3]$_DFF_P_  (.D(_0667_),
    .CK(clknet_4_0_0_wb_clk_i),
    .Q(net15),
    .QN(_0785_));
 DFF_X1 \wb_dat_o[4]$_DFF_P_  (.D(_0668_),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(net16),
    .QN(_0786_));
 DFF_X1 \wb_dat_o[5]$_DFF_P_  (.D(_0669_),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(net17),
    .QN(_0787_));
 DFF_X1 \wb_dat_o[6]$_DFF_P_  (.D(_0670_),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(net18),
    .QN(_0788_));
 DFF_X1 \wb_dat_o[7]$_DFF_P_  (.D(_0671_),
    .CK(clknet_4_2_0_wb_clk_i),
    .Q(net19),
    .QN(_0789_));
 DFFR_X1 \wb_inta_o$_DFF_PN0_  (.D(_0005_),
    .RN(net1),
    .CK(clknet_4_8_0_wb_clk_i),
    .Q(net20),
    .QN(_0672_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_69 ();
 BUF_X32 input1 (.A(net23),
    .Z(net1));
 BUF_X1 input2 (.A(scl_pad_i),
    .Z(net2));
 BUF_X1 input3 (.A(sda_pad_i),
    .Z(net3));
 BUF_X1 input4 (.A(wb_adr_i[2]),
    .Z(net4));
 BUF_X1 input5 (.A(wb_cyc_i),
    .Z(net5));
 BUF_X1 input6 (.A(wb_rst_i),
    .Z(net6));
 BUF_X1 input7 (.A(wb_stb_i),
    .Z(net7));
 BUF_X1 input8 (.A(wb_we_i),
    .Z(net8));
 BUF_X1 output9 (.A(net9),
    .Z(scl_padoen_o));
 BUF_X1 output10 (.A(net10),
    .Z(sda_padoen_o));
 BUF_X1 output11 (.A(net11),
    .Z(wb_ack_o));
 BUF_X1 output12 (.A(net12),
    .Z(wb_dat_o[0]));
 BUF_X1 output13 (.A(net13),
    .Z(wb_dat_o[1]));
 BUF_X1 output14 (.A(net14),
    .Z(wb_dat_o[2]));
 BUF_X1 output15 (.A(net15),
    .Z(wb_dat_o[3]));
 BUF_X1 output16 (.A(net16),
    .Z(wb_dat_o[4]));
 BUF_X1 output17 (.A(net17),
    .Z(wb_dat_o[5]));
 BUF_X1 output18 (.A(net18),
    .Z(wb_dat_o[6]));
 BUF_X1 output19 (.A(net19),
    .Z(wb_dat_o[7]));
 BUF_X1 output20 (.A(net20),
    .Z(wb_inta_o));
 LOGIC0_X1 _1470__21 (.Z(net21));
 LOGIC0_X1 _1471__22 (.Z(net22));
 CLKBUF_X3 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_0_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_1_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_2_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_3_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_4_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_5_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_6_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_7_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_8_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_9_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_10_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_11_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_12_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_13_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_14_0_wb_clk_i));
 CLKBUF_X3 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .Z(clknet_4_15_0_wb_clk_i));
 INV_X1 clkload0 (.A(clknet_4_0_0_wb_clk_i));
 INV_X2 clkload1 (.A(clknet_4_1_0_wb_clk_i));
 INV_X2 clkload2 (.A(clknet_4_2_0_wb_clk_i));
 INV_X4 clkload3 (.A(clknet_4_3_0_wb_clk_i));
 INV_X1 clkload4 (.A(clknet_4_4_0_wb_clk_i));
 INV_X2 clkload5 (.A(clknet_4_6_0_wb_clk_i));
 INV_X4 clkload6 (.A(clknet_4_7_0_wb_clk_i));
 CLKBUF_X1 clkload7 (.A(clknet_4_8_0_wb_clk_i));
 INV_X4 clkload8 (.A(clknet_4_9_0_wb_clk_i));
 INV_X2 clkload9 (.A(clknet_4_10_0_wb_clk_i));
 CLKBUF_X1 clkload10 (.A(clknet_4_11_0_wb_clk_i));
 INV_X2 clkload11 (.A(clknet_4_12_0_wb_clk_i));
 CLKBUF_X1 clkload12 (.A(clknet_4_13_0_wb_clk_i));
 INV_X2 clkload13 (.A(clknet_4_14_0_wb_clk_i));
 INV_X1 clkload14 (.A(clknet_4_15_0_wb_clk_i));
 CLKBUF_X1 hold1 (.A(arst_i),
    .Z(net23));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X8 FILLER_0_33 ();
 FILLCELL_X4 FILLER_0_41 ();
 FILLCELL_X8 FILLER_0_68 ();
 FILLCELL_X4 FILLER_0_96 ();
 FILLCELL_X1 FILLER_0_100 ();
 FILLCELL_X4 FILLER_0_141 ();
 FILLCELL_X2 FILLER_0_157 ();
 FILLCELL_X2 FILLER_0_168 ();
 FILLCELL_X32 FILLER_0_187 ();
 FILLCELL_X32 FILLER_0_219 ();
 FILLCELL_X8 FILLER_0_251 ();
 FILLCELL_X4 FILLER_0_259 ();
 FILLCELL_X1 FILLER_0_263 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_41 ();
 FILLCELL_X2 FILLER_1_45 ();
 FILLCELL_X1 FILLER_1_47 ();
 FILLCELL_X16 FILLER_1_85 ();
 FILLCELL_X4 FILLER_1_101 ();
 FILLCELL_X2 FILLER_1_105 ();
 FILLCELL_X8 FILLER_1_127 ();
 FILLCELL_X1 FILLER_1_135 ();
 FILLCELL_X8 FILLER_1_139 ();
 FILLCELL_X32 FILLER_1_160 ();
 FILLCELL_X32 FILLER_1_192 ();
 FILLCELL_X16 FILLER_1_224 ();
 FILLCELL_X4 FILLER_1_240 ();
 FILLCELL_X2 FILLER_1_244 ();
 FILLCELL_X1 FILLER_1_246 ();
 FILLCELL_X4 FILLER_1_250 ();
 FILLCELL_X2 FILLER_1_254 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_53 ();
 FILLCELL_X4 FILLER_2_74 ();
 FILLCELL_X2 FILLER_2_118 ();
 FILLCELL_X8 FILLER_2_157 ();
 FILLCELL_X2 FILLER_2_165 ();
 FILLCELL_X2 FILLER_2_192 ();
 FILLCELL_X1 FILLER_2_194 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X4 FILLER_3_25 ();
 FILLCELL_X2 FILLER_3_29 ();
 FILLCELL_X8 FILLER_3_51 ();
 FILLCELL_X2 FILLER_3_86 ();
 FILLCELL_X8 FILLER_3_91 ();
 FILLCELL_X2 FILLER_3_99 ();
 FILLCELL_X2 FILLER_3_111 ();
 FILLCELL_X1 FILLER_3_113 ();
 FILLCELL_X8 FILLER_3_124 ();
 FILLCELL_X4 FILLER_3_162 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X4 FILLER_3_170 ();
 FILLCELL_X1 FILLER_3_174 ();
 FILLCELL_X2 FILLER_3_179 ();
 FILLCELL_X1 FILLER_3_185 ();
 FILLCELL_X1 FILLER_3_198 ();
 FILLCELL_X2 FILLER_3_205 ();
 FILLCELL_X32 FILLER_3_211 ();
 FILLCELL_X8 FILLER_3_243 ();
 FILLCELL_X1 FILLER_3_251 ();
 FILLCELL_X8 FILLER_3_254 ();
 FILLCELL_X2 FILLER_3_262 ();
 FILLCELL_X8 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_9 ();
 FILLCELL_X1 FILLER_4_13 ();
 FILLCELL_X8 FILLER_4_34 ();
 FILLCELL_X2 FILLER_4_62 ();
 FILLCELL_X1 FILLER_4_86 ();
 FILLCELL_X4 FILLER_4_94 ();
 FILLCELL_X2 FILLER_4_98 ();
 FILLCELL_X2 FILLER_4_104 ();
 FILLCELL_X2 FILLER_4_109 ();
 FILLCELL_X1 FILLER_4_111 ();
 FILLCELL_X8 FILLER_4_152 ();
 FILLCELL_X4 FILLER_4_160 ();
 FILLCELL_X1 FILLER_4_164 ();
 FILLCELL_X8 FILLER_4_201 ();
 FILLCELL_X1 FILLER_4_229 ();
 FILLCELL_X16 FILLER_4_235 ();
 FILLCELL_X8 FILLER_4_251 ();
 FILLCELL_X4 FILLER_4_259 ();
 FILLCELL_X1 FILLER_4_263 ();
 FILLCELL_X2 FILLER_5_1 ();
 FILLCELL_X1 FILLER_5_3 ();
 FILLCELL_X1 FILLER_5_31 ();
 FILLCELL_X4 FILLER_5_39 ();
 FILLCELL_X2 FILLER_5_43 ();
 FILLCELL_X4 FILLER_5_59 ();
 FILLCELL_X2 FILLER_5_63 ();
 FILLCELL_X1 FILLER_5_65 ();
 FILLCELL_X4 FILLER_5_72 ();
 FILLCELL_X8 FILLER_5_79 ();
 FILLCELL_X1 FILLER_5_109 ();
 FILLCELL_X2 FILLER_5_131 ();
 FILLCELL_X1 FILLER_5_133 ();
 FILLCELL_X8 FILLER_5_171 ();
 FILLCELL_X4 FILLER_5_179 ();
 FILLCELL_X4 FILLER_5_188 ();
 FILLCELL_X2 FILLER_5_192 ();
 FILLCELL_X2 FILLER_5_209 ();
 FILLCELL_X32 FILLER_5_231 ();
 FILLCELL_X1 FILLER_5_263 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_20 ();
 FILLCELL_X1 FILLER_6_24 ();
 FILLCELL_X4 FILLER_6_28 ();
 FILLCELL_X8 FILLER_6_35 ();
 FILLCELL_X1 FILLER_6_57 ();
 FILLCELL_X8 FILLER_6_65 ();
 FILLCELL_X2 FILLER_6_73 ();
 FILLCELL_X4 FILLER_6_122 ();
 FILLCELL_X1 FILLER_6_126 ();
 FILLCELL_X1 FILLER_6_130 ();
 FILLCELL_X8 FILLER_6_142 ();
 FILLCELL_X16 FILLER_6_155 ();
 FILLCELL_X1 FILLER_6_194 ();
 FILLCELL_X2 FILLER_6_202 ();
 FILLCELL_X32 FILLER_6_228 ();
 FILLCELL_X4 FILLER_6_260 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_5 ();
 FILLCELL_X2 FILLER_7_30 ();
 FILLCELL_X1 FILLER_7_62 ();
 FILLCELL_X1 FILLER_7_68 ();
 FILLCELL_X1 FILLER_7_89 ();
 FILLCELL_X2 FILLER_7_93 ();
 FILLCELL_X1 FILLER_7_114 ();
 FILLCELL_X8 FILLER_7_125 ();
 FILLCELL_X4 FILLER_7_138 ();
 FILLCELL_X4 FILLER_7_169 ();
 FILLCELL_X2 FILLER_7_173 ();
 FILLCELL_X1 FILLER_7_175 ();
 FILLCELL_X2 FILLER_7_187 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X4 FILLER_7_257 ();
 FILLCELL_X2 FILLER_7_261 ();
 FILLCELL_X1 FILLER_7_263 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_9 ();
 FILLCELL_X16 FILLER_8_20 ();
 FILLCELL_X2 FILLER_8_36 ();
 FILLCELL_X2 FILLER_8_41 ();
 FILLCELL_X1 FILLER_8_43 ();
 FILLCELL_X1 FILLER_8_85 ();
 FILLCELL_X8 FILLER_8_103 ();
 FILLCELL_X2 FILLER_8_111 ();
 FILLCELL_X2 FILLER_8_123 ();
 FILLCELL_X1 FILLER_8_125 ();
 FILLCELL_X2 FILLER_8_142 ();
 FILLCELL_X8 FILLER_8_166 ();
 FILLCELL_X2 FILLER_8_174 ();
 FILLCELL_X1 FILLER_8_176 ();
 FILLCELL_X1 FILLER_8_197 ();
 FILLCELL_X1 FILLER_8_201 ();
 FILLCELL_X1 FILLER_8_208 ();
 FILLCELL_X16 FILLER_8_243 ();
 FILLCELL_X4 FILLER_8_259 ();
 FILLCELL_X1 FILLER_8_263 ();
 FILLCELL_X4 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_5 ();
 FILLCELL_X1 FILLER_9_7 ();
 FILLCELL_X2 FILLER_9_33 ();
 FILLCELL_X1 FILLER_9_66 ();
 FILLCELL_X2 FILLER_9_74 ();
 FILLCELL_X1 FILLER_9_80 ();
 FILLCELL_X2 FILLER_9_87 ();
 FILLCELL_X2 FILLER_9_112 ();
 FILLCELL_X1 FILLER_9_114 ();
 FILLCELL_X1 FILLER_9_118 ();
 FILLCELL_X4 FILLER_9_156 ();
 FILLCELL_X1 FILLER_9_160 ();
 FILLCELL_X4 FILLER_9_165 ();
 FILLCELL_X2 FILLER_9_192 ();
 FILLCELL_X1 FILLER_9_240 ();
 FILLCELL_X16 FILLER_9_243 ();
 FILLCELL_X4 FILLER_9_259 ();
 FILLCELL_X1 FILLER_9_263 ();
 FILLCELL_X4 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_5 ();
 FILLCELL_X2 FILLER_10_26 ();
 FILLCELL_X1 FILLER_10_35 ();
 FILLCELL_X2 FILLER_10_44 ();
 FILLCELL_X1 FILLER_10_55 ();
 FILLCELL_X1 FILLER_10_98 ();
 FILLCELL_X2 FILLER_10_188 ();
 FILLCELL_X2 FILLER_10_197 ();
 FILLCELL_X1 FILLER_10_203 ();
 FILLCELL_X2 FILLER_10_207 ();
 FILLCELL_X32 FILLER_10_222 ();
 FILLCELL_X8 FILLER_10_254 ();
 FILLCELL_X2 FILLER_10_262 ();
 FILLCELL_X1 FILLER_11_1 ();
 FILLCELL_X8 FILLER_11_5 ();
 FILLCELL_X2 FILLER_11_13 ();
 FILLCELL_X4 FILLER_11_19 ();
 FILLCELL_X2 FILLER_11_23 ();
 FILLCELL_X1 FILLER_11_25 ();
 FILLCELL_X2 FILLER_11_29 ();
 FILLCELL_X2 FILLER_11_63 ();
 FILLCELL_X1 FILLER_11_65 ();
 FILLCELL_X1 FILLER_11_72 ();
 FILLCELL_X1 FILLER_11_101 ();
 FILLCELL_X1 FILLER_11_105 ();
 FILLCELL_X2 FILLER_11_116 ();
 FILLCELL_X1 FILLER_11_118 ();
 FILLCELL_X8 FILLER_11_153 ();
 FILLCELL_X2 FILLER_11_161 ();
 FILLCELL_X1 FILLER_11_163 ();
 FILLCELL_X8 FILLER_11_167 ();
 FILLCELL_X2 FILLER_11_175 ();
 FILLCELL_X1 FILLER_11_216 ();
 FILLCELL_X16 FILLER_11_237 ();
 FILLCELL_X8 FILLER_11_253 ();
 FILLCELL_X2 FILLER_11_261 ();
 FILLCELL_X1 FILLER_11_263 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_24 ();
 FILLCELL_X1 FILLER_12_38 ();
 FILLCELL_X2 FILLER_12_66 ();
 FILLCELL_X1 FILLER_12_132 ();
 FILLCELL_X8 FILLER_12_135 ();
 FILLCELL_X1 FILLER_12_143 ();
 FILLCELL_X1 FILLER_12_148 ();
 FILLCELL_X1 FILLER_12_169 ();
 FILLCELL_X1 FILLER_12_190 ();
 FILLCELL_X1 FILLER_12_216 ();
 FILLCELL_X2 FILLER_12_222 ();
 FILLCELL_X16 FILLER_12_246 ();
 FILLCELL_X2 FILLER_12_262 ();
 FILLCELL_X2 FILLER_13_31 ();
 FILLCELL_X1 FILLER_13_33 ();
 FILLCELL_X2 FILLER_13_112 ();
 FILLCELL_X1 FILLER_13_121 ();
 FILLCELL_X4 FILLER_13_146 ();
 FILLCELL_X1 FILLER_13_170 ();
 FILLCELL_X4 FILLER_13_178 ();
 FILLCELL_X4 FILLER_13_185 ();
 FILLCELL_X2 FILLER_13_189 ();
 FILLCELL_X4 FILLER_13_196 ();
 FILLCELL_X1 FILLER_13_200 ();
 FILLCELL_X2 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_219 ();
 FILLCELL_X16 FILLER_13_224 ();
 FILLCELL_X2 FILLER_13_240 ();
 FILLCELL_X2 FILLER_13_262 ();
 FILLCELL_X2 FILLER_14_4 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_13 ();
 FILLCELL_X1 FILLER_14_15 ();
 FILLCELL_X1 FILLER_14_19 ();
 FILLCELL_X2 FILLER_14_23 ();
 FILLCELL_X2 FILLER_14_32 ();
 FILLCELL_X2 FILLER_14_39 ();
 FILLCELL_X1 FILLER_14_41 ();
 FILLCELL_X1 FILLER_14_59 ();
 FILLCELL_X1 FILLER_14_74 ();
 FILLCELL_X2 FILLER_14_82 ();
 FILLCELL_X2 FILLER_14_87 ();
 FILLCELL_X1 FILLER_14_98 ();
 FILLCELL_X4 FILLER_14_122 ();
 FILLCELL_X2 FILLER_14_126 ();
 FILLCELL_X1 FILLER_14_128 ();
 FILLCELL_X8 FILLER_14_136 ();
 FILLCELL_X4 FILLER_14_144 ();
 FILLCELL_X2 FILLER_14_148 ();
 FILLCELL_X2 FILLER_14_178 ();
 FILLCELL_X1 FILLER_14_180 ();
 FILLCELL_X1 FILLER_14_210 ();
 FILLCELL_X8 FILLER_14_255 ();
 FILLCELL_X1 FILLER_14_263 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_85 ();
 FILLCELL_X1 FILLER_15_98 ();
 FILLCELL_X1 FILLER_15_106 ();
 FILLCELL_X8 FILLER_15_151 ();
 FILLCELL_X4 FILLER_15_159 ();
 FILLCELL_X2 FILLER_15_163 ();
 FILLCELL_X2 FILLER_15_205 ();
 FILLCELL_X2 FILLER_15_211 ();
 FILLCELL_X1 FILLER_15_213 ();
 FILLCELL_X2 FILLER_15_217 ();
 FILLCELL_X1 FILLER_15_219 ();
 FILLCELL_X8 FILLER_15_223 ();
 FILLCELL_X1 FILLER_15_231 ();
 FILLCELL_X4 FILLER_15_236 ();
 FILLCELL_X1 FILLER_15_240 ();
 FILLCELL_X1 FILLER_15_247 ();
 FILLCELL_X1 FILLER_15_251 ();
 FILLCELL_X8 FILLER_15_256 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X1 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_18 ();
 FILLCELL_X1 FILLER_16_20 ();
 FILLCELL_X4 FILLER_16_32 ();
 FILLCELL_X2 FILLER_16_36 ();
 FILLCELL_X4 FILLER_16_49 ();
 FILLCELL_X2 FILLER_16_53 ();
 FILLCELL_X1 FILLER_16_55 ();
 FILLCELL_X2 FILLER_16_90 ();
 FILLCELL_X2 FILLER_16_99 ();
 FILLCELL_X4 FILLER_16_121 ();
 FILLCELL_X4 FILLER_16_130 ();
 FILLCELL_X1 FILLER_16_134 ();
 FILLCELL_X16 FILLER_16_147 ();
 FILLCELL_X8 FILLER_16_163 ();
 FILLCELL_X1 FILLER_16_171 ();
 FILLCELL_X1 FILLER_16_181 ();
 FILLCELL_X16 FILLER_16_184 ();
 FILLCELL_X1 FILLER_16_200 ();
 FILLCELL_X16 FILLER_16_221 ();
 FILLCELL_X4 FILLER_16_237 ();
 FILLCELL_X1 FILLER_16_241 ();
 FILLCELL_X2 FILLER_16_262 ();
 FILLCELL_X1 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_5 ();
 FILLCELL_X1 FILLER_17_26 ();
 FILLCELL_X1 FILLER_17_47 ();
 FILLCELL_X1 FILLER_17_53 ();
 FILLCELL_X1 FILLER_17_61 ();
 FILLCELL_X2 FILLER_17_66 ();
 FILLCELL_X2 FILLER_17_75 ();
 FILLCELL_X2 FILLER_17_97 ();
 FILLCELL_X1 FILLER_17_111 ();
 FILLCELL_X8 FILLER_17_117 ();
 FILLCELL_X4 FILLER_17_125 ();
 FILLCELL_X2 FILLER_17_129 ();
 FILLCELL_X1 FILLER_17_131 ();
 FILLCELL_X2 FILLER_17_152 ();
 FILLCELL_X16 FILLER_17_158 ();
 FILLCELL_X4 FILLER_17_174 ();
 FILLCELL_X2 FILLER_17_178 ();
 FILLCELL_X1 FILLER_17_180 ();
 FILLCELL_X8 FILLER_17_207 ();
 FILLCELL_X2 FILLER_17_215 ();
 FILLCELL_X1 FILLER_17_222 ();
 FILLCELL_X1 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_10 ();
 FILLCELL_X1 FILLER_18_16 ();
 FILLCELL_X1 FILLER_18_28 ();
 FILLCELL_X1 FILLER_18_36 ();
 FILLCELL_X1 FILLER_18_51 ();
 FILLCELL_X1 FILLER_18_54 ();
 FILLCELL_X1 FILLER_18_62 ();
 FILLCELL_X2 FILLER_18_84 ();
 FILLCELL_X2 FILLER_18_93 ();
 FILLCELL_X1 FILLER_18_102 ();
 FILLCELL_X4 FILLER_18_125 ();
 FILLCELL_X2 FILLER_18_129 ();
 FILLCELL_X1 FILLER_18_131 ();
 FILLCELL_X8 FILLER_18_137 ();
 FILLCELL_X4 FILLER_18_145 ();
 FILLCELL_X8 FILLER_18_176 ();
 FILLCELL_X4 FILLER_18_184 ();
 FILLCELL_X2 FILLER_18_206 ();
 FILLCELL_X1 FILLER_18_208 ();
 FILLCELL_X4 FILLER_18_212 ();
 FILLCELL_X2 FILLER_18_216 ();
 FILLCELL_X1 FILLER_18_218 ();
 FILLCELL_X4 FILLER_18_260 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X1 FILLER_19_50 ();
 FILLCELL_X2 FILLER_19_71 ();
 FILLCELL_X8 FILLER_19_95 ();
 FILLCELL_X1 FILLER_19_103 ();
 FILLCELL_X4 FILLER_19_124 ();
 FILLCELL_X1 FILLER_19_128 ();
 FILLCELL_X8 FILLER_19_149 ();
 FILLCELL_X4 FILLER_19_181 ();
 FILLCELL_X2 FILLER_19_185 ();
 FILLCELL_X1 FILLER_19_187 ();
 FILLCELL_X8 FILLER_19_191 ();
 FILLCELL_X4 FILLER_19_199 ();
 FILLCELL_X1 FILLER_19_203 ();
 FILLCELL_X2 FILLER_19_207 ();
 FILLCELL_X1 FILLER_19_228 ();
 FILLCELL_X1 FILLER_19_232 ();
 FILLCELL_X8 FILLER_19_253 ();
 FILLCELL_X2 FILLER_19_261 ();
 FILLCELL_X1 FILLER_19_263 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_9 ();
 FILLCELL_X1 FILLER_20_14 ();
 FILLCELL_X32 FILLER_20_61 ();
 FILLCELL_X4 FILLER_20_93 ();
 FILLCELL_X2 FILLER_20_97 ();
 FILLCELL_X1 FILLER_20_99 ();
 FILLCELL_X8 FILLER_20_108 ();
 FILLCELL_X1 FILLER_20_116 ();
 FILLCELL_X8 FILLER_20_121 ();
 FILLCELL_X1 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_155 ();
 FILLCELL_X2 FILLER_20_185 ();
 FILLCELL_X1 FILLER_20_194 ();
 FILLCELL_X2 FILLER_20_206 ();
 FILLCELL_X2 FILLER_20_235 ();
 FILLCELL_X2 FILLER_20_261 ();
 FILLCELL_X1 FILLER_20_263 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X16 FILLER_21_25 ();
 FILLCELL_X4 FILLER_21_51 ();
 FILLCELL_X2 FILLER_21_55 ();
 FILLCELL_X1 FILLER_21_77 ();
 FILLCELL_X2 FILLER_21_83 ();
 FILLCELL_X4 FILLER_21_94 ();
 FILLCELL_X2 FILLER_21_98 ();
 FILLCELL_X1 FILLER_21_100 ();
 FILLCELL_X16 FILLER_21_104 ();
 FILLCELL_X4 FILLER_21_120 ();
 FILLCELL_X1 FILLER_21_124 ();
 FILLCELL_X4 FILLER_21_155 ();
 FILLCELL_X1 FILLER_21_159 ();
 FILLCELL_X2 FILLER_21_167 ();
 FILLCELL_X2 FILLER_21_171 ();
 FILLCELL_X1 FILLER_21_180 ();
 FILLCELL_X1 FILLER_21_190 ();
 FILLCELL_X1 FILLER_21_199 ();
 FILLCELL_X1 FILLER_21_220 ();
 FILLCELL_X1 FILLER_21_229 ();
 FILLCELL_X1 FILLER_21_263 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_25 ();
 FILLCELL_X4 FILLER_22_30 ();
 FILLCELL_X2 FILLER_22_34 ();
 FILLCELL_X1 FILLER_22_36 ();
 FILLCELL_X4 FILLER_22_46 ();
 FILLCELL_X2 FILLER_22_50 ();
 FILLCELL_X1 FILLER_22_52 ();
 FILLCELL_X2 FILLER_22_66 ();
 FILLCELL_X1 FILLER_22_68 ();
 FILLCELL_X4 FILLER_22_72 ();
 FILLCELL_X4 FILLER_22_96 ();
 FILLCELL_X1 FILLER_22_100 ();
 FILLCELL_X2 FILLER_22_106 ();
 FILLCELL_X8 FILLER_22_114 ();
 FILLCELL_X4 FILLER_22_122 ();
 FILLCELL_X2 FILLER_22_150 ();
 FILLCELL_X1 FILLER_22_152 ();
 FILLCELL_X2 FILLER_22_173 ();
 FILLCELL_X1 FILLER_22_175 ();
 FILLCELL_X2 FILLER_22_184 ();
 FILLCELL_X2 FILLER_22_240 ();
 FILLCELL_X2 FILLER_22_262 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X2 FILLER_23_5 ();
 FILLCELL_X1 FILLER_23_27 ();
 FILLCELL_X1 FILLER_23_31 ();
 FILLCELL_X1 FILLER_23_39 ();
 FILLCELL_X4 FILLER_23_43 ();
 FILLCELL_X2 FILLER_23_47 ();
 FILLCELL_X1 FILLER_23_49 ();
 FILLCELL_X4 FILLER_23_126 ();
 FILLCELL_X2 FILLER_23_130 ();
 FILLCELL_X4 FILLER_23_137 ();
 FILLCELL_X16 FILLER_23_161 ();
 FILLCELL_X2 FILLER_23_177 ();
 FILLCELL_X1 FILLER_23_179 ();
 FILLCELL_X4 FILLER_23_259 ();
 FILLCELL_X1 FILLER_23_263 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X16 FILLER_24_49 ();
 FILLCELL_X4 FILLER_24_65 ();
 FILLCELL_X1 FILLER_24_108 ();
 FILLCELL_X2 FILLER_24_117 ();
 FILLCELL_X4 FILLER_24_139 ();
 FILLCELL_X2 FILLER_24_179 ();
 FILLCELL_X1 FILLER_24_181 ();
 FILLCELL_X1 FILLER_24_218 ();
 FILLCELL_X1 FILLER_24_237 ();
 FILLCELL_X1 FILLER_24_240 ();
 FILLCELL_X1 FILLER_24_245 ();
 FILLCELL_X2 FILLER_24_250 ();
 FILLCELL_X2 FILLER_24_261 ();
 FILLCELL_X1 FILLER_24_263 ();
 FILLCELL_X4 FILLER_25_1 ();
 FILLCELL_X1 FILLER_25_35 ();
 FILLCELL_X1 FILLER_25_44 ();
 FILLCELL_X4 FILLER_25_53 ();
 FILLCELL_X4 FILLER_25_61 ();
 FILLCELL_X1 FILLER_25_65 ();
 FILLCELL_X2 FILLER_25_111 ();
 FILLCELL_X1 FILLER_25_116 ();
 FILLCELL_X1 FILLER_25_123 ();
 FILLCELL_X8 FILLER_25_130 ();
 FILLCELL_X4 FILLER_25_138 ();
 FILLCELL_X2 FILLER_25_145 ();
 FILLCELL_X1 FILLER_25_147 ();
 FILLCELL_X8 FILLER_25_167 ();
 FILLCELL_X1 FILLER_25_186 ();
 FILLCELL_X1 FILLER_25_191 ();
 FILLCELL_X1 FILLER_25_210 ();
 FILLCELL_X1 FILLER_25_218 ();
 FILLCELL_X2 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_112 ();
 FILLCELL_X4 FILLER_26_119 ();
 FILLCELL_X2 FILLER_26_123 ();
 FILLCELL_X16 FILLER_26_145 ();
 FILLCELL_X8 FILLER_26_161 ();
 FILLCELL_X2 FILLER_26_169 ();
 FILLCELL_X4 FILLER_26_175 ();
 FILLCELL_X1 FILLER_26_179 ();
 FILLCELL_X1 FILLER_26_234 ();
 FILLCELL_X2 FILLER_26_262 ();
 FILLCELL_X16 FILLER_27_1 ();
 FILLCELL_X4 FILLER_27_17 ();
 FILLCELL_X2 FILLER_27_21 ();
 FILLCELL_X1 FILLER_27_64 ();
 FILLCELL_X2 FILLER_27_74 ();
 FILLCELL_X1 FILLER_27_80 ();
 FILLCELL_X1 FILLER_27_85 ();
 FILLCELL_X1 FILLER_27_99 ();
 FILLCELL_X16 FILLER_27_141 ();
 FILLCELL_X2 FILLER_27_157 ();
 FILLCELL_X4 FILLER_27_179 ();
 FILLCELL_X2 FILLER_27_183 ();
 FILLCELL_X1 FILLER_27_185 ();
 FILLCELL_X1 FILLER_27_192 ();
 FILLCELL_X1 FILLER_27_202 ();
 FILLCELL_X1 FILLER_27_211 ();
 FILLCELL_X2 FILLER_27_239 ();
 FILLCELL_X1 FILLER_27_241 ();
 FILLCELL_X1 FILLER_27_245 ();
 FILLCELL_X8 FILLER_27_252 ();
 FILLCELL_X4 FILLER_27_260 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X4 FILLER_28_17 ();
 FILLCELL_X1 FILLER_28_75 ();
 FILLCELL_X2 FILLER_28_80 ();
 FILLCELL_X1 FILLER_28_86 ();
 FILLCELL_X1 FILLER_28_115 ();
 FILLCELL_X2 FILLER_28_126 ();
 FILLCELL_X16 FILLER_28_148 ();
 FILLCELL_X8 FILLER_28_164 ();
 FILLCELL_X1 FILLER_28_223 ();
 FILLCELL_X1 FILLER_28_240 ();
 FILLCELL_X16 FILLER_28_246 ();
 FILLCELL_X2 FILLER_28_262 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X8 FILLER_29_33 ();
 FILLCELL_X2 FILLER_29_41 ();
 FILLCELL_X1 FILLER_29_43 ();
 FILLCELL_X4 FILLER_29_76 ();
 FILLCELL_X2 FILLER_29_80 ();
 FILLCELL_X1 FILLER_29_82 ();
 FILLCELL_X1 FILLER_29_91 ();
 FILLCELL_X32 FILLER_29_128 ();
 FILLCELL_X2 FILLER_29_160 ();
 FILLCELL_X1 FILLER_29_162 ();
 FILLCELL_X1 FILLER_29_220 ();
 FILLCELL_X2 FILLER_29_228 ();
 FILLCELL_X2 FILLER_29_237 ();
 FILLCELL_X8 FILLER_29_252 ();
 FILLCELL_X4 FILLER_29_260 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X16 FILLER_30_33 ();
 FILLCELL_X2 FILLER_30_49 ();
 FILLCELL_X1 FILLER_30_51 ();
 FILLCELL_X4 FILLER_30_74 ();
 FILLCELL_X2 FILLER_30_78 ();
 FILLCELL_X1 FILLER_30_80 ();
 FILLCELL_X32 FILLER_30_123 ();
 FILLCELL_X16 FILLER_30_155 ();
 FILLCELL_X8 FILLER_30_171 ();
 FILLCELL_X4 FILLER_30_179 ();
 FILLCELL_X2 FILLER_30_183 ();
 FILLCELL_X1 FILLER_30_185 ();
 FILLCELL_X2 FILLER_30_211 ();
 FILLCELL_X1 FILLER_30_231 ();
 FILLCELL_X8 FILLER_30_252 ();
 FILLCELL_X4 FILLER_30_260 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X8 FILLER_31_33 ();
 FILLCELL_X2 FILLER_31_41 ();
 FILLCELL_X8 FILLER_31_63 ();
 FILLCELL_X2 FILLER_31_71 ();
 FILLCELL_X1 FILLER_31_73 ();
 FILLCELL_X4 FILLER_31_98 ();
 FILLCELL_X32 FILLER_31_104 ();
 FILLCELL_X32 FILLER_31_136 ();
 FILLCELL_X16 FILLER_31_168 ();
 FILLCELL_X8 FILLER_31_184 ();
 FILLCELL_X1 FILLER_31_192 ();
 FILLCELL_X8 FILLER_31_196 ();
 FILLCELL_X2 FILLER_31_204 ();
 FILLCELL_X8 FILLER_31_208 ();
 FILLCELL_X1 FILLER_31_216 ();
 FILLCELL_X16 FILLER_31_237 ();
 FILLCELL_X8 FILLER_31_253 ();
 FILLCELL_X2 FILLER_31_261 ();
 FILLCELL_X1 FILLER_31_263 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X8 FILLER_32_193 ();
 FILLCELL_X2 FILLER_32_201 ();
 FILLCELL_X32 FILLER_32_223 ();
 FILLCELL_X8 FILLER_32_255 ();
 FILLCELL_X1 FILLER_32_263 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X4 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_168 ();
 FILLCELL_X32 FILLER_33_200 ();
 FILLCELL_X32 FILLER_33_232 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X16 FILLER_34_97 ();
 FILLCELL_X4 FILLER_34_113 ();
 FILLCELL_X1 FILLER_34_120 ();
 FILLCELL_X32 FILLER_34_124 ();
 FILLCELL_X32 FILLER_34_156 ();
 FILLCELL_X32 FILLER_34_188 ();
 FILLCELL_X32 FILLER_34_220 ();
 FILLCELL_X8 FILLER_34_252 ();
 FILLCELL_X4 FILLER_34_260 ();
endmodule
