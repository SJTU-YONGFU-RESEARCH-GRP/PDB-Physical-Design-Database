
* cell parameterized_freq_divider
* pin divide_value[13]
* pin duty_cycle[0]
* pin duty_cycle[4]
* pin duty_cycle[5]
* pin divide_value[2]
* pin duty_cycle[6]
* pin divide_value[4]
* pin divide_value[0]
* pin divide_value[1]
* pin divide_value[14]
* pin divide_value[7]
* pin divide_value[15]
* pin divide_value[12]
* pin divide_value[8]
* pin divide_value[9]
* pin divide_value[11]
* pin divide_value[10]
* pin clk_in
* pin rst_n
* pin enable
* pin clk_out
* pin divide_value[5]
* pin divide_value[3]
* pin divide_value[6]
* pin duty_cycle[3]
* pin duty_cycle[1]
* pin duty_cycle[2]
.SUBCKT parameterized_freq_divider 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
+ 19 20 21 1261 1404 1412 2463 2464 2465
* net 1 divide_value[13]
* net 2 duty_cycle[0]
* net 3 duty_cycle[4]
* net 4 duty_cycle[5]
* net 5 divide_value[2]
* net 6 duty_cycle[6]
* net 7 divide_value[4]
* net 8 divide_value[0]
* net 9 divide_value[1]
* net 10 divide_value[14]
* net 11 divide_value[7]
* net 12 divide_value[15]
* net 13 divide_value[12]
* net 14 divide_value[8]
* net 15 divide_value[9]
* net 16 divide_value[11]
* net 17 divide_value[10]
* net 18 clk_in
* net 19 rst_n
* net 20 enable
* net 21 clk_out
* net 1261 divide_value[5]
* net 1404 divide_value[3]
* net 1412 divide_value[6]
* net 2463 duty_cycle[3]
* net 2464 duty_cycle[1]
* net 2465 duty_cycle[2]
* cell instance $3 r0 *1 781.54,2.72
X$3 48 1 29 27 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $6 r0 *1 785.22,2.72
X$6 48 2 29 37 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $8 r0 *1 794.42,2.72
X$8 48 3 29 22 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $12 r0 *1 791.66,2.72
X$12 48 4 29 24 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $15 r0 *1 797.18,2.72
X$15 29 35 5 48 48 29 sky130_fd_sc_hd__dlymetal6s2s_1
* cell instance $18 m0 *1 799.02,8.16
X$18 48 6 29 63 48 29 sky130_fd_sc_hd__buf_2
* cell instance $21 r0 *1 802.24,2.72
X$21 48 7 34 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $24 r0 *1 807.3,2.72
X$24 48 8 29 32 48 29 sky130_fd_sc_hd__buf_2
* cell instance $27 r0 *1 809.14,2.72
X$27 29 31 9 48 48 29 sky130_fd_sc_hd__dlymetal6s2s_1
* cell instance $30 r0 *1 822.94,2.72
X$30 48 10 29 26 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $33 m0 *1 820.64,8.16
X$33 48 11 70 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $36 r0 *1 820.18,2.72
X$36 48 12 29 39 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $39 m0 *1 824.78,8.16
X$39 48 13 29 40 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $42 m0 *1 823.4,8.16
X$42 48 14 44 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $45 m0 *1 822.02,8.16
X$45 48 15 71 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $48 r0 *1 827.08,2.72
X$48 48 16 45 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $50 m0 *1 829.84,8.16
X$50 48 17 72 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $54 r0 *1 836.74,2.72
X$54 48 18 48 29 46 29 sky130_fd_sc_hd__buf_4
* cell instance $57 r0 *1 845.02,2.72
X$57 29 19 47 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $60 r0 *1 843.64,2.72
X$60 48 20 370 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $63 r0 *1 849.16,2.72
X$63 48 30 21 29 48 29 sky130_fd_sc_hd__clkbuf_1
* cell instance $78 r0 *1 802.24,84.32
X$78 48 22 462 968 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $80 r0 *1 754.4,13.6
X$80 48 22 39 137 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $82 m0 *1 750.72,8.16
X$82 48 22 26 50 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $84 m0 *1 766.82,8.16
X$84 48 22 40 57 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $87 r0 *1 763.6,2.72
X$87 48 22 27 134 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $89 m0 *1 795.34,78.88
X$89 48 22 206 23 791 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $91 m0 *1 790.28,89.76
X$91 48 22 440 1000 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $97 m0 *1 802.24,29.92
X$97 48 22 29 129 48 29 sky130_fd_sc_hd__buf_2
* cell instance $115 r0 *1 811.9,78.88
X$115 48 23 576 880 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $117 m0 *1 795.8,106.08
X$117 48 23 462 1356 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $121 r0 *1 2.3,845.92
X$121 29 2465 23 48 48 29 sky130_fd_sc_hd__buf_16
* cell instance $124 m0 *1 810.52,106.08
X$124 48 23 608 1243 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $126 m0 *1 756.24,19.04
X$126 48 23 26 141 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $128 m0 *1 761.76,8.16
X$128 48 23 39 86 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $132 r0 *1 813.28,13.6
X$132 48 23 29 68 48 29 sky130_fd_sc_hd__buf_2
* cell instance $134 m0 *1 778.32,8.16
X$134 48 23 27 91 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $151 m0 *1 747.5,19.04
X$151 48 24 26 150 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $153 m0 *1 748.42,8.16
X$153 48 24 27 81 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $155 m0 *1 764.52,8.16
X$155 48 24 40 56 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $157 m0 *1 751.64,24.48
X$157 48 24 39 176 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $159 m0 *1 792.58,78.88
X$159 48 24 462 844 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $161 r0 *1 794.42,73.44
X$161 48 24 781 806 29 352 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $163 r0 *1 790.28,29.92
X$163 48 24 29 77 48 29 sky130_fd_sc_hd__buf_2
* cell instance $167 m0 *1 776.02,8.16
X$167 48 24 28 41 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $172 r0 *1 754.86,2.72
X$172 48 25 48 29 36 29 sky130_fd_sc_hd__inv_1
* cell instance $174 r0 *1 760.84,8.16
X$174 29 53 25 38 86 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $191 r0 *1 761.3,2.72
X$191 48 33 26 38 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $193 r0 *1 750.72,24.48
X$193 48 63 26 221 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $196 m0 *1 822.02,19.04
X$196 48 26 84 145 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $199 m0 *1 822.48,24.48
X$199 48 26 84 146 191 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $201 m0 *1 824.32,24.48
X$201 48 180 26 48 182 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $203 m0 *1 793.5,13.6
X$203 48 101 26 99 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $207 r0 *1 783.38,8.16
X$207 48 102 26 42 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $224 r0 *1 758.08,19.04
X$224 48 206 27 156 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $227 m0 *1 750.72,19.04
X$227 48 63 27 152 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $231 r0 *1 823.4,8.16
X$231 48 45 72 27 40 84 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $233 r0 *1 822.48,19.04
X$233 48 175 27 174 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $235 r0 *1 804.08,13.6
X$235 48 102 27 65 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $237 m0 *1 793.96,19.04
X$237 48 101 27 128 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $248 m0 *1 799.48,29.92
X$248 48 101 28 244 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $250 r0 *1 826.16,8.16
X$250 48 45 29 28 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $253 m0 *1 823.4,19.04
X$253 48 146 72 28 40 29 175 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $256 r0 *1 804.08,2.72
X$256 48 33 28 64 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $258 m0 *1 811.9,8.16
X$258 48 68 28 87 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $261 r0 *1 776.94,19.04
X$261 48 143 28 142 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $264 r0 *1 783.84,13.6
X$264 48 129 28 116 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $268 r0 *1 810.06,13.6
X$268 48 102 28 120 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $270 m0 *1 826.16,29.92
X$270 48 255 28 254 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $272 m0 *1 821.56,29.92
X$272 48 28 67 212 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $5368 m0 *1 753.02,8.16
X$5368 48 33 39 51 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $5369 m0 *1 754.4,8.16
X$5369 29 107 54 53 52 154 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $5372 m0 *1 769.58,8.16
X$5372 29 133 58 57 41 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $5381 m0 *1 783.84,8.16
X$5381 29 59 61 93 43 60 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $5382 m0 *1 791.2,8.16
X$5382 29 117 119 99 62 166 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $5388 m0 *1 802.24,8.16
X$5388 29 43 66 64 65 89 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $5389 m0 *1 809.6,8.16
X$5389 48 33 67 69 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $5400 m0 *1 839.04,8.16
X$5400 29 47 30 46 375 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $6396 r0 *1 745.2,8.16
X$6396 48 49 48 29 83 29 sky130_fd_sc_hd__inv_1
* cell instance $6398 r0 *1 746.58,8.16
X$6398 29 49 82 50 81 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $6404 m0 *1 750.72,13.6
X$6404 48 105 48 29 104 29 sky130_fd_sc_hd__inv_1
* cell instance $6405 r0 *1 751.18,8.16
X$6405 29 105 106 51 83 36 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6407 m0 *1 753.02,13.6
X$6407 48 107 48 29 108 29 sky130_fd_sc_hd__inv_1
* cell instance $6408 m0 *1 754.4,13.6
X$6408 29 153 136 106 85 108 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6409 r0 *1 758.54,8.16
X$6409 48 73 48 29 85 29 sky130_fd_sc_hd__inv_1
* cell instance $6413 m0 *1 763.6,13.6
X$6413 48 54 48 29 55 29 sky130_fd_sc_hd__inv_1
* cell instance $6416 m0 *1 765.9,13.6
X$6416 29 109 132 110 112 74 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6417 r0 *1 766.36,8.16
X$6417 29 157 160 55 58 111 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6426 m0 *1 775.56,13.6
X$6426 48 113 48 29 74 29 sky130_fd_sc_hd__inv_1
* cell instance $6427 r0 *1 776.02,8.16
X$6427 29 113 60 42 91 90 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6429 m0 *1 777.4,13.6
X$6429 48 33 40 90 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6431 m0 *1 780.62,13.6
X$6431 29 115 93 96 76 116 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6432 r0 *1 785.68,8.16
X$6432 48 101 39 96 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6433 m0 *1 787.98,13.6
X$6433 48 77 67 76 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6435 r0 *1 788.44,8.16
X$6435 29 75 97 100 98 61 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6437 m0 *1 791.2,13.6
X$6437 48 117 48 29 100 29 sky130_fd_sc_hd__inv_1
* cell instance $6443 r0 *1 797.18,8.16
X$6443 29 98 92 94 95 78 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6445 m0 *1 798.1,13.6
X$6445 48 119 48 29 95 29 sky130_fd_sc_hd__inv_1
* cell instance $6447 m0 *1 800.4,13.6
X$6447 48 66 48 29 94 29 sky130_fd_sc_hd__inv_1
* cell instance $6453 m0 *1 804.08,13.6
X$6453 48 68 40 89 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6455 r0 *1 805,8.16
X$6455 29 78 88 69 79 87 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6456 m0 *1 806.38,13.6
X$6456 48 88 48 29 121 29 sky130_fd_sc_hd__inv_1
* cell instance $6458 m0 *1 808.22,13.6
X$6458 29 123 118 122 120 80 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $6459 r0 *1 812.36,8.16
X$6459 48 102 40 79 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6462 m0 *1 815.58,13.6
X$6462 48 68 67 80 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $6465 m0 *1 818.34,13.6
X$6465 48 70 44 71 39 29 114 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $6467 m0 *1 820.64,13.6
X$6467 48 71 29 103 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $7827 r0 *1 742.44,13.6
X$7827 29 140 138 139 82 104 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $7836 r0 *1 749.8,13.6
X$7836 29 139 177 150 137 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $7838 m0 *1 753.94,19.04
X$7838 48 153 48 29 151 29 sky130_fd_sc_hd__inv_1
* cell instance $7841 m0 *1 758.54,19.04
X$7841 29 154 110 156 198 141 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $7844 r0 *1 761.3,13.6
X$7844 48 136 48 29 135 29 sky130_fd_sc_hd__inv_1
* cell instance $7846 r0 *1 763.14,13.6
X$7846 29 52 73 134 56 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $7847 m0 *1 765.9,19.04
X$7847 48 157 48 29 158 29 sky130_fd_sc_hd__inv_1
* cell instance $7849 r0 *1 767.74,13.6
X$7849 48 109 48 29 111 29 sky130_fd_sc_hd__inv_1
* cell instance $7851 r0 *1 770.04,13.6
X$7851 48 133 48 29 112 29 sky130_fd_sc_hd__inv_1
* cell instance $7854 m0 *1 772.8,19.04
X$7854 48 161 48 29 159 29 sky130_fd_sc_hd__inv_1
* cell instance $7862 r0 *1 776.48,13.6
X$7862 29 161 131 132 115 59 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $7867 r0 *1 786.6,13.6
X$7867 48 75 48 29 130 29 sky130_fd_sc_hd__inv_1
* cell instance $7872 r0 *1 789.82,13.6
X$7872 48 37 29 101 48 29 sky130_fd_sc_hd__buf_2
* cell instance $7876 m0 *1 792.58,19.04
X$7876 48 129 67 166 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $7877 r0 *1 793.5,13.6
X$7877 48 77 103 62 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $7879 r0 *1 795.34,13.6
X$7879 29 165 126 128 127 168 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $7880 m0 *1 796.26,19.04
X$7880 48 77 125 127 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $7881 m0 *1 798.56,19.04
X$7881 48 129 103 168 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $7888 r0 *1 802.7,13.6
X$7888 48 92 48 29 124 29 sky130_fd_sc_hd__inv_1
* cell instance $7890 r0 *1 806.38,13.6
X$7890 48 33 103 122 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $7893 m0 *1 809.6,19.04
X$7893 48 118 48 29 170 29 sky130_fd_sc_hd__inv_1
* cell instance $7902 r0 *1 820.18,13.6
X$7902 48 44 29 125 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $7904 m0 *1 820.64,19.04
X$7904 48 145 114 147 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $7906 r0 *1 823.86,13.6
X$7906 48 72 29 67 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $9267 m0 *1 747.04,24.48
X$9267 29 194 196 177 176 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $9273 r0 *1 749.34,19.04
X$9273 29 218 224 138 152 151 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9279 m0 *1 760.38,24.48
X$9279 48 178 39 198 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $9282 r0 *1 761.3,19.04
X$9282 29 155 225 135 199 158 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9286 m0 *1 765.9,24.48
X$9286 48 143 40 199 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $9289 m0 *1 769.12,24.48
X$9289 48 201 48 29 200 29 sky130_fd_sc_hd__inv_1
* cell instance $9290 r0 *1 769.58,19.04
X$9290 29 201 162 160 142 159 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9298 m0 *1 776.94,24.48
X$9298 29 231 233 131 163 130 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9300 r0 *1 780.16,19.04
X$9300 48 143 67 163 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $9303 m0 *1 784.76,24.48
X$9303 29 275 204 235 164 97 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9309 r0 *1 790.74,19.04
X$9309 29 164 167 124 165 144 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9311 m0 *1 793.04,24.48
X$9311 29 238 197 240 203 242 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9313 r0 *1 799.02,19.04
X$9313 29 144 169 121 126 123 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9314 m0 *1 800.4,24.48
X$9314 48 169 48 29 202 29 sky130_fd_sc_hd__inv_1
* cell instance $9319 m0 *1 802.24,24.48
X$9319 29 179 195 170 197 248 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $9322 r0 *1 808.68,19.04
X$9322 48 33 125 246 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $9323 m0 *1 809.6,24.48
X$9323 48 68 103 193 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $9326 m0 *1 812.36,24.48
X$9326 48 102 67 249 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $9331 m0 *1 818.34,24.48
X$9331 48 192 84 180 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $9337 m0 *1 827.54,24.48
X$9337 48 189 188 181 29 48 190 29 sky130_fd_sc_hd__a21oi_1
* cell instance $9338 r0 *1 828,19.04
X$9338 48 190 148 149 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $9343 m0 *1 829.84,24.48
X$9343 48 186 40 48 187 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $9344 r0 *1 830.3,19.04
X$9344 29 148 173 172 174 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $9346 m0 *1 833.98,24.48
X$9346 29 185 184 183 182 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $9347 r0 *1 834.9,19.04
X$9347 48 173 149 185 48 171 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $10694 r0 *1 741.98,24.48
X$10694 29 213 214 194 221 140 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $10695 m0 *1 741.98,29.92
X$10695 29 270 215 220 196 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10697 m0 *1 747.04,29.92
X$10697 29 216 261 214 218 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10701 r0 *1 749.34,24.48
X$10701 48 217 48 29 219 29 sky130_fd_sc_hd__inv_1
* cell instance $10703 m0 *1 752.1,29.92
X$10703 29 222 223 205 224 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $10706 r0 *1 754.4,24.48
X$10706 48 63 39 220 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $10711 m0 *1 759,29.92
X$10711 48 206 29 33 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $10712 r0 *1 759,24.48
X$10712 48 155 48 29 205 29 sky130_fd_sc_hd__inv_1
* cell instance $10719 m0 *1 764.98,29.92
X$10719 29 279 207 226 200 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10721 r0 *1 766.82,24.48
X$10721 48 225 48 29 226 29 sky130_fd_sc_hd__inv_1
* cell instance $10723 m0 *1 769.58,29.92
X$10723 29 280 227 229 228 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10725 r0 *1 772.34,24.48
X$10725 48 162 48 29 229 29 sky130_fd_sc_hd__inv_1
* cell instance $10726 r0 *1 773.72,24.48
X$10726 48 231 48 29 228 29 sky130_fd_sc_hd__inv_1
* cell instance $10734 r0 *1 776.94,24.48
X$10734 48 63 29 143 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $10735 m0 *1 777.4,29.92
X$10735 48 208 48 29 232 29 sky130_fd_sc_hd__inv_1
* cell instance $10737 m0 *1 779.24,29.92
X$10737 48 209 48 29 230 29 sky130_fd_sc_hd__inv_1
* cell instance $10739 m0 *1 780.62,29.92
X$10739 29 208 209 167 237 236 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $10741 r0 *1 782.46,24.48
X$10741 48 233 48 29 234 29 sky130_fd_sc_hd__inv_1
* cell instance $10743 r0 *1 784.76,24.48
X$10743 48 143 103 235 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $10745 m0 *1 787.98,29.92
X$10745 48 210 48 29 236 29 sky130_fd_sc_hd__inv_1
* cell instance $10748 r0 *1 788.9,24.48
X$10748 29 210 239 202 238 179 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $10749 m0 *1 789.36,29.92
X$10749 48 143 125 237 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $10752 m0 *1 793.04,29.92
X$10752 48 101 40 240 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $10753 m0 *1 795.34,29.92
X$10753 48 129 125 242 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $10755 r0 *1 797.18,24.48
X$10755 29 241 290 211 243 245 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $10763 m0 *1 805,29.92
X$10763 48 178 29 102 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $10764 r0 *1 806.38,24.48
X$10764 48 195 48 29 211 29 sky130_fd_sc_hd__inv_1
* cell instance $10765 r0 *1 807.76,24.48
X$10765 29 248 252 246 249 193 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $10768 m0 *1 812.36,29.92
X$10768 48 252 48 29 250 29 sky130_fd_sc_hd__inv_1
* cell instance $10776 r0 *1 821.56,24.48
X$10776 48 191 39 257 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $10777 m0 *1 822.94,29.92
X$10777 48 67 146 255 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $10779 r0 *1 824.78,24.48
X$10779 29 258 251 256 257 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10780 m0 *1 824.78,29.92
X$10780 48 212 192 186 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $10784 r0 *1 829.38,24.48
X$10784 29 188 189 350 187 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $10786 m0 *1 829.84,29.92
X$10786 48 251 258 247 29 48 253 29 sky130_fd_sc_hd__a21oi_1
* cell instance $10791 r0 *1 836.28,24.48
X$10791 48 171 184 247 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $12138 r0 *1 742.44,29.92
X$12138 29 259 217 270 213 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $12142 m0 *1 747.04,35.36
X$12142 48 283 282 297 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $12143 r0 *1 747.04,29.92
X$12143 48 216 29 260 48 29 sky130_fd_sc_hd__buf_2
* cell instance $12147 m0 *1 748.42,35.36
X$12147 48 217 261 299 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $12148 r0 *1 748.88,29.92
X$12148 48 260 259 261 48 29 355 29 sky130_fd_sc_hd__o21ai_1
* cell instance $12149 m0 *1 749.8,35.36
X$12149 48 222 207 223 29 48 298 29 sky130_fd_sc_hd__a21o_1
* cell instance $12151 r0 *1 751.18,29.92
X$12151 48 260 223 261 29 48 262 29 sky130_fd_sc_hd__a21o_1
* cell instance $12152 m0 *1 752.56,35.36
X$12152 48 222 223 207 48 283 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $12154 r0 *1 755.78,29.92
X$12154 48 259 262 272 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $12155 m0 *1 755.78,35.36
X$12155 48 260 222 284 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $12158 r0 *1 757.62,29.92
X$12158 48 259 262 273 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $12159 m0 *1 758.08,35.36
X$12159 48 284 285 273 48 341 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $12161 m0 *1 759.92,35.36
X$12161 48 284 285 301 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $12166 m0 *1 761.76,35.36
X$12166 48 264 263 273 300 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $12168 r0 *1 762.22,29.92
X$12168 48 264 263 276 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $12169 m0 *1 763.6,35.36
X$12169 48 263 302 287 48 285 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $12170 r0 *1 763.6,29.92
X$12170 48 279 29 277 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $12171 m0 *1 766.36,35.36
X$12171 48 287 263 302 48 29 342 29 sky130_fd_sc_hd__o21ai_1
* cell instance $12172 r0 *1 766.36,29.92
X$12172 48 277 207 227 48 263 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $12173 m0 *1 768.2,35.36
X$12173 48 227 265 274 29 48 288 29 sky130_fd_sc_hd__a21oi_1
* cell instance $12176 r0 *1 770.5,29.92
X$12176 48 280 29 265 48 29 sky130_fd_sc_hd__buf_2
* cell instance $12177 m0 *1 770.5,35.36
X$12177 48 281 289 274 287 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $12186 r0 *1 774.64,29.92
X$12186 29 281 289 232 204 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $12189 m0 *1 779.7,35.36
X$12189 48 290 48 29 303 29 sky130_fd_sc_hd__inv_1
* cell instance $12190 r0 *1 780.16,29.92
X$12190 29 278 274 275 234 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $12192 m0 *1 782.92,35.36
X$12192 29 327 291 239 304 305 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $12197 m0 *1 790.28,35.36
X$12197 48 143 271 304 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $12201 r0 *1 793.5,29.92
X$12201 48 77 271 203 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $12203 r0 *1 795.8,29.92
X$12203 48 129 271 269 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $12204 m0 *1 796.26,35.36
X$12204 48 241 48 29 305 29 sky130_fd_sc_hd__inv_1
* cell instance $12206 r0 *1 798.1,29.92
X$12206 29 243 268 244 306 269 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $12207 m0 *1 799.48,35.36
X$12207 48 77 319 306 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $12215 r0 *1 805.46,29.92
X$12215 29 245 379 250 268 307 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $12216 m0 *1 805.46,35.36
X$12216 48 33 271 308 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $12217 m0 *1 807.76,35.36
X$12217 29 307 292 308 267 309 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $12218 r0 *1 812.82,29.92
X$12218 48 102 103 267 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $12224 r0 *1 817.42,29.92
X$12224 48 70 29 271 48 29 sky130_fd_sc_hd__buf_2
* cell instance $12226 r0 *1 819.26,29.92
X$12226 48 125 70 452 266 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $12228 m0 *1 821.1,35.36
X$12228 48 266 103 312 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $12230 r0 *1 821.56,29.92
X$12230 48 266 103 146 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $12234 m0 *1 827.08,35.36
X$12234 48 294 293 181 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $12240 m0 *1 829.84,35.36
X$12240 29 295 293 311 254 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $12243 r0 *1 833.52,29.92
X$12243 29 47 183 46 381 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $12245 m0 *1 835.36,35.36
X$12245 29 47 172 46 310 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $13587 m0 *1 743.36,40.8
X$13587 48 260 297 353 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $13589 m0 *1 744.74,40.8
X$13589 48 215 354 339 48 29 356 29 sky130_fd_sc_hd__o21ai_1
* cell instance $13590 r0 *1 745.2,35.36
X$13590 48 299 48 29 313 29 sky130_fd_sc_hd__inv_1
* cell instance $13593 m0 *1 747.04,40.8
X$13593 29 219 355 283 339 299 282 48 48 29 sky130_fd_sc_hd__a32oi_4
* cell instance $13597 r0 *1 747.5,35.36
X$13597 48 215 313 298 314 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $13599 r0 *1 750.26,35.36
X$13599 48 222 277 282 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $13601 r0 *1 752.1,35.36
X$13601 48 277 338 337 336 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $13603 r0 *1 754.4,35.36
X$13603 48 474 436 335 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $13604 r0 *1 755.78,35.36
X$13604 29 29 315 357 340 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $13605 m0 *1 757.16,40.8
X$13605 29 342 358 333 286 276 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $13607 r0 *1 758.54,35.36
X$13607 48 316 288 317 48 29 334 29 sky130_fd_sc_hd__o21ai_1
* cell instance $13609 r0 *1 760.84,35.36
X$13609 29 315 333 286 276 301 259 48 48 29 sky130_fd_sc_hd__o311ai_2
* cell instance $13610 m0 *1 764.98,40.8
X$13610 48 332 29 348 48 29 sky130_fd_sc_hd__buf_2
* cell instance $13611 r0 *1 766.82,35.36
X$13611 48 278 274 277 265 302 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $13612 m0 *1 766.82,40.8
X$13612 48 265 278 316 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $13613 m0 *1 768.2,40.8
X$13613 48 345 29 360 48 29 sky130_fd_sc_hd__buf_2
* cell instance $13614 r0 *1 769.58,35.36
X$13614 48 278 274 289 48 264 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $13615 m0 *1 770.04,40.8
X$13615 48 289 281 318 29 48 317 29 sky130_fd_sc_hd__a21oi_1
* cell instance $13616 m0 *1 771.88,40.8
X$13616 48 347 330 331 29 48 343 29 sky130_fd_sc_hd__a21oi_1
* cell instance $13618 r0 *1 773.26,35.36
X$13618 48 281 278 289 48 29 331 29 sky130_fd_sc_hd__o21ai_1
* cell instance $13624 m0 *1 774.64,40.8
X$13624 48 330 331 346 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $13626 r0 *1 775.56,35.36
X$13626 48 274 48 29 330 29 sky130_fd_sc_hd__inv_1
* cell instance $13627 m0 *1 776.02,40.8
X$13627 29 362 468 303 364 363 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $13628 r0 *1 776.94,35.36
X$13628 29 332 318 230 329 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $13629 r0 *1 781.54,35.36
X$13629 48 327 48 29 329 29 sky130_fd_sc_hd__inv_1
* cell instance $13633 r0 *1 784.3,35.36
X$13633 48 291 48 29 328 29 sky130_fd_sc_hd__inv_1
* cell instance $13634 m0 *1 784.3,40.8
X$13634 29 411 369 326 365 367 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $13635 r0 *1 785.68,35.36
X$13635 48 101 67 326 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13638 r0 *1 788.9,35.36
X$13638 48 129 319 367 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13640 m0 *1 791.66,40.8
X$13640 29 366 371 325 369 372 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $13651 r0 *1 802.7,35.36
X$13651 48 292 48 29 325 29 sky130_fd_sc_hd__inv_1
* cell instance $13652 r0 *1 804.08,35.36
X$13652 48 102 125 324 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13653 m0 *1 804.08,40.8
X$13653 48 33 319 376 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13655 m0 *1 806.38,40.8
X$13655 48 68 271 377 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13657 r0 *1 808.68,35.36
X$13657 48 68 125 309 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $13661 m0 *1 810.98,40.8
X$13661 48 379 48 29 380 29 sky130_fd_sc_hd__inv_1
* cell instance $13668 r0 *1 818.34,35.36
X$13668 29 192 103 125 271 323 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $13671 m0 *1 821.1,40.8
X$13671 29 384 387 390 322 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $13672 r0 *1 822.94,35.36
X$13672 48 192 67 322 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $13673 m0 *1 825.7,40.8
X$13673 48 388 384 386 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $13675 r0 *1 826.62,35.36
X$13675 48 387 386 295 48 294 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $13677 r0 *1 828.46,35.36
X$13677 29 320 296 389 253 48 48 29 sky130_fd_sc_hd__o21bai_4
* cell instance $13685 m0 *1 831.22,40.8
X$13685 48 385 172 378 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $13686 m0 *1 834.44,40.8
X$13686 48 296 382 381 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $13687 r0 *1 835.36,35.36
X$13687 48 296 378 310 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $13691 m0 *1 837.2,40.8
X$13691 48 320 351 352 29 48 375 29 sky130_fd_sc_hd__a21oi_1
* cell instance $13692 r0 *1 838.58,35.36
X$13692 48 296 374 321 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $13696 m0 *1 840.42,40.8
X$13696 48 351 373 370 48 320 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $13701 r0 *1 843.64,35.36
X$13701 29 47 350 46 321 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $15034 m0 *1 732.78,46.24
X$15034 29 391 428 426 392 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $15040 m0 *1 740.6,46.24
X$15040 48 392 401 414 48 29 431 29 sky130_fd_sc_hd__o21ai_1
* cell instance $15042 m0 *1 742.44,46.24
X$15042 29 391 260 298 395 393 394 48 48 29 sky130_fd_sc_hd__o311a_2
* cell instance $15043 r0 *1 742.9,40.8
X$15043 48 353 260 298 29 48 394 29 sky130_fd_sc_hd__a21oi_1
* cell instance $15044 r0 *1 744.74,40.8
X$15044 29 313 354 215 298 334 339 48 48 29 sky130_fd_sc_hd__o311ai_0
* cell instance $15046 m0 *1 747.04,46.24
X$15046 29 277 393 222 260 337 338 48 48 29 sky130_fd_sc_hd__o2111ai_2
* cell instance $15050 r0 *1 747.96,40.8
X$15050 29 339 457 335 215 403 356 48 48 29 sky130_fd_sc_hd__a311oi_4
* cell instance $15051 m0 *1 752.56,46.24
X$15051 29 358 222 404 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $15052 r0 *1 757.62,40.8
X$15052 48 340 315 48 407 29 29 sky130_fd_sc_hd__and2_2
* cell instance $15054 r0 *1 760.84,40.8
X$15054 29 340 333 286 300 272 341 48 48 29 sky130_fd_sc_hd__o311a_1
* cell instance $15055 m0 *1 762.68,46.24
X$15055 48 316 397 416 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $15056 m0 *1 764.06,46.24
X$15056 29 343 477 346 486 265 417 48 48 29 sky130_fd_sc_hd__a32oi_4
* cell instance $15058 r0 *1 765.44,40.8
X$15058 48 398 344 359 343 48 396 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $15059 r0 *1 768.66,40.8
X$15059 48 265 346 344 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $15060 r0 *1 770.04,40.8
X$15060 48 318 348 361 48 29 333 29 sky130_fd_sc_hd__a21o_2
* cell instance $15061 r0 *1 773.26,40.8
X$15061 48 318 348 349 29 48 410 29 sky130_fd_sc_hd__a21oi_1
* cell instance $15066 m0 *1 774.64,46.24
X$15066 29 29 410 417 264 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $15067 r0 *1 775.1,40.8
X$15067 29 345 349 328 362 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $15070 m0 *1 778.32,46.24
X$15070 48 143 319 364 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $15072 r0 *1 780.62,40.8
X$15072 29 363 409 380 411 366 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $15077 m0 *1 787.52,46.24
X$15077 29 446 444 408 445 399 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $15080 r0 *1 789.36,40.8
X$15080 48 77 368 365 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $15084 r0 *1 795.8,40.8
X$15084 48 371 48 29 408 29 sky130_fd_sc_hd__inv_1
* cell instance $15085 m0 *1 796.72,46.24
X$15085 48 101 103 443 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $15095 r0 *1 802.24,40.8
X$15095 29 372 441 376 324 377 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $15099 m0 *1 805.46,46.24
X$15099 48 441 48 29 442 29 sky130_fd_sc_hd__inv_1
* cell instance $15102 m0 *1 810.52,46.24
X$15102 48 31 29 440 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $15108 m0 *1 816.04,46.24
X$15108 29 2466 405 439 31 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $15109 r0 *1 816.04,40.8
X$15109 29 2468 406 32 31 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $15110 r0 *1 820.64,40.8
X$15110 48 405 406 147 383 351 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $15112 r0 *1 823.4,40.8
X$15112 48 147 351 323 48 29 389 29 sky130_fd_sc_hd__o21ai_1
* cell instance $15116 m0 *1 825.7,46.24
X$15116 48 400 438 437 29 48 388 29 sky130_fd_sc_hd__a21oi_1
* cell instance $15118 r0 *1 826.62,40.8
X$15118 29 438 400 421 312 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $15126 m0 *1 831.22,46.24
X$15126 48 350 48 29 435 29 sky130_fd_sc_hd__inv_1
* cell instance $15128 r0 *1 832.14,40.8
X$15128 48 434 183 382 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $15129 m0 *1 832.6,46.24
X$15129 48 424 423 402 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $15130 m0 *1 833.98,46.24
X$15130 29 47 311 46 433 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $15131 r0 *1 835.36,40.8
X$15131 48 402 350 374 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $15134 m0 *1 843.18,46.24
X$15134 48 421 311 350 390 29 432 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $16466 m0 *1 727.72,51.68
X$16466 48 403 407 426 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16467 r0 *1 729.56,46.24
X$16467 48 426 453 412 29 48 600 29 sky130_fd_sc_hd__o21a_2
* cell instance $16468 m0 *1 730.02,51.68
X$16468 48 487 493 447 48 453 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $16470 m0 *1 732.32,51.68
X$16470 29 429 490 489 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $16473 r0 *1 733.7,46.24
X$16473 48 391 404 413 427 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $16475 r0 *1 736.46,46.24
X$16475 29 277 395 429 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $16476 m0 *1 742.44,51.68
X$16476 48 391 404 413 491 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $16477 m0 *1 744.28,51.68
X$16477 48 491 528 473 545 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $16480 m0 *1 747.04,51.68
X$16480 29 401 260 298 395 393 394 48 48 29 sky130_fd_sc_hd__o311ai_2
* cell instance $16485 r0 *1 747.96,46.24
X$16485 48 391 404 588 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16487 r0 *1 750.72,46.24
X$16487 48 456 48 29 413 29 sky130_fd_sc_hd__clkbuf_2
* cell instance $16489 m0 *1 753.02,51.68
X$16489 29 314 474 457 334 436 48 48 29 sky130_fd_sc_hd__and4b_1
* cell instance $16490 r0 *1 753.48,46.24
X$16490 29 415 448 336 396 458 48 48 29 sky130_fd_sc_hd__nor4b_2
* cell instance $16491 m0 *1 756.7,51.68
X$16491 48 475 416 334 29 48 337 29 sky130_fd_sc_hd__a21o_1
* cell instance $16492 r0 *1 759,46.24
X$16492 48 475 416 436 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $16493 m0 *1 759.46,51.68
X$16493 48 281 286 333 29 48 488 29 sky130_fd_sc_hd__o21a_2
* cell instance $16495 r0 *1 760.84,46.24
X$16495 48 476 404 415 414 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $16497 m0 *1 762.68,51.68
X$16497 48 348 281 397 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $16498 r0 *1 763.14,46.24
X$16498 48 338 337 277 48 458 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $16499 m0 *1 764.06,51.68
X$16499 29 486 477 359 265 448 417 48 48 29 sky130_fd_sc_hd__o41ai_4
* cell instance $16501 r0 *1 765.44,46.24
X$16501 48 449 397 317 29 498 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $16503 r0 *1 769.12,46.24
X$16503 48 360 348 417 265 29 398 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $16505 r0 *1 772.34,46.24
X$16505 48 348 360 265 347 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $16511 r0 *1 774.64,46.24
X$16511 48 349 450 418 48 29 361 29 sky130_fd_sc_hd__o21bai_1
* cell instance $16513 m0 *1 775.1,51.68
X$16513 48 349 360 478 29 48 449 29 sky130_fd_sc_hd__a21oi_1
* cell instance $16516 m0 *1 777.86,51.68
X$16516 29 500 478 521 469 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $16517 r0 *1 778.32,46.24
X$16517 48 360 48 29 450 29 sky130_fd_sc_hd__inv_1
* cell instance $16520 r0 *1 781.08,46.24
X$16520 48 468 48 29 469 29 sky130_fd_sc_hd__inv_1
* cell instance $16523 m0 *1 783.84,51.68
X$16523 29 520 485 409 451 518 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $16525 r0 *1 786.6,46.24
X$16525 48 143 368 451 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $16531 m0 *1 792.58,51.68
X$16531 48 101 125 563 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16534 m0 *1 794.88,51.68
X$16534 48 77 574 471 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16535 r0 *1 795.34,46.24
X$16535 29 445 470 443 471 472 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $16536 m0 *1 797.18,51.68
X$16536 48 129 368 472 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16543 m0 *1 802.24,51.68
X$16543 29 399 484 442 470 466 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $16545 r0 *1 803.62,46.24
X$16545 48 206 368 467 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16546 r0 *1 805.92,46.24
X$16546 29 466 463 467 465 464 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $16547 m0 *1 809.6,51.68
X$16547 48 68 319 464 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $16549 m0 *1 812.36,51.68
X$16549 48 368 34 319 539 383 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $16554 m0 *1 815.58,51.68
X$16554 48 440 462 383 452 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $16558 m0 *1 819.72,51.68
X$16558 48 461 125 459 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $16559 r0 *1 820.64,46.24
X$16559 48 271 323 461 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $16560 r0 *1 822.02,46.24
X$16560 29 460 419 480 459 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $16564 m0 *1 826.16,51.68
X$16564 48 256 48 29 483 29 sky130_fd_sc_hd__inv_1
* cell instance $16565 r0 *1 826.62,46.24
X$16565 48 420 419 437 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $16570 r0 *1 828.92,46.24
X$16570 48 311 48 29 422 29 sky130_fd_sc_hd__inv_1
* cell instance $16572 m0 *1 829.84,51.68
X$16572 48 296 482 479 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $16573 r0 *1 830.3,46.24
X$16573 48 311 390 421 423 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $16575 m0 *1 831.68,51.68
X$16575 48 172 48 29 455 29 sky130_fd_sc_hd__inv_1
* cell instance $16577 r0 *1 833.06,46.24
X$16577 48 423 435 455 424 29 434 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $16578 m0 *1 833.06,51.68
X$16578 29 47 256 46 479 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $16580 r0 *1 835.82,46.24
X$16580 48 454 422 425 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $16581 r0 *1 839.04,46.24
X$16581 48 296 425 433 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $16585 m0 *1 842.72,51.68
X$16585 48 480 183 256 172 29 481 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $16587 r0 *1 843.64,46.24
X$16587 48 432 481 430 634 29 48 373 29 sky130_fd_sc_hd__and4_1
* cell instance $17648 r0 *1 717.14,51.68
X$17648 29 525 526 507 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $17652 r0 *1 727.26,51.68
X$17652 48 404 413 511 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $17654 r0 *1 730.48,51.68
X$17654 48 489 527 512 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $17656 r0 *1 733.24,51.68
X$17656 29 490 429 513 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $17657 r0 *1 743.36,51.68
X$17657 48 487 447 392 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $17658 r0 *1 744.74,51.68
X$17658 48 413 392 404 401 29 48 473 29 sky130_fd_sc_hd__and4_1
* cell instance $17662 r0 *1 747.96,51.68
X$17662 48 494 404 413 492 48 547 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $17663 r0 *1 750.26,51.68
X$17663 29 29 493 514 447 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $17664 r0 *1 752.56,51.68
X$17664 29 395 337 474 48 48 29 sky130_fd_sc_hd__nand2b_2
* cell instance $17666 r0 *1 756.24,51.68
X$17666 29 396 525 448 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $17668 r0 *1 760.84,51.68
X$17668 48 412 495 496 643 29 48 29 sky130_fd_sc_hd__nand3b_1
* cell instance $17669 r0 *1 763.6,51.68
X$17669 48 278 531 498 29 48 529 29 sky130_fd_sc_hd__o21a_2
* cell instance $17670 r0 *1 766.82,51.68
X$17670 48 281 348 500 360 48 612 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $17671 r0 *1 769.12,51.68
X$17671 48 499 316 397 523 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $17672 r0 *1 770.96,51.68
X$17672 48 475 571 348 29 497 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $17673 r0 *1 774.18,51.68
X$17673 48 360 500 501 534 48 499 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $17677 r0 *1 776.48,51.68
X$17677 48 500 478 522 48 418 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $17679 r0 *1 780.16,51.68
X$17679 48 520 48 29 521 29 sky130_fd_sc_hd__inv_1
* cell instance $17683 r0 *1 784.76,51.68
X$17683 48 485 48 29 519 29 sky130_fd_sc_hd__inv_1
* cell instance $17685 r0 *1 786.6,51.68
X$17685 48 446 48 29 518 29 sky130_fd_sc_hd__inv_1
* cell instance $17688 r0 *1 789.36,51.68
X$17688 48 444 48 29 517 29 sky130_fd_sc_hd__inv_1
* cell instance $17697 r0 *1 804.08,51.68
X$17697 48 484 48 29 516 29 sky130_fd_sc_hd__inv_1
* cell instance $17699 r0 *1 807.3,51.68
X$17699 48 102 271 465 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $17700 r0 *1 809.6,51.68
X$17700 48 463 48 29 515 29 sky130_fd_sc_hd__inv_1
* cell instance $17702 r0 *1 812.82,51.68
X$17702 48 34 29 574 48 29 sky130_fd_sc_hd__buf_2
* cell instance $17706 r0 *1 816.96,51.68
X$17706 48 462 48 29 439 29 sky130_fd_sc_hd__inv_1
* cell instance $17707 r0 *1 818.34,51.68
X$17707 48 452 271 48 510 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $17709 r0 *1 822.02,51.68
X$17709 48 509 556 508 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $17711 r0 *1 824.78,51.68
X$17711 48 554 508 460 48 420 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $17713 r0 *1 827.54,51.68
X$17713 48 502 483 482 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $17717 r0 *1 830.76,51.68
X$17717 48 183 172 385 502 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $17718 r0 *1 832.6,51.68
X$17718 48 423 504 435 503 29 385 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $17719 r0 *1 834.9,51.68
X$17719 48 504 503 505 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $17720 r0 *1 836.28,51.68
X$17720 48 390 421 505 454 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $17721 r0 *1 838.12,51.68
X$17721 48 505 421 506 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $18397 m0 *1 725.42,57.12
X$18397 48 413 404 527 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $18398 m0 *1 728.64,57.12
X$18398 29 527 544 489 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $18401 m0 *1 734.16,57.12
X$18401 48 404 413 586 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $18403 m0 *1 737.38,57.12
X$18403 29 512 602 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $18405 m0 *1 742.44,57.12
X$18405 29 545 546 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $18407 m0 *1 747.04,57.12
X$18407 29 491 548 528 473 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $18408 m0 *1 753.02,57.12
X$18408 48 549 29 447 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $18409 m0 *1 755.78,57.12
X$18409 29 488 476 529 530 550 48 48 29 sky130_fd_sc_hd__nor4_4
* cell instance $18410 m0 *1 763.6,57.12
X$18410 29 278 530 498 531 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $18411 m0 *1 769.58,57.12
X$18411 29 523 338 533 532 48 48 29 sky130_fd_sc_hd__a21boi_2
* cell instance $18414 m0 *1 774.64,57.12
X$18414 48 500 360 536 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $18416 m0 *1 776.48,57.12
X$18416 29 534 522 537 519 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $18418 m0 *1 782.46,57.12
X$18418 29 537 558 517 557 559 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $18419 m0 *1 789.82,57.12
X$18419 48 560 48 29 561 29 sky130_fd_sc_hd__inv_1
* cell instance $18421 m0 *1 791.66,57.12
X$18421 29 564 567 563 565 594 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $18426 m0 *1 803.16,57.12
X$18426 48 37 271 659 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $18429 m0 *1 809.6,57.12
X$18429 48 68 368 566 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $18434 m0 *1 818.8,57.12
X$18434 48 562 319 323 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $18435 m0 *1 821.1,57.12
X$18435 29 556 554 540 510 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $18436 m0 *1 825.7,57.12
X$18436 48 183 48 29 555 29 sky130_fd_sc_hd__inv_1
* cell instance $18440 m0 *1 829.84,57.12
X$18440 48 421 48 29 541 29 sky130_fd_sc_hd__inv_1
* cell instance $18442 m0 *1 831.68,57.12
X$18442 48 390 541 424 582 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $18443 m0 *1 833.98,57.12
X$18443 48 480 540 503 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $18444 m0 *1 835.36,57.12
X$18444 29 47 421 46 552 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $19095 r0 *1 716.68,57.12
X$19095 48 569 524 513 48 661 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $19096 r0 *1 718.52,57.12
X$19096 48 577 602 546 48 29 579 29 sky130_fd_sc_hd__o21ai_1
* cell instance $19100 r0 *1 720.36,57.12
X$19100 29 583 526 525 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $19101 r0 *1 726.34,57.12
X$19101 48 524 569 489 583 29 585 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $19102 r0 *1 728.64,57.12
X$19102 48 427 547 584 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19106 r0 *1 733.7,57.12
X$19106 29 586 543 428 511 48 48 29 sky130_fd_sc_hd__o21bai_4
* cell instance $19108 r0 *1 741.06,57.12
X$19108 29 447 525 487 476 48 490 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $19113 r0 *1 749.8,57.12
X$19113 48 403 357 590 493 624 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $19114 r0 *1 752.56,57.12
X$19114 29 415 476 404 391 48 412 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $19116 r0 *1 760.84,57.12
X$19116 29 529 530 551 48 48 29 sky130_fd_sc_hd__nor2_8
* cell instance $19117 r0 *1 768.2,57.12
X$19117 29 281 550 333 286 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $19118 r0 *1 774.18,57.12
X$19118 48 572 535 523 29 474 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $19122 r0 *1 777.4,57.12
X$19122 48 522 573 570 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $19123 r0 *1 778.78,57.12
X$19123 48 536 538 449 29 475 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $19124 r0 *1 782,57.12
X$19124 48 522 534 595 29 48 538 29 sky130_fd_sc_hd__a21oi_1
* cell instance $19126 r0 *1 784.3,57.12
X$19126 48 558 48 29 596 29 sky130_fd_sc_hd__inv_1
* cell instance $19127 r0 *1 785.68,57.12
X$19127 48 63 574 557 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19129 r0 *1 788.44,57.12
X$19129 29 559 560 516 564 575 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $19130 r0 *1 795.8,57.12
X$19130 48 77 576 565 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19132 r0 *1 798.56,57.12
X$19132 29 575 592 515 567 591 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $19136 r0 *1 805.92,57.12
X$19136 48 206 574 607 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19137 r0 *1 808.22,57.12
X$19137 48 178 319 589 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19138 r0 *1 810.52,57.12
X$19138 48 35 576 539 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $19149 r0 *1 830.76,57.12
X$19149 48 541 424 390 48 553 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $19150 r0 *1 832.6,57.12
X$19150 48 296 553 582 29 48 581 29 sky130_fd_sc_hd__a21oi_1
* cell instance $19154 r0 *1 837.66,57.12
X$19154 48 296 29 542 48 29 sky130_fd_sc_hd__buf_2
* cell instance $19155 r0 *1 839.5,57.12
X$19155 48 542 506 552 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $19156 r0 *1 840.88,57.12
X$19156 48 542 647 580 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $19826 m0 *1 714.84,62.56
X$19826 48 568 613 543 48 614 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $19827 m0 *1 716.68,62.56
X$19827 48 597 507 598 489 29 48 578 29 sky130_fd_sc_hd__a31oi_1
* cell instance $19829 m0 *1 719.44,62.56
X$19829 29 569 568 583 524 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $19830 m0 *1 725.42,62.56
X$19830 48 615 583 764 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $19831 m0 *1 728.64,62.56
X$19831 48 616 600 599 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $19832 m0 *1 730.94,62.56
X$19832 48 412 392 514 601 617 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $19834 m0 *1 734.16,62.56
X$19834 29 639 618 619 602 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $19835 m0 *1 740.14,62.56
X$19835 29 493 447 476 48 526 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $19838 m0 *1 747.5,62.56
X$19838 29 528 588 496 413 495 412 48 48 29 sky130_fd_sc_hd__o2111a_1
* cell instance $19839 m0 *1 751.64,62.56
X$19839 48 765 549 415 476 29 48 456 29 sky130_fd_sc_hd__and4_1
* cell instance $19840 m0 *1 754.86,62.56
X$19840 29 493 403 549 407 48 495 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $19841 m0 *1 762.68,62.56
X$19841 48 359 477 360 29 593 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $19842 m0 *1 765.9,62.56
X$19842 29 531 612 570 532 603 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $19843 m0 *1 770.5,62.56
X$19843 48 348 534 611 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $19844 m0 *1 771.88,62.56
X$19844 48 499 532 533 29 48 571 29 sky130_fd_sc_hd__a21oi_1
* cell instance $19847 m0 *1 774.64,62.56
X$19847 48 532 570 603 48 610 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $19849 m0 *1 778.78,62.56
X$19849 29 609 595 653 596 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $19854 m0 *1 794.42,62.56
X$19854 48 129 574 594 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19856 m0 *1 797.64,62.56
X$19856 48 592 48 29 604 29 sky130_fd_sc_hd__inv_1
* cell instance $19857 m0 *1 799.02,62.56
X$19857 48 35 29 608 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $19859 m0 *1 802.24,62.56
X$19859 48 129 576 660 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $19862 m0 *1 805.92,62.56
X$19862 29 591 656 607 589 566 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $19864 m0 *1 813.74,62.56
X$19864 48 539 440 574 462 29 674 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $19867 m0 *1 818.34,62.56
X$19867 48 562 319 48 587 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $19868 m0 *1 821.56,62.56
X$19868 29 606 650 605 587 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $19875 m0 *1 832.14,62.56
X$19875 29 633 605 540 480 48 424 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $19877 m0 *1 837.2,62.56
X$19877 29 47 390 46 581 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $20528 r0 *1 712.08,62.56
X$20528 48 636 489 635 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $20529 r0 *1 713.46,62.56
X$20529 29 615 507 637 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $20533 r0 *1 723.58,62.56
X$20533 48 407 403 601 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $20534 r0 *1 725.88,62.56
X$20534 48 621 403 662 48 29 638 29 sky130_fd_sc_hd__o21ai_1
* cell instance $20535 r0 *1 727.72,62.56
X$20535 29 621 622 427 513 407 547 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $20536 r0 *1 730.94,62.56
X$20536 48 427 547 623 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $20539 r0 *1 733.24,62.56
X$20539 29 619 640 623 585 48 48 29 sky130_fd_sc_hd__and3_4
* cell instance $20540 r0 *1 737.38,62.56
X$20540 29 600 619 641 412 48 48 29 sky130_fd_sc_hd__o21bai_4
* cell instance $20541 r0 *1 744.28,62.56
X$20541 48 412 514 642 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $20542 r0 *1 745.66,62.56
X$20542 29 496 495 414 431 643 48 618 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $20546 r0 *1 755.32,62.56
X$20546 48 590 625 391 48 494 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $20547 r0 *1 757.16,62.56
X$20547 48 626 593 627 497 29 48 549 29 sky130_fd_sc_hd__and4_1
* cell instance $20549 r0 *1 760.84,62.56
X$20549 48 497 627 29 645 48 29 sky130_fd_sc_hd__and2_4
* cell instance $20550 r0 *1 764.06,62.56
X$20550 29 646 648 359 628 682 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $20551 r0 *1 771.42,62.56
X$20551 48 348 475 571 627 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $20552 r0 *1 773.72,62.56
X$20552 48 522 595 535 603 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $20556 r0 *1 775.56,62.56
X$20556 48 611 536 630 716 48 629 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $20557 r0 *1 778.78,62.56
X$20557 48 595 48 29 630 29 sky130_fd_sc_hd__inv_1
* cell instance $20558 r0 *1 780.16,62.56
X$20558 48 534 595 501 48 573 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $20559 r0 *1 782.92,62.56
X$20559 48 752 29 652 48 29 sky130_fd_sc_hd__buf_2
* cell instance $20560 r0 *1 784.76,62.56
X$20560 48 63 576 680 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $20566 r0 *1 796.26,62.56
X$20566 48 77 440 655 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $20567 r0 *1 798.56,62.56
X$20567 48 77 608 657 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $20568 r0 *1 800.86,62.56
X$20568 29 677 675 659 657 660 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $20574 r0 *1 809.6,62.56
X$20574 48 656 48 29 658 29 sky130_fd_sc_hd__inv_1
* cell instance $20578 r0 *1 816.04,62.56
X$20578 48 368 574 631 562 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $20581 r0 *1 822.94,62.56
X$20581 48 650 606 654 29 48 509 29 sky130_fd_sc_hd__a21oi_1
* cell instance $20583 r0 *1 826.62,62.56
X$20583 48 480 48 29 651 29 sky130_fd_sc_hd__inv_1
* cell instance $20588 r0 *1 831.68,62.56
X$20588 29 47 480 46 649 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $20591 r0 *1 843.64,62.56
X$20591 29 47 605 46 580 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $21254 m0 *1 707.48,68
X$21254 29 683 635 751 489 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $21255 m0 *1 713.46,68
X$21255 48 661 636 543 507 29 684 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $21256 m0 *1 716.22,68
X$21256 48 704 620 579 29 48 687 29 sky130_fd_sc_hd__and3_2
* cell instance $21258 m0 *1 719.44,68
X$21258 29 577 615 524 569 602 546 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $21259 m0 *1 729.56,68
X$21259 29 568 513 619 623 48 696 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $21260 m0 *1 737.38,68
X$21260 48 401 487 447 492 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $21261 m0 *1 739.22,68
X$21261 29 600 616 577 48 48 29 sky130_fd_sc_hd__nor2_8
* cell instance $21263 m0 *1 747.04,68
X$21263 29 685 642 357 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $21264 m0 *1 753.02,68
X$21264 29 686 357 403 493 487 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $21265 m0 *1 757.62,68
X$21265 29 626 497 593 627 48 625 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $21266 m0 *1 765.44,68
X$21266 48 360 359 477 626 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $21268 m0 *1 768.2,68
X$21268 29 663 418 682 477 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $21270 m0 *1 774.64,68
X$21270 29 663 595 664 501 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $21271 m0 *1 780.62,68
X$21271 48 609 29 501 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $21272 m0 *1 783.38,68
X$21272 48 665 48 29 681 29 sky130_fd_sc_hd__inv_1
* cell instance $21273 m0 *1 784.76,68
X$21273 29 653 679 561 680 666 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $21274 m0 *1 792.12,68
X$21274 48 679 48 29 678 29 sky130_fd_sc_hd__inv_1
* cell instance $21276 m0 *1 794.42,68
X$21276 29 666 676 604 677 667 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $21280 m0 *1 803.62,68
X$21280 29 667 699 658 675 717 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $21284 m0 *1 814.2,68
X$21284 48 674 368 673 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $21285 m0 *1 817.42,68
X$21285 29 672 668 644 673 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $21287 m0 *1 822.94,68
X$21287 48 669 668 654 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $21289 m0 *1 826.16,68
X$21289 48 632 651 670 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $21291 m0 *1 829.84,68
X$21291 48 540 605 633 632 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $21293 m0 *1 832.6,68
X$21293 48 542 670 649 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $21296 m0 *1 838.58,68
X$21296 48 633 605 647 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $21297 m0 *1 841.8,68
X$21297 48 671 605 540 644 29 634 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $21298 m0 *1 844.1,68
X$21298 29 47 706 46 707 48 48 29 sky130_fd_sc_hd__dfrtp_4
* cell instance $21941 r0 *1 701.96,68
X$21941 48 639 48 29 689 29 sky130_fd_sc_hd__inv_1
* cell instance $21942 r0 *1 703.34,68
X$21942 48 637 29 702 48 29 sky130_fd_sc_hd__buf_2
* cell instance $21944 r0 *1 705.64,68
X$21944 48 689 691 703 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $21945 r0 *1 707.02,68
X$21945 29 690 692 543 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $21946 r0 *1 713,68
X$21946 29 543 692 693 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $21951 r0 *1 723.58,68
X$21951 29 568 727 489 692 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $21952 r0 *1 729.56,68
X$21952 29 641 392 695 601 694 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $21954 r0 *1 733.24,68
X$21954 48 412 392 514 29 48 622 29 sky130_fd_sc_hd__a21oi_1
* cell instance $21956 r0 *1 735.54,68
X$21956 29 636 548 708 705 598 544 48 48 29 sky130_fd_sc_hd__o2111ai_4
* cell instance $21957 r0 *1 745.2,68
X$21957 29 697 710 551 447 493 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $21962 r0 *1 750.26,68
X$21962 29 624 686 616 412 625 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $21963 r0 *1 757.62,68
X$21963 48 593 626 48 712 29 29 sky130_fd_sc_hd__and2_2
* cell instance $21966 r0 *1 761.3,68
X$21966 29 625 496 590 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $21968 r0 *1 765.9,68
X$21968 29 646 663 648 286 629 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $21969 r0 *1 773.72,68
X$21969 29 29 534 682 500 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $21973 r0 *1 776.02,68
X$21973 48 652 664 501 48 716 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $21974 r0 *1 777.86,68
X$21974 29 500 610 698 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $21977 r0 *1 790.28,68
X$21977 48 143 608 722 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $21980 r0 *1 793.04,68
X$21980 48 719 48 29 721 29 sky130_fd_sc_hd__inv_1
* cell instance $21983 r0 *1 795.8,68
X$21983 48 63 178 37 723 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $21984 r0 *1 797.64,68
X$21984 48 63 48 29 720 29 sky130_fd_sc_hd__inv_1
* cell instance $21990 r0 *1 801.78,68
X$21990 48 699 48 29 718 29 sky130_fd_sc_hd__inv_1
* cell instance $21991 r0 *1 803.16,68
X$21991 48 129 608 742 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $21994 r0 *1 808.22,68
X$21994 29 717 715 777 740 739 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $21996 r0 *1 816.04,68
X$21996 48 576 608 714 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $21998 r0 *1 819.26,68
X$21998 48 799 773 672 48 669 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $22000 r0 *1 822.02,68
X$22000 48 390 48 29 713 29 sky130_fd_sc_hd__inv_1
* cell instance $22008 r0 *1 832.14,68
X$22008 48 605 48 29 711 29 sky130_fd_sc_hd__inv_1
* cell instance $22009 r0 *1 833.52,68
X$22009 29 47 540 46 735 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $22011 r0 *1 843.64,68
X$22011 48 701 542 709 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22012 r0 *1 845.02,68
X$22012 48 706 542 707 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22675 m0 *1 699.66,73.44
X$22675 48 687 688 702 48 29 768 29 sky130_fd_sc_hd__o21ai_1
* cell instance $22676 m0 *1 701.5,73.44
X$22676 48 639 683 749 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22677 m0 *1 702.88,73.44
X$22677 48 702 724 747 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22679 m0 *1 704.72,73.44
X$22679 48 689 725 637 821 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $22680 m0 *1 706.56,73.44
X$22680 48 691 750 693 29 48 724 29 sky130_fd_sc_hd__a21oi_1
* cell instance $22681 m0 *1 708.4,73.44
X$22681 48 635 489 751 48 29 750 29 sky130_fd_sc_hd__a21o_2
* cell instance $22682 m0 *1 711.62,73.44
X$22682 48 577 546 751 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22683 m0 *1 713,73.44
X$22683 48 636 543 578 704 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $22684 m0 *1 714.84,73.44
X$22684 48 584 619 578 48 29 763 29 sky130_fd_sc_hd__o21ai_1
* cell instance $22685 m0 *1 716.68,73.44
X$22685 48 447 403 357 493 48 694 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $22687 m0 *1 719.44,73.44
X$22687 29 725 704 620 579 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $22688 m0 *1 723.12,73.44
X$22688 48 543 568 636 513 48 620 29 29 sky130_fd_sc_hd__nand4b_1
* cell instance $22690 m0 *1 727.26,73.44
X$22690 29 727 577 546 602 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $22691 m0 *1 733.24,73.44
X$22691 29 754 824 780 708 726 48 755 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $22693 m0 *1 743.36,73.44
X$22693 29 597 728 695 710 697 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $22695 m0 *1 747.04,73.44
X$22695 29 728 695 710 524 697 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $22696 m0 *1 754.86,73.44
X$22696 29 496 756 710 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $22697 m0 *1 759,73.44
X$22697 29 550 710 488 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $22699 m0 *1 764.06,73.44
X$22699 29 534 784 729 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $22701 m0 *1 774.64,73.44
X$22701 29 29 753 48 572 535 48 sky130_fd_sc_hd__nor2_2
* cell instance $22702 m0 *1 776.94,73.44
X$22702 48 664 652 730 29 48 533 29 sky130_fd_sc_hd__a21oi_1
* cell instance $22704 m0 *1 779.7,73.44
X$22704 48 652 730 664 29 48 535 29 sky130_fd_sc_hd__a21o_1
* cell instance $22705 m0 *1 782.46,73.44
X$22705 29 752 664 678 681 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $22707 m0 *1 787.52,73.44
X$22707 29 665 748 676 722 721 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $22709 m0 *1 795.8,73.44
X$22709 48 745 791 723 29 48 781 29 sky130_fd_sc_hd__a21oi_1
* cell instance $22710 m0 *1 797.64,73.44
X$22710 48 720 731 746 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22714 m0 *1 802.24,73.44
X$22714 29 743 741 778 655 742 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $22715 m0 *1 809.6,73.44
X$22715 48 178 368 740 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $22716 m0 *1 811.9,73.44
X$22716 48 68 574 739 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $22718 m0 *1 815.12,73.44
X$22718 48 631 574 48 738 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $22719 m0 *1 818.34,73.44
X$22719 29 737 839 700 772 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $22720 m0 *1 822.94,73.44
X$22720 29 771 770 736 439 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $22721 m0 *1 827.54,73.44
X$22721 48 706 48 29 736 29 sky130_fd_sc_hd__inv_1
* cell instance $22725 m0 *1 830.3,73.44
X$22725 48 540 48 29 732 29 sky130_fd_sc_hd__inv_1
* cell instance $22727 m0 *1 832.14,73.44
X$22727 48 504 732 733 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $22728 m0 *1 835.36,73.44
X$22728 48 542 733 735 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $22729 m0 *1 836.74,73.44
X$22729 29 47 700 46 709 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $22730 m0 *1 846.4,73.44
X$22730 29 701 671 706 734 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $23368 r0 *1 690,73.44
X$23368 48 693 683 757 29 48 793 29 sky130_fd_sc_hd__a21oi_1
* cell instance $23369 r0 *1 691.84,73.44
X$23369 29 757 796 683 693 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $23373 r0 *1 694.14,73.44
X$23373 48 683 757 767 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $23374 r0 *1 695.52,73.44
X$23374 48 758 744 797 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $23376 r0 *1 697.82,73.44
X$23376 29 769 768 689 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $23377 r0 *1 703.8,73.44
X$23377 48 759 760 820 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $23379 r0 *1 705.64,73.44
X$23379 48 689 690 775 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $23380 r0 *1 707.02,73.44
X$23380 48 703 776 760 29 48 803 29 sky130_fd_sc_hd__a21oi_1
* cell instance $23381 r0 *1 708.86,73.44
X$23381 29 744 760 759 725 761 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $23382 r0 *1 712.08,73.44
X$23382 48 687 637 639 29 761 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $23383 r0 *1 715.3,73.44
X$23383 48 684 762 614 48 29 691 29 sky130_fd_sc_hd__o21bai_1
* cell instance $23384 r0 *1 718.06,73.44
X$23384 29 29 685 758 763 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $23388 r0 *1 720.36,73.44
X$23388 48 639 763 685 810 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $23389 r0 *1 722.2,73.44
X$23389 48 639 758 687 850 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $23390 r0 *1 724.04,73.44
X$23390 29 779 810 687 764 755 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $23391 r0 *1 728.64,73.44
X$23391 48 764 29 788 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $23396 r0 *1 733.7,73.44
X$23396 29 546 602 780 569 577 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $23398 r0 *1 741.52,73.44
X$23398 29 551 756 726 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $23402 r0 *1 751.64,73.44
X$23402 48 765 48 29 493 29 sky130_fd_sc_hd__buf_4
* cell instance $23403 r0 *1 754.4,73.44
X$23403 29 488 754 550 514 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $23405 r0 *1 760.84,73.44
X$23405 48 407 642 662 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $23406 r0 *1 762.22,73.44
X$23406 48 785 729 698 783 29 48 765 29 sky130_fd_sc_hd__and4_1
* cell instance $23407 r0 *1 765.44,73.44
X$23407 29 902 663 784 812 790 628 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $23411 r0 *1 775.1,73.44
X$23411 29 753 501 783 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $23412 r0 *1 785.22,73.44
X$23412 48 811 48 29 782 29 sky130_fd_sc_hd__buf_4
* cell instance $23415 r0 *1 788.9,73.44
X$23415 48 748 48 29 808 29 sky130_fd_sc_hd__inv_1
* cell instance $23418 r0 *1 797.64,73.44
X$23418 29 719 804 718 743 805 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $23422 r0 *1 805,73.44
X$23422 48 37 319 778 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $23424 r0 *1 807.76,73.44
X$23424 48 440 48 29 731 29 sky130_fd_sc_hd__inv_1
* cell instance $23426 r0 *1 810.06,73.44
X$23426 48 206 576 777 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $23428 r0 *1 812.82,73.44
X$23428 48 715 48 29 802 29 sky130_fd_sc_hd__inv_1
* cell instance $23429 r0 *1 814.2,73.44
X$23429 48 766 714 631 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $23432 r0 *1 816.96,73.44
X$23432 48 774 801 773 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $23433 r0 *1 819.26,73.44
X$23433 29 772 766 439 731 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $23434 r0 *1 823.86,73.44
X$23434 48 770 771 798 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $23446 r0 *1 845.48,73.44
X$23446 48 700 48 29 734 29 sky130_fd_sc_hd__inv_1
* cell instance $24103 m0 *1 687.7,78.88
X$24103 48 702 786 789 834 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $24104 m0 *1 689.54,78.88
X$24104 48 787 693 816 794 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $24106 m0 *1 691.84,78.88
X$24106 48 788 726 817 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $24107 m0 *1 693.22,78.88
X$24107 48 836 788 688 693 48 837 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $24108 m0 *1 695.52,78.88
X$24108 48 750 757 786 789 48 1010 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $24109 m0 *1 698.74,78.88
X$24109 48 702 759 760 29 48 800 29 sky130_fd_sc_hd__a21oi_1
* cell instance $24110 m0 *1 700.58,78.88
X$24110 48 639 747 758 48 955 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $24111 m0 *1 702.42,78.88
X$24111 48 749 693 788 725 639 822 29 48 29 sky130_fd_sc_hd__a32oi_1
* cell instance $24112 m0 *1 705.64,78.88
X$24112 29 760 759 725 858 761 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $24113 m0 *1 713.46,78.88
X$24113 48 810 725 788 29 48 807 29 sky130_fd_sc_hd__a21oi_1
* cell instance $24115 m0 *1 716.22,78.88
X$24115 48 597 598 513 507 29 613 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $24117 m0 *1 719.44,78.88
X$24117 29 755 639 637 787 48 809 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $24118 m0 *1 727.26,78.88
X$24118 48 851 29 787 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $24119 m0 *1 730.02,78.88
X$24119 29 883 617 638 696 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $24120 m0 *1 733.7,78.88
X$24120 48 599 29 636 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $24121 m0 *1 736.46,78.88
X$24121 29 705 780 1011 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $24123 m0 *1 747.04,78.88
X$24123 29 493 712 814 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $24124 m0 *1 757.16,78.88
X$24124 29 852 645 712 698 928 825 48 48 29 sky130_fd_sc_hd__a2111oi_2
* cell instance $24125 m0 *1 762.68,78.88
X$24125 29 590 813 783 698 729 48 48 29 sky130_fd_sc_hd__nand4b_2
* cell instance $24126 m0 *1 768.2,78.88
X$24126 48 830 501 652 782 48 812 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $24127 m0 *1 770.5,78.88
X$24127 29 29 652 628 501 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $24128 m0 *1 772.8,78.88
X$24128 48 849 826 848 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $24130 m0 *1 774.64,78.88
X$24130 29 790 730 829 782 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $24132 m0 *1 781.08,78.88
X$24132 29 847 572 868 846 48 48 29 sky130_fd_sc_hd__a21boi_2
* cell instance $24133 m0 *1 785.22,78.88
X$24133 29 811 730 808 845 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $24137 m0 *1 797.18,78.88
X$24137 48 720 791 745 48 806 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $24138 m0 *1 799.02,78.88
X$24138 48 804 48 29 843 29 sky130_fd_sc_hd__inv_1
* cell instance $24143 m0 *1 803.16,78.88
X$24143 29 805 842 802 741 884 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $24147 m0 *1 815.58,78.88
X$24147 29 801 799 792 738 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $24150 m0 *1 821.56,78.88
X$24150 48 737 798 839 29 48 841 29 sky130_fd_sc_hd__a21o_1
* cell instance $24156 m0 *1 830.76,78.88
X$24156 29 47 644 46 838 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $24157 m0 *1 839.96,78.88
X$24157 29 47 792 46 835 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $24158 m0 *1 849.16,78.88
X$24158 48 700 833 792 795 29 430 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $24793 r0 *1 683.56,78.88
X$24793 48 815 690 767 873 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $24794 r0 *1 685.86,78.88
X$24794 48 815 744 767 29 48 816 29 sky130_fd_sc_hd__a21oi_1
* cell instance $24795 r0 *1 687.7,78.88
X$24795 48 789 786 854 817 29 48 818 29 sky130_fd_sc_hd__a31oi_1
* cell instance $24796 r0 *1 690,78.88
X$24796 48 683 818 834 693 815 48 853 29 29 sky130_fd_sc_hd__o2111ai_1
* cell instance $24800 r0 *1 693.22,78.88
X$24800 48 793 796 797 48 908 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $24801 r0 *1 695.06,78.88
X$24801 48 787 690 858 767 857 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $24803 r0 *1 698.74,78.88
X$24803 29 788 840 819 823 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $24804 r0 *1 702.42,78.88
X$24804 48 819 823 821 859 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $24807 r0 *1 705.64,78.88
X$24807 29 915 822 786 820 821 789 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $24808 r0 *1 708.86,78.88
X$24808 29 1037 803 859 822 48 48 29 sky130_fd_sc_hd__nor3b_2
* cell instance $24809 r0 *1 713.46,78.88
X$24809 48 860 823 637 29 757 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $24811 r0 *1 717.14,78.88
X$24811 48 856 809 972 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $24812 r0 *1 719.44,78.88
X$24812 48 861 755 862 48 29 823 29 sky130_fd_sc_hd__or3_2
* cell instance $24816 r0 *1 722.2,78.88
X$24816 29 687 787 639 856 883 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $24818 r0 *1 730.48,78.88
X$24818 29 29 824 48 710 695 48 sky130_fd_sc_hd__nor2_2
* cell instance $24821 r0 *1 733.7,78.88
X$24821 29 708 898 754 824 780 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $24823 r0 *1 741.98,78.88
X$24823 29 756 551 854 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $24827 r0 *1 752.1,78.88
X$24827 29 551 901 728 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $24829 r0 *1 758.54,78.88
X$24829 48 864 29 487 48 29 sky130_fd_sc_hd__buf_2
* cell instance $24831 r0 *1 760.84,78.88
X$24831 29 783 698 864 813 729 48 48 29 sky130_fd_sc_hd__and4b_1
* cell instance $24833 r0 *1 764.98,78.88
X$24833 29 782 830 866 648 828 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $24835 r0 *1 773.26,78.88
X$24835 48 828 827 892 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $24839 r0 *1 775.56,78.88
X$24839 48 782 829 730 29 48 828 29 sky130_fd_sc_hd__a21o_1
* cell instance $24840 r0 *1 778.32,78.88
X$24840 48 830 829 891 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $24842 r0 *1 780.62,78.88
X$24842 29 847 830 829 782 652 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $24846 r0 *1 788.9,78.88
X$24846 29 845 887 843 746 889 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $24847 r0 *1 796.26,78.88
X$24847 48 887 48 29 888 29 sky130_fd_sc_hd__inv_1
* cell instance $24854 r0 *1 805.92,78.88
X$24854 48 842 48 29 885 29 sky130_fd_sc_hd__inv_1
* cell instance $24855 r0 *1 807.3,78.88
X$24855 48 178 574 882 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $24856 r0 *1 809.6,78.88
X$24856 48 206 608 881 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $24861 r0 *1 816.96,78.88
X$24861 29 878 917 833 877 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $24862 r0 *1 821.56,78.88
X$24862 48 766 608 875 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $24865 r0 *1 827.08,78.88
X$24865 48 644 48 29 869 29 sky130_fd_sc_hd__inv_1
* cell instance $24870 r0 *1 828.92,78.88
X$24870 48 870 869 831 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $24871 r0 *1 832.14,78.88
X$24871 48 542 831 838 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $24872 r0 *1 833.52,78.88
X$24872 48 869 711 870 48 29 504 29 sky130_fd_sc_hd__or3_2
* cell instance $24873 r0 *1 836.28,78.88
X$24873 29 874 633 644 832 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $24877 r0 *1 841.8,78.88
X$24877 48 542 871 835 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $24879 r0 *1 843.64,78.88
X$24879 29 47 795 46 910 48 48 29 sky130_fd_sc_hd__dfrtp_2
* cell instance $25533 m0 *1 684.48,84.32
X$25533 48 815 767 690 48 893 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $25534 m0 *1 686.32,84.32
X$25534 48 894 840 834 906 48 29 29 sky130_fd_sc_hd__or3b_1
* cell instance $25535 m0 *1 689.54,84.32
X$25535 48 856 702 836 894 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $25537 m0 *1 691.84,84.32
X$25537 48 856 702 855 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $25538 m0 *1 693.22,84.32
X$25538 48 815 908 857 29 48 895 29 sky130_fd_sc_hd__a21oi_1
* cell instance $25539 m0 *1 695.06,84.32
X$25539 29 683 789 786 788 48 909 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $25540 m0 *1 699.66,84.32
X$25540 48 840 800 858 48 912 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $25541 m0 *1 701.5,84.32
X$25541 29 29 836 48 819 823 48 sky130_fd_sc_hd__nor2_2
* cell instance $25543 m0 *1 704.26,84.32
X$25543 48 820 688 858 48 29 914 29 sky130_fd_sc_hd__o21ai_1
* cell instance $25545 m0 *1 706.56,84.32
X$25545 48 702 639 758 820 48 876 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $25546 m0 *1 708.86,84.32
X$25546 48 915 815 775 29 48 897 29 sky130_fd_sc_hd__a21oi_1
* cell instance $25549 m0 *1 713.46,84.32
X$25549 29 759 879 861 963 807 883 48 48 29 sky130_fd_sc_hd__o2111ai_2
* cell instance $25551 m0 *1 719.44,84.32
X$25551 29 755 760 861 862 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $25552 m0 *1 723.12,84.32
X$25552 48 755 788 687 810 29 48 921 29 sky130_fd_sc_hd__or4_2
* cell instance $25553 m0 *1 726.34,84.32
X$25553 48 763 685 851 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $25555 m0 *1 729.1,84.32
X$25555 48 447 493 695 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $25556 m0 *1 731.4,84.32
X$25556 48 754 824 705 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $25558 m0 *1 734.16,84.32
X$25558 29 645 863 937 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $25559 m0 *1 744.28,84.32
X$25559 29 447 900 487 785 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $25561 m0 *1 747.04,84.32
X$25561 29 863 645 890 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $25562 m0 *1 757.16,84.32
X$25562 29 900 927 569 852 865 939 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $25563 m0 *1 766.82,84.32
X$25563 48 729 813 783 785 48 825 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $25565 m0 *1 769.58,84.32
X$25565 48 828 827 943 929 29 48 29 sky130_fd_sc_hd__nor3b_1
* cell instance $25566 m0 *1 772.34,84.32
X$25566 48 902 828 926 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $25569 m0 *1 774.64,84.32
X$25569 48 830 926 925 29 48 867 29 sky130_fd_sc_hd__a21oi_1
* cell instance $25570 m0 *1 776.48,84.32
X$25570 29 827 891 868 846 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $25571 m0 *1 782.46,84.32
X$25571 29 29 868 48 866 829 48 sky130_fd_sc_hd__nor2_2
* cell instance $25573 m0 *1 785.22,84.32
X$25573 48 924 48 29 830 29 sky130_fd_sc_hd__buf_4
* cell instance $25575 m0 *1 788.44,84.32
X$25575 48 923 48 29 920 29 sky130_fd_sc_hd__inv_1
* cell instance $25577 m0 *1 790.28,84.32
X$25577 48 143 462 976 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $25579 m0 *1 792.58,84.32
X$25579 29 889 974 885 971 886 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $25583 m0 *1 803.16,84.32
X$25583 48 37 574 965 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $25585 m0 *1 806.38,84.32
X$25585 29 884 958 881 882 880 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $25588 m0 *1 815.12,84.32
X$25588 48 919 576 877 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $25590 m0 *1 818.8,84.32
X$25590 48 917 878 918 29 48 774 29 sky130_fd_sc_hd__a21oi_1
* cell instance $25593 m0 *1 822.02,84.32
X$25593 48 916 841 904 29 48 918 29 sky130_fd_sc_hd__a21o_1
* cell instance $25594 m0 *1 824.78,84.32
X$25594 29 916 904 795 875 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $25597 m0 *1 830.3,84.32
X$25597 48 700 706 832 870 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $25598 m0 *1 832.14,84.32
X$25598 29 2467 874 706 700 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $25600 m0 *1 837.66,84.32
X$25600 48 874 795 952 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $25601 m0 *1 840.88,84.32
X$25601 48 792 48 29 913 29 sky130_fd_sc_hd__inv_1
* cell instance $25603 m0 *1 842.72,84.32
X$25603 48 542 911 872 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $25604 m0 *1 844.1,84.32
X$25604 29 47 833 46 872 48 48 29 sky130_fd_sc_hd__dfrtp_1
* cell instance $26240 r0 *1 684.94,84.32
X$26240 48 893 873 951 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $26241 r0 *1 686.32,84.32
X$26241 48 906 29 931 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $26242 r0 *1 689.08,84.32
X$26242 48 893 853 837 1007 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $26243 r0 *1 690.92,84.32
X$26243 29 894 840 907 834 48 48 29 sky130_fd_sc_hd__nor3b_4
* cell instance $26247 r0 *1 697.82,84.32
X$26247 29 912 954 787 896 836 702 48 48 29 sky130_fd_sc_hd__o32ai_1
* cell instance $26248 r0 *1 701.04,84.32
X$26248 29 930 896 955 914 897 788 48 48 29 sky130_fd_sc_hd__o221a_1
* cell instance $26250 r0 *1 705.64,84.32
X$26250 29 29 744 896 787 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $26253 r0 *1 709.32,84.32
X$26253 48 776 29 759 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $26254 r0 *1 712.08,84.32
X$26254 29 788 962 898 750 961 966 48 48 29 sky130_fd_sc_hd__a2111oi_0
* cell instance $26255 r0 *1 715.3,84.32
X$26255 29 898 970 819 936 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $26256 r0 *1 718.98,84.32
X$26256 48 972 29 786 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $26260 r0 *1 721.74,84.32
X$26260 48 850 876 935 896 815 48 977 29 29 sky130_fd_sc_hd__a311oi_1
* cell instance $26261 r0 *1 724.96,84.32
X$26261 48 978 48 29 922 29 sky130_fd_sc_hd__buf_4
* cell instance $26263 r0 *1 728.18,84.32
X$26263 29 978 860 936 985 779 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $26267 r0 *1 733.24,84.32
X$26267 29 577 979 938 899 602 546 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $26268 r0 *1 743.36,84.32
X$26268 48 865 939 1086 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $26269 r0 *1 745.66,84.32
X$26269 29 712 863 487 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $26274 r0 *1 750.26,84.32
X$26274 29 698 901 980 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $26277 r0 *1 761.3,84.32
X$26277 48 783 785 729 29 48 928 29 sky130_fd_sc_hd__a21o_1
* cell instance $26278 r0 *1 764.06,84.32
X$26278 29 939 652 944 867 848 48 48 29 sky130_fd_sc_hd__nor4b_2
* cell instance $26279 r0 *1 769.58,84.32
X$26279 48 942 929 827 828 48 946 29 29 sky130_fd_sc_hd__a22oi_1
* cell instance $26280 r0 *1 772.34,84.32
X$26280 48 782 946 903 48 29 944 29 sky130_fd_sc_hd__a21boi_1
* cell instance $26284 r0 *1 775.1,84.32
X$26284 48 942 929 830 48 903 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $26285 r0 *1 776.94,84.32
X$26285 48 782 902 1045 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $26286 r0 *1 778.32,84.32
X$26286 29 847 532 846 868 48 48 29 sky130_fd_sc_hd__a21bo_1
* cell instance $26288 r0 *1 782.46,84.32
X$26288 29 924 829 920 888 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $26290 r0 *1 788.44,84.32
X$26290 29 923 973 974 976 975 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $26297 r0 *1 804.54,84.32
X$26297 29 969 1018 965 968 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $26298 r0 *1 809.14,84.32
X$26298 48 958 48 29 964 29 sky130_fd_sc_hd__inv_1
* cell instance $26303 r0 *1 816.04,84.32
X$26303 48 608 440 462 919 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $26304 r0 *1 817.88,84.32
X$26304 29 957 987 455 941 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $26305 r0 *1 822.48,84.32
X$26305 29 948 992 483 688 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $26313 r0 *1 838.58,84.32
X$26313 48 833 795 874 953 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $26314 r0 *1 840.42,84.32
X$26314 48 542 952 910 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $26318 r0 *1 843.64,84.32
X$26318 48 950 905 911 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $26319 r0 *1 846.86,84.32
X$26319 48 795 700 706 950 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $26321 r0 *1 849.16,84.32
X$26321 48 833 48 29 905 29 sky130_fd_sc_hd__inv_1
* cell instance $27250 m0 *1 684.02,89.76
X$27250 29 990 932 981 930 1128 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $27252 r0 *1 684.94,89.76
X$27252 29 1129 1104 1006 690 895 794 48 48 29 sky130_fd_sc_hd__a311oi_2
* cell instance $27253 r0 *1 690.46,89.76
X$27253 48 855 750 990 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $27255 m0 *1 691.84,89.76
X$27255 29 932 931 854 797 758 982 48 48 29 sky130_fd_sc_hd__a2111oi_2
* cell instance $27259 r0 *1 695.98,89.76
X$27259 29 1024 991 909 1010 854 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $27260 m0 *1 697.36,89.76
X$27260 29 788 922 991 750 836 933 48 48 29 sky130_fd_sc_hd__o2111ai_4
* cell instance $27261 r0 *1 699.2,89.76
X$27261 29 1009 702 787 954 914 688 48 48 29 sky130_fd_sc_hd__a32o_1
* cell instance $27263 r0 *1 703.34,89.76
X$27263 48 702 898 750 1028 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $27266 r0 *1 706.56,89.76
X$27266 29 983 1012 1011 1008 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $27268 m0 *1 707.94,89.76
X$27268 29 933 922 758 858 48 959 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $27270 r0 *1 714.38,89.76
X$27270 29 984 970 1030 1011 983 48 48 29 sky130_fd_sc_hd__a2bb2oi_4
* cell instance $27271 m0 *1 715.76,89.76
X$27271 48 890 1013 934 963 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $27275 m0 *1 719.44,89.76
X$27275 48 861 862 999 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $27277 m0 *1 720.82,89.76
X$27277 29 809 933 856 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $27278 r0 *1 724.04,89.76
X$27278 29 984 921 809 856 1174 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $27279 m0 *1 724.96,89.76
X$27279 29 779 789 860 936 985 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $27280 r0 *1 728.64,89.76
X$27280 48 935 688 787 775 29 1035 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $27283 m0 *1 732.78,89.76
X$27283 29 862 814 937 980 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $27284 r0 *1 733.24,89.76
X$27284 29 936 862 1003 48 48 29 sky130_fd_sc_hd__nand2b_2
* cell instance $27285 m0 *1 736.46,89.76
X$27285 29 979 814 934 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $27288 r0 *1 738.76,89.76
X$27288 29 1004 940 861 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $27290 m0 *1 747.04,89.76
X$27290 29 940 1004 1003 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $27294 r0 *1 750.26,89.76
X$27294 29 901 698 1013 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $27296 m0 *1 753.48,89.76
X$27296 29 729 1005 940 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $27298 r0 *1 760.84,89.76
X$27298 29 782 827 1036 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $27299 m0 *1 763.6,89.76
X$27299 29 783 813 901 729 48 48 29 sky130_fd_sc_hd__nand3b_4
* cell instance $27300 m0 *1 770.96,89.76
X$27300 48 790 652 945 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $27301 r0 *1 770.96,89.76
X$27301 48 830 942 1014 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $27302 r0 *1 772.34,89.76
X$27302 29 865 652 826 849 867 944 48 48 29 sky130_fd_sc_hd__o41a_1
* cell instance $27305 m0 *1 774.64,89.76
X$27305 48 782 892 947 29 48 849 29 sky130_fd_sc_hd__a21oi_1
* cell instance $27306 r0 *1 776.48,89.76
X$27306 29 902 866 1015 1002 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $27307 m0 *1 776.48,89.76
X$27307 48 943 827 790 986 48 947 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $27310 m0 *1 781.08,89.76
X$27310 29 1015 1002 782 830 48 646 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $27312 r0 *1 784.3,89.76
X$27312 48 866 1002 1047 29 48 1016 29 sky130_fd_sc_hd__a21oi_1
* cell instance $27314 r0 *1 786.6,89.76
X$27314 48 1017 1016 942 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $27320 m0 *1 792.58,89.76
X$27320 48 973 48 29 1001 29 sky130_fd_sc_hd__inv_1
* cell instance $27323 m0 *1 794.42,89.76
X$27323 29 971 967 998 844 1000 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $27324 r0 *1 794.88,89.76
X$27324 48 37 368 998 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $27325 r0 *1 797.18,89.76
X$27325 29 975 1034 997 1033 1124 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $27328 m0 *1 802.24,89.76
X$27328 29 886 997 964 967 1019 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $27329 r0 *1 804.54,89.76
X$27329 48 1018 48 29 1033 29 sky130_fd_sc_hd__inv_1
* cell instance $27330 r0 *1 805.92,89.76
X$27330 48 68 440 1071 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $27331 r0 *1 807.3,89.76
X$27331 48 33 462 1069 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $27336 m0 *1 811.9,89.76
X$27336 29 996 995 435 960 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $27343 r0 *1 816.96,89.76
X$27343 48 995 957 987 29 48 1032 29 sky130_fd_sc_hd__a21o_1
* cell instance $27344 m0 *1 818.34,89.76
X$27344 48 957 948 994 996 48 956 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $27347 r0 *1 820.64,89.76
X$27347 29 1049 1029 541 1031 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $27349 m0 *1 822.02,89.76
X$27349 48 992 948 993 29 48 988 29 sky130_fd_sc_hd__a21oi_1
* cell instance $27351 r0 *1 825.24,89.76
X$27351 48 956 1020 1021 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $27355 r0 *1 828,89.76
X$27355 29 745 1062 1021 989 1060 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $27363 m0 *1 838.12,89.76
X$27363 48 953 913 871 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $27366 m0 *1 841.34,89.76
X$27366 48 913 905 949 832 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $27367 r0 *1 841.34,89.76
X$27367 48 1058 1022 989 48 1027 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $27368 m0 *1 843.18,89.76
X$27368 48 795 48 29 949 29 sky130_fd_sc_hd__inv_1
* cell instance $27371 r0 *1 844.1,89.76
X$27371 29 989 1025 905 1026 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $27374 r0 *1 848.7,89.76
X$27374 29 1156 1055 706 1023 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $28330 m0 *1 691.84,95.2
X$28330 48 1024 48 29 981 29 sky130_fd_sc_hd__buf_4
* cell instance $28333 m0 *1 694.6,95.2
X$28333 29 991 909 1010 1076 854 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $28334 m0 *1 702.42,95.2
X$28334 29 982 744 1037 688 1038 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $28335 m0 *1 705.64,95.2
X$28335 29 933 1038 922 775 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $28337 m0 *1 709.78,95.2
X$28337 29 1039 1028 962 815 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $28338 m0 *1 713.92,95.2
X$28338 48 898 819 936 961 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $28339 m0 *1 715.76,95.2
X$28339 48 819 1003 963 1077 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $28343 m0 *1 719.44,95.2
X$28343 48 759 999 966 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $28346 m0 *1 720.82,95.2
X$28346 29 809 1078 856 999 1107 921 48 48 29 sky130_fd_sc_hd__o2111ai_2
* cell instance $28348 m0 *1 728.18,95.2
X$28348 48 935 1136 787 981 29 1040 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $28349 m0 *1 730.48,95.2
X$28349 48 1041 1035 1040 977 29 48 1080 29 sky130_fd_sc_hd__or4_2
* cell instance $28352 m0 *1 737.84,95.2
X$28352 48 940 980 938 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $28353 m0 *1 739.22,95.2
X$28353 29 546 602 1004 899 577 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $28355 m0 *1 747.04,95.2
X$28355 29 546 602 1079 1043 577 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $28358 m0 *1 754.4,95.2
X$28358 29 29 927 48 1042 1043 48 sky130_fd_sc_hd__nor2_2
* cell instance $28359 m0 *1 756.7,95.2
X$28359 29 927 852 900 939 865 598 48 48 29 sky130_fd_sc_hd__o221a_2
* cell instance $28360 m0 *1 760.84,95.2
X$28360 29 902 830 1044 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $28361 m0 *1 770.96,95.2
X$28361 48 943 945 1036 1044 29 48 785 29 sky130_fd_sc_hd__and4_1
* cell instance $28365 m0 *1 774.64,95.2
X$28365 48 943 827 790 1045 48 925 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $28366 m0 *1 776.94,95.2
X$28366 29 1002 1046 866 1001 48 48 29 sky130_fd_sc_hd__ha_4
* cell instance $28367 m0 *1 786.14,95.2
X$28367 29 1017 986 830 1016 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $28368 m0 *1 788.44,95.2
X$28368 29 1074 1047 1075 1073 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $28369 m0 *1 793.04,95.2
X$28369 29 1075 1046 1125 1122 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $28375 m0 *1 802.24,95.2
X$28375 48 969 48 29 1072 29 sky130_fd_sc_hd__inv_1
* cell instance $28376 m0 *1 803.62,95.2
X$28376 29 1127 1070 1069 1068 1071 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $28377 m0 *1 810.98,95.2
X$28377 48 102 608 1068 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $28378 m0 *1 812.36,95.2
X$28378 29 994 1048 555 1067 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $28380 m0 *1 817.42,95.2
X$28380 48 994 1032 1048 29 48 993 29 sky130_fd_sc_hd__a21o_1
* cell instance $28382 m0 *1 821.1,95.2
X$28382 48 1049 1050 1064 1161 48 1020 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $28383 m0 *1 823.4,95.2
X$28383 48 1120 1050 1203 29 48 1065 29 sky130_fd_sc_hd__a21oi_1
* cell instance $28384 m0 *1 825.24,95.2
X$28384 48 1066 1049 1029 29 48 1063 29 sky130_fd_sc_hd__a21o_1
* cell instance $28385 m0 *1 828,95.2
X$28385 48 1061 1052 1062 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $28389 m0 *1 829.84,95.2
X$28389 48 1051 1021 1200 29 48 1060 29 sky130_fd_sc_hd__a21oi_1
* cell instance $28390 m0 *1 831.68,95.2
X$28390 48 1053 1097 1157 29 48 1202 29 sky130_fd_sc_hd__a21oi_1
* cell instance $28394 m0 *1 841.8,95.2
X$28394 48 1027 1025 1059 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $28395 m0 *1 844.1,95.2
X$28395 29 1100 1058 949 1056 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $28397 m0 *1 849.62,95.2
X$28397 48 1055 1057 1054 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $29049 r0 *1 684.94,95.2
X$29049 48 1008 1081 1105 48 1104 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $29050 r0 *1 686.78,95.2
X$29050 48 854 48 29 1105 29 sky130_fd_sc_hd__buf_4
* cell instance $29053 r0 *1 691.84,95.2
X$29053 48 1008 1081 1166 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $29057 r0 *1 695.52,95.2
X$29057 29 909 1082 1010 991 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $29059 r0 *1 698.28,95.2
X$29059 29 1006 1082 854 1083 1135 1039 48 48 29 sky130_fd_sc_hd__a41oi_2
* cell instance $29062 r0 *1 705.64,95.2
X$29062 48 1038 1136 1037 48 29 1106 29 sky130_fd_sc_hd__a21o_2
* cell instance $29063 r0 *1 708.86,95.2
X$29063 29 1083 1078 879 1077 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $29064 r0 *1 712.54,95.2
X$29064 29 879 1081 1078 1077 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $29066 r0 *1 715.3,95.2
X$29066 48 970 984 1012 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $29067 r0 *1 716.68,95.2
X$29067 29 809 856 983 819 936 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $29069 r0 *1 724.04,95.2
X$29069 48 1085 1108 1084 776 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $29070 r0 *1 725.88,95.2
X$29070 48 985 1108 1085 1084 29 1107 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $29072 r0 *1 729.1,95.2
X$29072 29 921 1443 966 1110 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $29074 r0 *1 733.24,95.2
X$29074 29 1086 1079 1113 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $29075 r0 *1 743.36,95.2
X$29075 48 1079 1086 1084 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $29079 r0 *1 751.18,95.2
X$29079 48 544 548 1087 636 1114 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $29081 r0 *1 755.78,95.2
X$29081 29 1117 1088 495 496 412 1089 48 48 29 sky130_fd_sc_hd__o41a_2
* cell instance $29083 r0 *1 760.84,95.2
X$29083 29 783 813 1042 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $29084 r0 *1 770.96,95.2
X$29084 48 790 1014 943 29 48 826 29 sky130_fd_sc_hd__a21oi_1
* cell instance $29085 r0 *1 772.8,95.2
X$29085 29 1002 1093 1092 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $29087 r0 *1 782.92,95.2
X$29087 29 846 1093 1002 48 48 29 sky130_fd_sc_hd__nand2b_2
* cell instance $29088 r0 *1 786.14,95.2
X$29088 48 1002 1095 1074 1017 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $29090 r0 *1 788.44,95.2
X$29090 48 102 462 1211 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $29091 r0 *1 790.74,95.2
X$29091 29 1170 1122 1123 1121 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29093 r0 *1 795.8,95.2
X$29093 48 1034 48 29 1125 29 sky130_fd_sc_hd__inv_1
* cell instance $29095 r0 *1 798.1,95.2
X$29095 29 1124 1126 1096 1072 1127 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $29098 r0 *1 806.38,95.2
X$29098 48 1126 48 29 1123 29 sky130_fd_sc_hd__inv_1
* cell instance $29103 r0 *1 813.28,95.2
X$29103 48 32 29 462 48 29 sky130_fd_sc_hd__buf_2
* cell instance $29108 r0 *1 820.64,95.2
X$29108 29 1050 1120 422 1090 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29109 r0 *1 825.24,95.2
X$29109 48 956 1065 988 48 1051 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $29110 r0 *1 827.08,95.2
X$29110 29 1097 1053 732 1119 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29112 r0 *1 831.68,95.2
X$29112 29 1116 1115 711 1118 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29113 r0 *1 836.28,95.2
X$29113 29 1098 1099 913 1240 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29114 r0 *1 840.88,95.2
X$29114 48 1099 1098 1059 29 48 1199 29 sky130_fd_sc_hd__a21oi_1
* cell instance $29117 r0 *1 843.64,95.2
X$29117 48 1100 1054 1101 48 1022 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $29119 r0 *1 847.32,95.2
X$29119 29 1057 1101 734 1112 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29121 r0 *1 852.38,95.2
X$29121 29 1103 1237 1109 1102 1111 1154 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $29760 m0 *1 684.94,100.64
X$29760 48 1128 1129 1130 951 48 29 1163 29 sky130_fd_sc_hd__o211a_2
* cell instance $29761 m0 *1 688.62,100.64
X$29761 48 1129 1130 951 48 1162 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $29763 m0 *1 691.84,100.64
X$29763 48 1166 1131 1006 1165 1130 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $29766 m0 *1 695.06,100.64
X$29766 48 1133 1132 1105 29 1131 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $29769 m0 *1 702.88,100.64
X$29769 48 1134 1181 1135 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $29770 m0 *1 704.26,100.64
X$29770 29 1133 1038 1037 1136 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $29773 m0 *1 711.62,100.64
X$29773 29 959 1132 896 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $29775 m0 *1 716.68,100.64
X$29775 48 861 1013 934 1137 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $29777 m0 *1 719.44,100.64
X$29777 48 1137 48 29 1169 29 sky130_fd_sc_hd__inv_1
* cell instance $29780 m0 *1 720.82,100.64
X$29780 48 860 48 29 819 29 sky130_fd_sc_hd__buf_4
* cell instance $29781 m0 *1 723.58,100.64
X$29781 48 1085 1084 1171 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $29782 m0 *1 724.96,100.64
X$29782 48 786 1138 789 1311 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $29783 m0 *1 726.8,100.64
X$29783 48 1138 1113 985 1174 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $29785 m0 *1 729.1,100.64
X$29785 48 1138 1113 1207 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $29787 m0 *1 732.32,100.64
X$29787 48 640 1085 1084 1139 1110 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $29789 m0 *1 736,100.64
X$29789 48 1136 48 29 688 29 sky130_fd_sc_hd__buf_4
* cell instance $29791 m0 *1 740.6,100.64
X$29791 29 548 636 544 762 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $29793 m0 *1 747.04,100.64
X$29793 29 29 927 899 1086 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $29796 m0 *1 749.34,100.64
X$29796 29 544 548 636 1140 48 1141 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $29797 m0 *1 757.16,100.64
X$29797 29 813 783 1445 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $29798 m0 *1 767.28,100.64
X$29798 48 1178 1092 1251 1087 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $29799 m0 *1 769.12,100.64
X$29799 48 1091 1036 1177 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $29801 m0 *1 772.8,100.64
X$29801 48 1142 1094 1175 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $29805 m0 *1 774.64,100.64
X$29805 48 1176 1143 1091 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $29806 m0 *1 776.02,100.64
X$29806 29 1093 1173 1172 1144 1215 48 48 29 sky130_fd_sc_hd__fa_2
* cell instance $29808 m0 *1 784.76,100.64
X$29808 48 1095 1074 1047 29 48 1015 29 sky130_fd_sc_hd__a21o_1
* cell instance $29809 m0 *1 787.52,100.64
X$29809 29 1212 1073 1170 1309 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29810 m0 *1 792.12,100.64
X$29810 48 1075 48 29 1144 29 sky130_fd_sc_hd__inv_1
* cell instance $29811 m0 *1 793.5,100.64
X$29811 48 101 440 1209 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $29813 m0 *1 796.72,100.64
X$29813 48 1168 48 29 1121 29 sky130_fd_sc_hd__inv_1
* cell instance $29815 m0 *1 798.56,100.64
X$29815 48 101 576 1206 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $29817 m0 *1 800.4,100.64
X$29817 48 1145 48 29 1167 29 sky130_fd_sc_hd__inv_1
* cell instance $29829 m0 *1 809.6,100.64
X$29829 48 206 440 1164 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $29835 m0 *1 816.5,100.64
X$29835 29 1064 1204 713 1146 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29838 m0 *1 822.48,100.64
X$29838 29 1161 1066 651 1160 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29840 m0 *1 827.54,100.64
X$29840 48 1097 1116 1159 1061 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $29844 m0 *1 829.84,100.64
X$29844 29 1159 1147 869 1158 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $29845 m0 *1 834.44,100.64
X$29845 48 1116 1147 1115 29 48 1157 29 sky130_fd_sc_hd__a21o_1
* cell instance $29849 m0 *1 843.18,100.64
X$29849 48 1057 1156 1100 1098 48 1052 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $29852 m0 *1 850.08,100.64
X$29852 48 1190 1026 1155 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $29853 m0 *1 851.46,100.64
X$29853 48 1148 48 29 1112 29 sky130_fd_sc_hd__inv_1
* cell instance $29854 m0 *1 852.84,100.64
X$29854 29 1154 1155 1026 1056 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $29858 m0 *1 857.44,100.64
X$29858 29 1153 1197 1196 1056 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $29859 m0 *1 861.12,100.64
X$29859 48 1152 1109 1148 1150 29 48 29 sky130_fd_sc_hd__nand3b_1
* cell instance $29860 m0 *1 863.88,100.64
X$29860 48 1056 1149 1151 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30793 m0 *1 678.96,106.08
X$30793 48 1179 907 1253 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30795 m0 *1 682.18,106.08
X$30795 48 1030 726 1217 48 1179 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $30796 m0 *1 685.4,106.08
X$30796 29 1253 769 1281 1192 1218 1235 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $30799 r0 *1 686.78,100.64
X$30799 48 1132 931 1235 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30800 r0 *1 688.16,100.64
X$30800 29 1192 769 1193 1007 1009 1179 48 48 29 sky130_fd_sc_hd__o2111a_1
* cell instance $30802 m0 *1 689.54,106.08
X$30802 48 1105 931 1180 1193 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $30804 m0 *1 691.84,106.08
X$30804 48 1030 1217 1254 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30805 r0 *1 692.3,100.64
X$30805 29 1239 1180 907 1105 1132 1133 48 48 29 sky130_fd_sc_hd__o2111a_1
* cell instance $30809 m0 *1 693.22,106.08
X$30809 29 726 1272 1106 1198 907 1219 48 48 29 sky130_fd_sc_hd__a2111oi_0
* cell instance $30810 r0 *1 696.44,100.64
X$30810 48 1219 769 1007 48 29 1195 29 sky130_fd_sc_hd__o21ai_1
* cell instance $30811 m0 *1 696.44,106.08
X$30811 48 1083 1241 1134 29 48 1217 29 sky130_fd_sc_hd__o21a_2
* cell instance $30812 r0 *1 698.28,100.64
X$30812 48 1134 1241 1030 1083 1180 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $30813 m0 *1 699.66,106.08
X$30813 29 1274 1258 1030 1081 1135 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $30815 r0 *1 701.96,100.64
X$30815 48 1134 1181 1030 1083 1198 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $30816 m0 *1 704.26,106.08
X$30816 48 933 819 922 1241 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $30819 r0 *1 705.64,100.64
X$30819 48 933 1182 922 1181 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $30821 m0 *1 706.56,106.08
X$30821 48 1134 1241 1244 1169 1221 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $30822 r0 *1 707.48,100.64
X$30822 48 933 922 759 29 1244 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $30823 m0 *1 709.32,106.08
X$30823 48 1255 1221 1223 1222 1219 1220 48 29 29 sky130_fd_sc_hd__o221ai_1
* cell instance $30825 r0 *1 711.62,100.64
X$30825 29 1134 1183 789 786 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $30826 m0 *1 712.54,106.08
X$30826 29 688 1201 819 1222 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $30827 r0 *1 717.6,100.64
X$30827 48 786 789 1183 29 48 1201 29 sky130_fd_sc_hd__a21o_1
* cell instance $30830 m0 *1 719.44,106.08
X$30830 48 819 934 1201 1255 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $30835 r0 *1 720.82,100.64
X$30835 48 896 959 1246 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30836 m0 *1 721.28,106.08
X$30836 48 1246 29 1219 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $30838 r0 *1 724.04,100.64
X$30838 48 1184 1171 1182 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30839 m0 *1 724.04,106.08
X$30839 48 1256 1207 1171 1108 29 48 1183 29 sky130_fd_sc_hd__or4_2
* cell instance $30841 r0 *1 726.34,100.64
X$30841 29 1113 1184 1138 48 860 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $30842 m0 *1 727.26,106.08
X$30842 48 762 1257 935 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30843 m0 *1 728.64,106.08
X$30843 48 789 786 1224 1085 29 1278 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $30844 m0 *1 731.4,106.08
X$30844 29 1277 1278 1113 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $30846 r0 *1 733.24,100.64
X$30846 48 696 1185 985 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $30847 r0 *1 735.54,100.64
X$30847 48 1210 1136 48 29 29 sky130_fd_sc_hd__clkinv_2
* cell instance $30850 m0 *1 737.84,106.08
X$30850 29 29 1210 48 933 922 48 sky130_fd_sc_hd__nor2_2
* cell instance $30851 r0 *1 738.3,100.64
X$30851 48 1210 29 815 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $30852 m0 *1 740.14,106.08
X$30852 48 1258 29 1067 48 29 sky130_fd_sc_hd__clkinv_4
* cell instance $30854 r0 *1 741.52,100.64
X$30854 29 1138 1213 1186 1141 48 48 29 sky130_fd_sc_hd__mux2_2
* cell instance $30856 m0 *1 743.82,106.08
X$30856 48 933 922 1276 1287 1226 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $30857 r0 *1 745.66,100.64
X$30857 29 1213 1085 1186 1141 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $30859 m0 *1 747.04,106.08
X$30859 48 1226 1216 1225 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30863 m0 *1 750.26,106.08
X$30863 48 1228 1227 1213 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30864 m0 *1 751.64,106.08
X$30864 48 1178 1259 1227 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30865 m0 *1 753.02,106.08
X$30865 48 1228 1360 1186 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30866 r0 *1 753.94,100.64
X$30866 48 1114 1228 48 1216 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $30867 m0 *1 754.4,106.08
X$30867 48 1187 1273 1259 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30870 r0 *1 757.62,100.64
X$30870 48 1187 1088 1252 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30871 m0 *1 758.08,106.08
X$30871 48 1142 1178 1288 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30872 r0 *1 759,100.64
X$30872 48 783 785 1005 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30873 m0 *1 759.46,106.08
X$30873 48 1142 1178 1088 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30876 r0 *1 761.3,100.64
X$30876 29 1043 1044 1087 1177 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $30877 m0 *1 761.76,106.08
X$30877 48 1273 1187 1140 1251 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $30878 m0 *1 763.6,106.08
X$30878 29 1044 943 1228 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $30880 r0 *1 765.44,100.64
X$30880 29 1188 1044 945 1036 48 813 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $30881 m0 *1 769.58,106.08
X$30881 48 1172 29 1273 48 29 sky130_fd_sc_hd__buf_2
* cell instance $30882 m0 *1 771.42,106.08
X$30882 48 1260 48 29 1187 29 sky130_fd_sc_hd__buf_4
* cell instance $30883 r0 *1 773.26,100.64
X$30883 29 1188 1092 1143 1176 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $30888 m0 *1 774.64,106.08
X$30888 29 943 1092 1175 1143 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $30889 r0 *1 779.24,100.64
X$30889 48 1095 48 29 1173 29 sky130_fd_sc_hd__inv_1
* cell instance $30890 m0 *1 780.62,106.08
X$30890 29 1229 1089 1271 1214 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $30892 r0 *1 781.54,100.64
X$30892 48 1073 48 29 1215 29 sky130_fd_sc_hd__inv_1
* cell instance $30894 r0 *1 783.38,100.64
X$30894 29 1260 1095 1212 1250 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $30900 m0 *1 788.44,106.08
X$30900 48 37 608 1249 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30901 r0 *1 790.28,100.64
X$30901 29 1214 1247 1211 1209 48 48 29 sky130_fd_sc_hd__ha_2
* cell instance $30903 m0 *1 791.2,106.08
X$30903 29 1270 1269 1249 1248 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $30904 r0 *1 795.8,100.64
X$30904 48 1189 48 29 1208 29 sky130_fd_sc_hd__inv_1
* cell instance $30905 r0 *1 797.18,100.64
X$30905 29 1168 1189 1070 1206 1167 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $30906 m0 *1 798.1,106.08
X$30906 48 178 440 1308 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30914 m0 *1 803.16,106.08
X$30914 29 32 37 1230 1245 1229 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $30917 r0 *1 805.92,100.64
X$30917 48 178 576 1205 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30918 r0 *1 808.22,100.64
X$30918 29 1019 1096 1164 1205 1243 48 48 29 sky130_fd_sc_hd__fa_1
* cell instance $30926 r0 *1 822.02,100.64
X$30926 48 1064 1063 1204 29 48 1203 29 sky130_fd_sc_hd__a21o_1
* cell instance $30928 m0 *1 824.32,106.08
X$30928 48 1158 1231 1242 48 29 1268 29 sky130_fd_sc_hd__o21ai_1
* cell instance $30931 m0 *1 826.62,106.08
X$30931 48 1190 1158 1242 1231 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $30940 r0 *1 829.84,100.64
X$30940 48 1061 1199 1202 48 1200 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $30943 m0 *1 833.98,106.08
X$30943 48 1262 1303 1304 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30945 m0 *1 835.36,106.08
X$30945 48 1267 29 1240 48 29 sky130_fd_sc_hd__buf_2
* cell instance $30946 m0 *1 837.2,106.08
X$30946 29 1420 1111 1295 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $30948 m0 *1 841.34,106.08
X$30948 48 1383 29 48 1267 29 sky130_fd_sc_hd__inv_2
* cell instance $30952 m0 *1 843.18,106.08
X$30952 29 1237 1026 1232 1262 1238 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $30955 r0 *1 845.02,100.64
X$30955 48 1111 48 29 1238 29 sky130_fd_sc_hd__inv_1
* cell instance $30959 m0 *1 849.16,106.08
X$30959 48 1194 1026 1296 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $30962 m0 *1 852.38,106.08
X$30962 48 1232 1111 1103 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30964 m0 *1 853.76,106.08
X$30964 48 1191 1263 1102 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30966 r0 *1 855.14,100.64
X$30966 48 1026 1111 1197 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $30970 r0 *1 856.52,100.64
X$30970 48 1111 1026 1196 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30973 m0 *1 859.28,106.08
X$30973 29 1266 1337 1236 1150 1229 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $30974 r0 *1 859.74,100.64
X$30974 48 1148 1109 1152 1190 48 1236 29 29 sky130_fd_sc_hd__nand4b_1
* cell instance $30975 m0 *1 862.5,106.08
X$30975 48 1151 1194 1301 1191 1335 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $30976 r0 *1 862.96,100.64
X$30976 48 1191 1194 1152 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $30977 m0 *1 864.8,106.08
X$30977 48 1264 1149 1109 1233 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $30978 r0 *1 866.18,100.64
X$30978 48 1264 1109 1234 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $30980 m0 *1 867.56,106.08
X$30980 29 1265 1233 1299 1148 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $30981 r0 *1 868.48,100.64
X$30981 48 1191 29 48 1056 29 sky130_fd_sc_hd__inv_2
* cell instance $32010 r0 *1 681.26,106.08
X$32010 48 907 1198 1389 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32012 r0 *1 683.1,106.08
X$32012 48 1165 907 1030 1331 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $32013 r0 *1 684.94,106.08
X$32013 48 1165 1254 1105 48 1279 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $32014 r0 *1 686.78,106.08
X$32014 48 1067 931 1280 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32015 r0 *1 688.16,106.08
X$32015 29 1391 1280 1331 1128 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $32016 r0 *1 691.84,106.08
X$32016 29 1105 1282 981 931 1132 1133 48 48 29 sky130_fd_sc_hd__a2111oi_0
* cell instance $32020 r0 *1 695.06,106.08
X$32020 48 1282 1239 1272 937 48 29 1340 29 sky130_fd_sc_hd__o31ai_1
* cell instance $32021 r0 *1 697.82,106.08
X$32021 29 1106 1218 1076 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $32023 r0 *1 702.88,106.08
X$32023 48 1134 890 759 934 29 1285 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $32025 r0 *1 705.64,106.08
X$32025 29 1284 1343 1134 934 1283 1285 48 48 29 sky130_fd_sc_hd__a311oi_4
* cell instance $32026 r0 *1 715.3,106.08
X$32026 29 1223 759 688 1169 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $32027 r0 *1 718.98,106.08
X$32027 48 1003 1244 1316 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32032 r0 *1 720.82,106.08
X$32032 48 1003 980 1347 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32033 r0 *1 722.2,106.08
X$32033 48 1311 1286 1224 29 48 1350 29 sky130_fd_sc_hd__a21o_1
* cell instance $32034 r0 *1 724.96,106.08
X$32034 29 1351 1311 896 1224 1286 959 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $32036 r0 *1 728.64,106.08
X$32036 48 786 789 1256 29 48 1286 29 sky130_fd_sc_hd__a21o_1
* cell instance $32041 r0 *1 733.7,106.08
X$32041 29 29 1184 48 1042 1224 48 sky130_fd_sc_hd__nor2_2
* cell instance $32043 r0 *1 737.84,106.08
X$32043 29 1355 640 1210 762 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $32044 r0 *1 743.82,106.08
X$32044 48 688 1276 1357 1287 1411 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $32045 r0 *1 746.58,106.08
X$32045 48 1313 762 1358 29 48 1402 29 sky130_fd_sc_hd__a21oi_1
* cell instance $32050 r0 *1 748.88,106.08
X$32050 29 1276 1257 727 1319 1141 1314 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $32051 r0 *1 752.1,106.08
X$32051 48 1359 1273 48 1319 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $32052 r0 *1 755.32,106.08
X$32052 48 1259 1288 1273 1117 48 1360 29 29 sky130_fd_sc_hd__a22oi_1
* cell instance $32053 r0 *1 758.08,106.08
X$32053 48 1089 1187 1361 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $32055 r0 *1 760.84,106.08
X$32055 29 1288 1257 1117 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $32056 r0 *1 764.98,106.08
X$32056 48 1142 1089 1405 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $32058 r0 *1 767.74,106.08
X$32058 48 1273 1187 29 48 1143 29 sky130_fd_sc_hd__nor2b_2
* cell instance $32059 r0 *1 770.96,106.08
X$32059 29 1187 1176 1194 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $32063 r0 *1 781.08,106.08
X$32063 29 1271 1178 1214 48 1176 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $32066 r0 *1 788.44,106.08
X$32066 48 1289 1312 1307 1310 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $32067 r0 *1 790.28,106.08
X$32067 29 1401 1309 1208 1269 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $32069 r0 *1 795.8,106.08
X$32069 48 1214 48 29 1245 29 sky130_fd_sc_hd__inv_1
* cell instance $32070 r0 *1 797.18,106.08
X$32070 29 1248 1145 1308 1356 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $32080 r0 *1 816.04,106.08
X$32080 48 1291 1306 1290 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32081 r0 *1 817.42,106.08
X$32081 48 1305 1292 1348 48 1349 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $32084 r0 *1 822.02,106.08
X$32084 48 1325 1346 1290 48 29 1294 29 sky130_fd_sc_hd__o21ai_1
* cell instance $32085 r0 *1 823.86,106.08
X$32085 29 1303 1242 1293 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $32090 r0 *1 830.3,106.08
X$32090 48 1190 1242 1345 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32091 r0 *1 831.68,106.08
X$32091 29 1268 1295 1304 1267 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $32092 r0 *1 839.96,106.08
X$32092 29 1327 1341 1267 1302 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $32097 r0 *1 847.78,106.08
X$32097 29 1149 1296 1111 1262 1338 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $32098 r0 *1 852.38,106.08
X$32098 48 1232 1296 1338 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32099 r0 *1 853.76,106.08
X$32099 48 1026 48 29 1263 29 sky130_fd_sc_hd__inv_1
* cell instance $32105 r0 *1 857.9,106.08
X$32105 48 1190 1148 1109 1152 1337 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $32106 r0 *1 860.66,106.08
X$32106 48 1297 1149 1301 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32107 r0 *1 862.04,106.08
X$32107 48 1335 1336 1333 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32108 r0 *1 865.26,106.08
X$32108 48 1384 1300 1264 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32109 r0 *1 866.64,106.08
X$32109 48 1334 1336 1299 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32113 r0 *1 871.7,106.08
X$32113 48 1191 1298 1334 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32114 r0 *1 873.08,106.08
X$32114 29 1329 1265 1330 1429 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $32754 m0 *1 678.96,111.52
X$32754 29 1390 1389 1332 1128 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $32755 m0 *1 682.64,111.52
X$32755 48 1217 1008 1362 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32756 m0 *1 685.86,111.52
X$32756 29 907 1332 1105 1362 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $32757 m0 *1 688.16,111.52
X$32757 48 726 1391 1627 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32760 m0 *1 691.84,111.52
X$32760 48 1008 1315 1363 48 1393 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $32761 m0 *1 695.06,111.52
X$32761 48 1363 1315 1283 1131 1364 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $32762 m0 *1 698.28,111.52
X$32762 48 1076 1106 1219 726 1315 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $32763 m0 *1 701.04,111.52
X$32763 48 1219 1135 815 1182 1342 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $32764 m0 *1 703.34,111.52
X$32764 29 1394 1365 1220 1395 1366 48 48 29 sky130_fd_sc_hd__nor4b_2
* cell instance $32765 m0 *1 708.86,111.52
X$32765 48 1076 1106 1221 1365 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $32766 m0 *1 710.7,111.52
X$32766 48 1133 981 1316 1132 29 1397 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $32768 m0 *1 713.92,111.52
X$32768 29 1343 1284 934 759 1367 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $32769 m0 *1 717.14,111.52
X$32769 48 1368 861 1342 29 48 1549 29 sky130_fd_sc_hd__a21oi_1
* cell instance $32771 m0 *1 719.44,111.52
X$32771 48 1222 1316 1368 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32772 m0 *1 720.82,111.52
X$32772 48 1369 1222 1106 726 29 1275 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $32773 m0 *1 723.58,111.52
X$32773 48 890 934 1369 1367 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $32775 m0 *1 725.88,111.52
X$32775 29 1399 1350 1351 1277 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $32777 m0 *1 731.4,111.52
X$32777 29 1317 1076 1225 1219 1106 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $32778 m0 *1 736,111.52
X$32778 29 1258 1433 1434 1317 48 1318 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $32779 m0 *1 743.82,111.52
X$32779 48 933 922 1402 48 1357 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $32782 m0 *1 747.04,111.52
X$32782 48 762 1140 1403 1257 29 1313 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $32783 m0 *1 749.8,111.52
X$32783 29 1256 762 1216 1436 1370 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $32784 m0 *1 754.4,111.52
X$32784 48 1252 727 1314 29 48 1359 29 sky130_fd_sc_hd__a21oi_1
* cell instance $32785 m0 *1 756.24,111.52
X$32785 48 1361 1273 1320 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32786 m0 *1 759.46,111.52
X$32786 48 1320 1288 1273 1117 29 1370 48 29 sky130_fd_sc_hd__a22o_1
* cell instance $32788 m0 *1 763.14,111.52
X$32788 29 1176 1371 1092 1143 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $32789 m0 *1 765.44,111.52
X$32789 48 1405 48 29 1140 29 sky130_fd_sc_hd__buf_4
* cell instance $32790 m0 *1 768.2,111.52
X$32790 48 1044 1188 48 1372 29 29 sky130_fd_sc_hd__and2_2
* cell instance $32792 m0 *1 771.88,111.52
X$32792 48 1371 1188 1373 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $32794 m0 *1 774.64,111.52
X$32794 29 1176 1187 1377 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $32795 m0 *1 784.76,111.52
X$32795 48 1094 29 1178 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $32797 m0 *1 787.98,111.52
X$32797 29 1094 1250 1401 1437 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $32798 m0 *1 792.58,111.52
X$32798 48 1374 1257 1118 29 48 1322 29 sky130_fd_sc_hd__a21oi_1
* cell instance $32799 m0 *1 794.42,111.52
X$32799 48 1375 1321 1354 1289 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $32800 m0 *1 796.26,111.52
X$32800 48 1376 1322 1353 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32801 m0 *1 797.64,111.52
X$32801 48 1398 1118 1374 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32805 m0 *1 802.24,111.52
X$32805 48 1377 1230 1354 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32806 m0 *1 803.62,111.52
X$32806 48 1262 1232 1323 48 29 1396 29 sky130_fd_sc_hd__o21ai_1
* cell instance $32807 m0 *1 805.46,111.52
X$32807 48 1323 1118 1306 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32809 m0 *1 809.6,111.52
X$32809 48 1378 1379 48 1346 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $32812 m0 *1 814.2,111.52
X$32812 48 1324 1380 1348 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32813 m0 *1 815.58,111.52
X$32813 29 1392 1305 1306 1380 1352 1324 48 48 29 sky130_fd_sc_hd__o41ai_1
* cell instance $32815 m0 *1 819.26,111.52
X$32815 48 1470 1352 1381 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32817 m0 *1 822.94,111.52
X$32817 48 1432 1293 1506 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32818 m0 *1 826.16,111.52
X$32818 48 1242 1325 1344 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $32822 m0 *1 831.22,111.52
X$32822 48 1232 1325 1388 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32824 m0 *1 833.06,111.52
X$32824 48 1324 1303 1302 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $32825 m0 *1 834.44,111.52
X$32825 48 1240 1327 1302 48 1326 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $32826 m0 *1 837.66,111.52
X$32826 48 1305 1573 1382 48 29 1339 29 sky130_fd_sc_hd__o21ai_1
* cell instance $32827 m0 *1 839.5,111.52
X$32827 29 1383 1450 1421 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $32828 m0 *1 849.62,111.52
X$32828 29 1328 1111 1431 1423 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $32829 m0 *1 853.76,111.52
X$32829 48 1190 1377 1328 48 1298 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $32832 m0 *1 858.36,111.52
X$32832 48 1190 1328 1297 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $32833 m0 *1 859.74,111.52
X$32833 29 1336 1498 1190 1328 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $32835 m0 *1 862.5,111.52
X$32835 29 1149 1492 1300 1384 48 48 29 sky130_fd_sc_hd__a21boi_2
* cell instance $32837 m0 *1 867.1,111.52
X$32837 29 1387 1023 1266 1329 1385 1386 48 48 29 sky130_fd_sc_hd__a221oi_2
* cell instance $32838 m0 *1 872.62,111.52
X$32838 48 1148 1234 1333 1330 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $33415 r0 *1 682.64,111.52
X$33415 48 1279 1165 1008 29 48 1456 29 sky130_fd_sc_hd__a21boi_0
* cell instance $33416 r0 *1 685.4,111.52
X$33416 48 1008 1217 1494 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33418 r0 *1 687.24,111.52
X$33418 29 1362 1067 1105 1460 1497 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $33421 r0 *1 695.52,111.52
X$33421 48 1008 1067 1217 29 48 1461 29 sky130_fd_sc_hd__a21oi_1
* cell instance $33423 r0 *1 697.82,111.52
X$33423 29 1655 1406 1132 1407 1195 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $33424 r0 *1 701.04,111.52
X$33424 48 981 1133 1406 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33425 r0 *1 702.42,111.52
X$33425 48 1133 981 1465 1132 29 1395 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $33427 r0 *1 705.64,111.52
X$33427 29 1407 1363 1275 1039 48 48 29 sky130_fd_sc_hd__nor3b_2
* cell instance $33428 r0 *1 710.24,111.52
X$33428 48 934 1244 1465 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33429 r0 *1 711.62,111.52
X$33429 48 890 1347 1284 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $33430 r0 *1 713,111.52
X$33430 29 1222 1223 937 1408 48 1363 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $33432 r0 *1 720.82,111.52
X$33432 48 1347 934 1244 48 29 1408 29 sky130_fd_sc_hd__o21ai_1
* cell instance $33433 r0 *1 722.66,111.52
X$33433 48 1165 1277 1350 48 29 1442 29 sky130_fd_sc_hd__o21ai_1
* cell instance $33434 r0 *1 724.5,111.52
X$33434 29 1277 1440 1013 1108 48 48 1350 29 sky130_fd_sc_hd__or4b_1
* cell instance $33436 r0 *1 729.1,111.52
X$33436 48 1257 981 1133 1410 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $33439 r0 *1 733.24,111.52
X$33439 48 1218 1409 1410 29 1469 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $33440 r0 *1 736.46,111.52
X$33440 48 1314 1219 1409 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33442 r0 *1 738.3,111.52
X$33442 48 1411 1225 1433 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $33443 r0 *1 740.6,111.52
X$33443 48 1225 1411 1434 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33447 r0 *1 744.28,111.52
X$33447 29 1178 1481 1444 1355 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $33449 r0 *1 747.96,111.52
X$33449 48 1178 1435 1314 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $33450 r0 *1 749.34,111.52
X$33450 48 1444 1227 1413 762 1436 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $33451 r0 *1 752.1,111.52
X$33451 48 1473 1273 1403 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $33453 r0 *1 756.24,111.52
X$33453 48 1142 1178 1089 1414 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $33454 r0 *1 758.08,111.52
X$33454 48 1117 1414 1474 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $33457 r0 *1 761.76,111.52
X$33457 48 1089 1142 1435 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $33458 r0 *1 764.06,111.52
X$33458 29 1321 1480 1287 48 48 29 sky130_fd_sc_hd__nor2_8
* cell instance $33459 r0 *1 771.42,111.52
X$33459 29 1036 1372 1375 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $33461 r0 *1 777.4,111.52
X$33461 48 1438 1415 1439 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33462 r0 *1 778.78,111.52
X$33462 29 2469 1142 1214 1271 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $33463 r0 *1 783.38,111.52
X$33463 29 1371 1321 1188 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $33466 r0 *1 788.44,111.52
X$33466 29 1271 1437 1270 1247 48 48 29 sky130_fd_sc_hd__ha_1
* cell instance $33467 r0 *1 793.04,111.52
X$33467 48 1417 1484 1416 1478 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $33468 r0 *1 794.88,111.52
X$33468 48 1699 1752 1400 1477 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $33470 r0 *1 797.18,111.52
X$33470 48 1376 29 1190 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $33471 r0 *1 799.94,111.52
X$33471 48 1398 1418 1419 29 48 1476 29 sky130_fd_sc_hd__a21oi_1
* cell instance $33473 r0 *1 801.78,111.52
X$33473 48 1354 1307 1472 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $33474 r0 *1 804.08,111.52
X$33474 48 1376 1119 1118 1419 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $33475 r0 *1 805.92,111.52
X$33475 48 1321 29 1305 48 29 sky130_fd_sc_hd__buf_2
* cell instance $33477 r0 *1 808.22,111.52
X$33477 29 1380 1378 1379 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $33482 r0 *1 816.5,111.52
X$33482 48 1346 1290 1508 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $33483 r0 *1 817.88,111.52
X$33483 48 1158 1349 1242 1348 1305 1470 29 48 29 sky130_fd_sc_hd__a32oi_1
* cell instance $33485 r0 *1 822.02,111.52
X$33485 48 1537 1346 1290 1448 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $33486 r0 *1 824.32,111.52
X$33486 48 1352 1290 1432 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33489 r0 *1 828,111.52
X$33489 48 1324 1303 1448 1294 1449 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $33491 r0 *1 830.76,111.52
X$33491 48 1325 1388 1345 48 1420 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $33492 r0 *1 833.98,111.52
X$33492 48 1327 1291 1240 1303 48 1451 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $33493 r0 *1 836.28,111.52
X$33493 29 1381 1420 1421 1295 48 1818 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $33494 r0 *1 840.88,111.52
X$33494 29 29 1452 48 1326 1341 48 sky130_fd_sc_hd__nor2_2
* cell instance $33496 r0 *1 843.64,111.52
X$33496 48 1341 1326 1466 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $33499 r0 *1 848.7,111.52
X$33499 48 1452 1421 1464 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $33500 r0 *1 850.08,111.52
X$33500 48 1422 1111 1431 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $33502 r0 *1 851.92,111.52
X$33502 48 1421 1452 1423 29 48 1462 29 sky130_fd_sc_hd__a21boi_0
* cell instance $33503 r0 *1 854.68,111.52
X$33503 48 1500 1491 1474 29 48 1425 29 sky130_fd_sc_hd__a21o_1
* cell instance $33505 r0 *1 857.44,111.52
X$33505 29 1454 1424 1425 1300 1384 1190 1153 48 48 29 sky130_fd_sc_hd__a222oi_1
* cell instance $33507 r0 *1 862.04,111.52
X$33507 29 1336 1426 1194 1191 1455 48 48 29 sky130_fd_sc_hd__nor4_4
* cell instance $33510 r0 *1 871.24,111.52
X$33510 48 1230 48 29 1459 29 sky130_fd_sc_hd__inv_1
* cell instance $33511 r0 *1 872.62,111.52
X$33511 48 1430 1426 1429 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $33513 r0 *1 874.46,111.52
X$33513 48 1427 1428 1429 29 48 1457 29 sky130_fd_sc_hd__a21oi_1
* cell instance $34142 m0 *1 681.26,116.96
X$34142 29 1680 931 1128 1456 1165 1390 48 48 29 sky130_fd_sc_hd__o32a_1
* cell instance $34143 m0 *1 684.94,116.96
X$34143 48 1494 1131 1283 48 1495 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $34149 m0 *1 692.3,116.96
X$34149 29 1497 1008 1105 1132 981 1133 48 48 29 sky130_fd_sc_hd__a2111oi_2
* cell instance $34153 m0 *1 698.28,116.96
X$34153 29 1258 1132 1133 981 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $34155 m0 *1 704.72,116.96
X$34155 48 1406 1195 1499 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34157 m0 *1 707.94,116.96
X$34157 48 1132 1223 981 1133 48 1366 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $34158 m0 *1 711.16,116.96
X$34158 48 934 1347 1547 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34160 m0 *1 713,116.96
X$34160 29 1479 1397 861 1218 1222 1244 48 48 29 sky130_fd_sc_hd__a41oi_2
* cell instance $34162 m0 *1 719.44,116.96
X$34162 48 861 1013 1369 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $34165 m0 *1 720.82,116.96
X$34165 48 1440 1406 1399 1441 1502 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $34166 m0 *1 724.04,116.96
X$34166 48 1067 1441 1277 1503 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $34169 m0 *1 727.72,116.96
X$34169 29 1407 1219 1218 1468 1443 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $34170 m0 *1 735.54,116.96
X$34170 29 1469 1080 1551 1355 1481 1067 48 48 29 sky130_fd_sc_hd__a221oi_4
* cell instance $34174 m0 *1 747.04,116.96
X$34174 48 1444 1227 1358 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $34177 m0 *1 748.42,116.96
X$34177 48 762 1178 1471 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $34178 m0 *1 751.64,116.96
X$34178 48 1480 815 1471 1513 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $34179 m0 *1 753.48,116.96
X$34179 48 1178 1444 1252 48 1473 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $34181 m0 *1 756.24,116.96
X$34181 48 1435 29 1444 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34182 m0 *1 759,116.96
X$34182 48 1370 1474 1413 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34183 m0 *1 760.38,116.96
X$34183 48 1435 1194 1475 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $34184 m0 *1 761.76,116.96
X$34184 29 29 1289 1139 1445 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $34185 m0 *1 764.06,116.96
X$34185 48 1291 1474 1507 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $34186 m0 *1 765.44,116.96
X$34186 48 1483 1438 1736 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34203 m0 *1 778.78,116.96
X$34203 48 1412 29 319 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34204 m0 *1 781.54,116.96
X$34204 48 1261 29 368 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34215 m0 *1 793.5,116.96
X$34215 29 1447 1262 1478 1417 1446 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $34216 m0 *1 798.1,116.96
X$34216 48 1416 1119 1446 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $34221 m0 *1 802.24,116.96
X$34221 29 1447 1353 1417 1418 1242 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $34222 m0 *1 809.6,116.96
X$34222 48 1118 1379 1510 1509 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $34224 m0 *1 812.36,116.96
X$34224 48 1373 29 1450 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34227 m0 *1 817.42,116.96
X$34227 29 1488 1508 1487 1352 1392 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $34230 m0 *1 823.4,116.96
X$34230 29 1506 1488 1380 1505 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $34234 m0 *1 829.84,116.96
X$34234 48 1303 1324 1294 1448 48 1467 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $34235 m0 *1 833.06,116.96
X$34235 29 29 1448 1327 1294 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $34236 m0 *1 835.36,116.96
X$34236 48 1240 1449 1451 48 1382 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $34237 m0 *1 837.2,116.96
X$34237 48 1576 1618 1291 29 1463 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $34238 m0 *1 840.42,116.96
X$34238 48 1326 1341 1472 29 1504 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $34240 m0 *1 844.56,116.96
X$34240 48 1421 1466 1453 1501 29 48 29 sky130_fd_sc_hd__nor3b_1
* cell instance $34241 m0 *1 847.32,116.96
X$34241 48 1421 1452 1453 29 48 1490 29 sky130_fd_sc_hd__a21oi_1
* cell instance $34242 m0 *1 849.16,116.96
X$34242 29 1423 1421 1452 1455 1490 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $34247 m0 *1 857.9,116.96
X$34247 29 1526 1194 1300 1498 1613 1561 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $34249 m0 *1 868.02,116.96
X$34249 48 1430 1426 1492 1496 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $34251 m0 *1 870.78,116.96
X$34251 29 1492 1458 1426 1430 1520 1521 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $34936 r0 *1 681.72,116.96
X$34936 29 1008 1511 1217 1131 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $34937 r0 *1 685.4,116.96
X$34937 29 1495 1511 1393 1568 1569 48 1523 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $34941 r0 *1 695.06,116.96
X$34941 29 1165 1105 1546 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $34948 r0 *1 718.98,116.96
X$34948 48 1258 29 1165 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34952 r0 *1 721.74,116.96
X$34952 48 1184 980 1441 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34953 r0 *1 723.12,116.96
X$34953 48 1165 1277 1350 1579 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $34954 r0 *1 725.42,116.96
X$34954 48 1407 1219 1528 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $34958 r0 *1 733.24,116.96
X$34958 48 640 1443 1529 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $34960 r0 *1 736,116.96
X$34960 29 1469 1067 1530 1080 1355 1481 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $34961 r0 *1 739.68,116.96
X$34961 29 1482 1593 1480 1258 1532 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $34965 r0 *1 747.5,116.96
X$34965 48 1257 48 29 1533 29 sky130_fd_sc_hd__inv_1
* cell instance $34967 r0 *1 749.34,116.96
X$34967 48 1513 1319 48 1482 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $34970 r0 *1 753.94,116.96
X$34970 29 1257 1232 1444 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $34972 r0 *1 759,116.96
X$34972 48 1483 1554 1535 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $34974 r0 *1 760.84,116.96
X$34974 48 1140 29 1376 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34976 r0 *1 764.06,116.96
X$34976 29 1372 1036 1638 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $34986 r0 *1 779.7,116.96
X$34986 48 1404 29 576 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $34994 r0 *1 788.44,116.96
X$34994 29 29 1514 48 1321 1354 48 sky130_fd_sc_hd__nor2_2
* cell instance $34995 r0 *1 790.74,116.96
X$34995 29 29 1475 1515 1373 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $34996 r0 *1 793.04,116.96
X$34996 48 1118 1516 1378 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $34997 r0 *1 794.42,116.96
X$34997 48 1517 1599 1543 48 1544 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $34998 r0 *1 797.64,116.96
X$34998 48 1446 1398 1376 1476 29 48 1292 29 sky130_fd_sc_hd__a31oi_1
* cell instance $34999 r0 *1 799.94,116.96
X$34999 48 1484 48 29 1119 29 sky130_fd_sc_hd__clkinvlp_4
* cell instance $35003 r0 *1 802.7,116.96
X$35003 48 1484 1416 1418 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35005 r0 *1 804.54,116.96
X$35005 48 1416 1485 1396 1486 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $35006 r0 *1 806.38,116.96
X$35006 48 1396 1194 1305 1485 29 1542 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $35007 r0 *1 808.68,116.96
X$35007 48 1510 1379 1644 1540 29 1541 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $35009 r0 *1 811.9,116.96
X$35009 48 1509 1486 1287 29 1538 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $35012 r0 *1 816.04,116.96
X$35012 48 1509 1291 1486 48 29 1539 29 sky130_fd_sc_hd__o21ai_1
* cell instance $35021 r0 *1 830.3,116.96
X$35021 48 1449 1305 1240 1467 48 1536 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $35022 r0 *1 832.6,116.96
X$35022 48 1450 1383 1327 1534 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $35023 r0 *1 834.44,116.96
X$35023 48 1327 1344 1450 1489 1667 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $35024 r0 *1 837.2,116.96
X$35024 48 1291 1327 1344 1559 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $35025 r0 *1 839.04,116.96
X$35025 48 1324 1489 1303 29 48 1531 29 sky130_fd_sc_hd__a21oi_1
* cell instance $35029 r0 *1 843.64,116.96
X$35029 29 1452 1422 1423 1615 1567 48 1336 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $35030 r0 *1 853.3,116.96
X$35030 29 1519 1336 1462 1501 48 48 29 sky130_fd_sc_hd__o21bai_2
* cell instance $35034 r0 *1 857.44,116.96
X$35034 48 1500 1111 1491 1424 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $35036 r0 *1 859.74,116.96
X$35036 48 1336 1190 1328 29 48 1526 29 sky130_fd_sc_hd__a21oi_1
* cell instance $35038 r0 *1 862.04,116.96
X$35038 29 1430 1455 1525 1056 48 48 29 sky130_fd_sc_hd__a21boi_4
* cell instance $35039 r0 *1 868.94,116.96
X$35039 48 1524 1234 1496 48 1522 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $35041 r0 *1 871.24,116.96
X$35041 29 1459 1493 1426 1430 1520 1521 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $35681 m0 *1 680.8,122.4
X$35681 48 931 1165 1179 48 29 1569 29 sky130_fd_sc_hd__or3_2
* cell instance $35682 m0 *1 683.56,122.4
X$35682 48 1165 1179 931 29 1568 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $35684 m0 *1 687.7,122.4
X$35684 29 1495 1612 1511 1393 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $35686 m0 *1 691.84,122.4
X$35686 29 1281 1163 1545 48 1570 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $35687 m0 *1 698.28,122.4
X$35687 29 1461 1545 1274 1364 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $35688 m0 *1 701.96,122.4
X$35688 48 1546 1274 1461 48 1616 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $35689 m0 *1 704.72,122.4
X$35689 48 1340 1394 1547 1590 29 48 29 sky130_fd_sc_hd__nand3b_1
* cell instance $35690 m0 *1 707.48,122.4
X$35690 29 1394 1548 1547 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $35693 m0 *1 713,122.4
X$35693 48 1503 1502 1658 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35694 m0 *1 714.38,122.4
X$35694 48 1502 1503 1479 1549 29 1577 48 29 sky130_fd_sc_hd__a22o_1
* cell instance $35695 m0 *1 717.6,122.4
X$35695 48 1479 1549 1550 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35697 m0 *1 719.44,122.4
X$35697 48 1185 1503 1502 29 48 1623 29 sky130_fd_sc_hd__a21oi_1
* cell instance $35698 m0 *1 721.28,122.4
X$35698 29 1578 1184 1442 1579 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $35699 m0 *1 724.96,122.4
X$35699 48 1442 1579 1582 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35700 m0 *1 726.34,122.4
X$35700 48 1529 1218 1528 48 29 1660 29 sky130_fd_sc_hd__a21o_2
* cell instance $35701 m0 *1 729.56,122.4
X$35701 48 1218 1528 1624 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35704 m0 *1 732.32,122.4
X$35704 48 1530 29 1552 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $35705 m0 *1 735.08,122.4
X$35705 48 1551 941 1690 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35706 m0 *1 736.46,122.4
X$35706 48 1444 1552 1512 48 29 1553 29 sky130_fd_sc_hd__o21ai_1
* cell instance $35708 m0 *1 738.76,122.4
X$35708 48 1480 1552 1583 29 48 1626 29 sky130_fd_sc_hd__a21oi_1
* cell instance $35709 m0 *1 740.6,122.4
X$35709 48 1583 29 1512 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $35710 m0 *1 743.36,122.4
X$35710 48 1532 1482 1258 1480 29 48 1584 29 sky130_fd_sc_hd__or4_2
* cell instance $35712 m0 *1 747.04,122.4
X$35712 29 29 1041 48 1140 1533 48 sky130_fd_sc_hd__nor2_2
* cell instance $35713 m0 *1 749.34,122.4
X$35713 48 1355 1533 1532 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $35717 m0 *1 755.32,122.4
X$35717 48 1480 48 29 1324 29 sky130_fd_sc_hd__buf_4
* cell instance $35718 m0 *1 758.08,122.4
X$35718 48 1444 48 29 1262 29 sky130_fd_sc_hd__buf_4
* cell instance $35719 m0 *1 760.84,122.4
X$35719 48 1376 1474 1483 48 1555 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $35720 m0 *1 764.06,122.4
X$35720 48 1555 1554 1586 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $35722 m0 *1 766.36,122.4
X$35722 29 1377 1480 1140 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $35723 m0 *1 770.5,122.4
X$35723 29 1595 1291 1639 1031 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $35725 m0 *1 774.64,122.4
X$35725 48 1507 1438 1625 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $35726 m0 *1 777.86,122.4
X$35726 29 1485 1516 1556 1312 48 48 29 sky130_fd_sc_hd__xnor3_2
* cell instance $35727 m0 *1 786.6,122.4
X$35727 29 1556 1312 1379 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $35728 m0 *1 796.72,122.4
X$35728 29 1262 1417 1484 1510 1557 48 48 29 sky130_fd_sc_hd__o31ai_2
* cell instance $35732 m0 *1 803.16,122.4
X$35732 29 1732 1585 1510 1379 1194 1321 48 48 29 sky130_fd_sc_hd__o41ai_1
* cell instance $35734 m0 *1 807.3,122.4
X$35734 29 1558 1416 1638 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $35735 m0 *1 813.28,122.4
X$35735 29 1622 1509 1486 1450 1377 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $35736 m0 *1 816.96,122.4
X$35736 29 1581 1604 1580 1539 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $35740 m0 *1 823.86,122.4
X$35740 48 1352 1293 1538 48 29 1605 29 sky130_fd_sc_hd__a21boi_1
* cell instance $35741 m0 *1 826.62,122.4
X$35741 48 1537 1352 1538 1606 29 48 29 sky130_fd_sc_hd__nor3b_1
* cell instance $35744 m0 *1 830.3,122.4
X$35744 48 1646 1534 1536 48 29 1566 29 sky130_fd_sc_hd__a21o_2
* cell instance $35746 m0 *1 833.98,122.4
X$35746 48 1489 1344 1576 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $35748 m0 *1 835.82,122.4
X$35748 48 1240 1647 1575 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35750 m0 *1 838.12,122.4
X$35750 48 1305 1559 1575 1573 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $35751 m0 *1 839.96,122.4
X$35751 48 1531 1327 1559 1489 1609 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $35752 m0 *1 843.18,122.4
X$35752 48 1518 1571 1572 48 29 1423 29 sky130_fd_sc_hd__or3_2
* cell instance $35754 m0 *1 846.4,122.4
X$35754 48 1466 1609 1567 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35756 m0 *1 848.24,122.4
X$35756 29 1453 1464 1339 48 1560 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $35757 m0 *1 853.3,122.4
X$35757 48 1453 29 1026 48 29 sky130_fd_sc_hd__buf_2
* cell instance $35758 m0 *1 855.14,122.4
X$35758 48 1566 1026 1614 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $35762 m0 *1 857.9,122.4
X$35762 48 1026 1561 1491 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $35764 m0 *1 859.74,122.4
X$35764 29 29 1560 1821 1377 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $35766 m0 *1 862.5,122.4
X$35766 29 29 1525 48 1194 1336 48 sky130_fd_sc_hd__nor2_2
* cell instance $35768 m0 *1 865.26,122.4
X$35768 48 1562 48 29 1563 29 sky130_fd_sc_hd__inv_1
* cell instance $35770 m0 *1 867.1,122.4
X$35770 48 1563 1056 1565 48 29 1520 29 sky130_fd_sc_hd__a21o_2
* cell instance $35771 m0 *1 870.32,122.4
X$35771 29 1564 1148 1427 1458 1454 1493 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $35773 m0 *1 880.9,122.4
X$35773 48 1520 1521 1611 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $36372 r0 *1 681.72,122.4
X$36372 48 1568 1569 1652 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36373 r0 *1 683.1,122.4
X$36373 48 1568 1128 1569 48 1587 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $36375 r0 *1 686.78,122.4
X$36375 29 1612 1527 1588 1587 1460 48 1657 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $36379 r0 *1 696.9,122.4
X$36379 48 1628 1162 1620 48 29 1589 29 sky130_fd_sc_hd__o21ai_1
* cell instance $36380 r0 *1 698.74,122.4
X$36380 48 1274 1461 1617 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $36382 r0 *1 701.5,122.4
X$36382 48 1617 29 1619 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $36385 r0 *1 705.64,122.4
X$36385 48 1590 1552 1591 1577 29 1620 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $36386 r0 *1 707.94,122.4
X$36386 48 1530 1591 1577 48 29 1574 29 sky130_fd_sc_hd__or3_2
* cell instance $36387 r0 *1 710.7,122.4
X$36387 48 937 1547 1394 1723 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $36389 r0 *1 713.46,122.4
X$36389 48 1551 1658 1588 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36390 r0 *1 714.84,122.4
X$36390 48 1630 1550 1527 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36391 r0 *1 716.22,122.4
X$36391 48 1479 1549 48 1632 29 29 sky130_fd_sc_hd__and2_2
* cell instance $36392 r0 *1 718.98,122.4
X$36392 48 1503 1502 1185 29 48 1631 29 sky130_fd_sc_hd__a21o_1
* cell instance $36396 r0 *1 722.66,122.4
X$36396 29 1725 1550 1591 1552 1578 1623 48 48 29 sky130_fd_sc_hd__a2111o_1
* cell instance $36397 r0 *1 726.8,122.4
X$36397 29 1661 1140 1631 1632 1552 1591 48 48 29 sky130_fd_sc_hd__o41ai_1
* cell instance $36400 r0 *1 731.4,122.4
X$36400 48 1184 1582 1662 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36402 r0 *1 733.24,122.4
X$36402 48 1592 1633 1663 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36403 r0 *1 734.62,122.4
X$36403 48 1592 1630 1665 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36405 r0 *1 736.92,122.4
X$36405 48 1691 1666 1634 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $36406 r0 *1 739.22,122.4
X$36406 48 1551 941 1635 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $36407 r0 *1 740.6,122.4
X$36407 29 1584 1593 1318 48 1591 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $36408 r0 *1 747.04,122.4
X$36408 48 1475 1594 1636 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36411 r0 *1 748.42,122.4
X$36411 48 1593 1584 1594 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36414 r0 *1 751.18,122.4
X$36414 29 1882 1413 1669 1670 1637 1444 48 48 29 sky130_fd_sc_hd__o41a_1
* cell instance $36416 r0 *1 755.78,122.4
X$36416 29 29 1592 1108 1445 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $36418 r0 *1 759,122.4
X$36418 48 1592 1438 1554 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36420 r0 *1 760.84,122.4
X$36420 29 29 1592 48 1375 1515 48 sky130_fd_sc_hd__nor2_2
* cell instance $36421 r0 *1 763.14,122.4
X$36421 29 1287 1224 1638 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $36422 r0 *1 767.28,122.4
X$36422 48 1445 1638 1514 29 48 1185 29 sky130_fd_sc_hd__and3_2
* cell instance $36424 r0 *1 770.5,122.4
X$36424 48 1475 29 1291 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $36425 r0 *1 773.26,122.4
X$36425 48 1639 1625 1675 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36428 r0 *1 774.64,122.4
X$36428 29 1595 1438 1312 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $36429 r0 *1 784.76,122.4
X$36429 48 1291 1641 1477 29 48 1556 29 sky130_fd_sc_hd__o21a_2
* cell instance $36431 r0 *1 788.44,122.4
X$36431 48 1596 1597 1598 29 48 1641 29 sky130_fd_sc_hd__a21oi_1
* cell instance $36432 r0 *1 790.28,122.4
X$36432 48 1597 1598 1678 1698 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $36433 r0 *1 792.12,122.4
X$36433 48 1262 1679 1417 48 1557 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $36434 r0 *1 793.96,122.4
X$36434 48 1517 1543 1323 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $36435 r0 *1 796.26,122.4
X$36435 48 1323 1599 1700 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $36436 r0 *1 798.56,122.4
X$36436 29 1643 1544 1585 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $36439 r0 *1 804.54,122.4
X$36439 29 1600 1701 1485 1396 1643 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $36440 r0 *1 809.14,122.4
X$36440 48 1542 1644 1676 48 29 1601 29 sky130_fd_sc_hd__o21ai_1
* cell instance $36442 r0 *1 811.9,122.4
X$36442 48 1585 48 29 1540 29 sky130_fd_sc_hd__clkinvlp_4
* cell instance $36445 r0 *1 816.04,122.4
X$36445 48 1602 1603 1558 1604 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $36446 r0 *1 817.88,122.4
X$36446 48 1305 1581 1621 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $36447 r0 *1 819.26,122.4
X$36447 29 1672 1604 1580 1538 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $36448 r0 *1 822.94,122.4
X$36448 48 1538 1558 1671 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $36450 r0 *1 828,122.4
X$36450 48 1605 1606 1646 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $36453 r0 *1 829.38,122.4
X$36453 48 1489 1305 1467 29 48 1668 29 sky130_fd_sc_hd__a21oi_1
* cell instance $36454 r0 *1 831.22,122.4
X$36454 48 1450 1489 1291 1327 1344 1607 29 48 29 sky130_fd_sc_hd__a311o_1
* cell instance $36455 r0 *1 834.9,122.4
X$36455 48 1667 1647 1607 48 1608 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $36456 r0 *1 838.12,122.4
X$36456 48 1240 1303 1618 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $36457 r0 *1 839.5,122.4
X$36457 48 1609 1381 1421 1648 29 48 1664 29 sky130_fd_sc_hd__a31oi_1
* cell instance $36461 r0 *1 843.64,122.4
X$36461 29 1571 1518 1572 1609 1463 48 1615 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $36462 r0 *1 853.3,122.4
X$36462 29 1648 1614 1610 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $36465 r0 *1 859.28,122.4
X$36465 48 1377 1560 1714 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $36466 r0 *1 861.58,122.4
X$36466 29 1650 1613 1821 1562 1561 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $36467 r0 *1 866.18,122.4
X$36467 48 1610 1650 48 1524 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $36471 r0 *1 871.24,122.4
X$36471 29 1521 1056 1563 1565 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $36472 r0 *1 874.92,122.4
X$36472 29 1656 1524 1611 1457 1234 1496 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $36473 r0 *1 878.14,122.4
X$36473 48 1454 1493 1653 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $36474 r0 *1 879.52,122.4
X$36474 48 1520 1521 1428 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37110 m0 *1 682.18,127.84
X$37110 29 1612 1768 1574 1545 1627 1680 48 48 29 sky130_fd_sc_hd__a221oi_2
* cell instance $37111 m0 *1 687.7,127.84
X$37111 29 1545 1680 1681 1612 1574 1627 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $37113 m0 *1 691.84,127.84
X$37113 29 1688 1655 1523 1163 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $37115 m0 *1 697.82,127.84
X$37115 48 1162 1620 1628 48 1887 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $37116 m0 *1 700.58,127.84
X$37116 29 1720 1684 1616 1629 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $37117 m0 *1 704.26,127.84
X$37117 48 1162 1628 1499 1686 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $37118 m0 *1 706.1,127.84
X$37118 48 1591 1530 1577 1590 1685 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $37121 m0 *1 711.16,127.84
X$37121 48 1723 1552 1591 1577 29 1629 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $37123 m0 *1 714.38,127.84
X$37123 29 1726 1632 1551 1630 1631 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $37127 m0 *1 720.36,127.84
X$37127 29 1725 1688 1689 1744 1578 1570 48 48 29 sky130_fd_sc_hd__o32ai_4
* cell instance $37128 m0 *1 730.48,127.84
X$37128 29 1578 1728 1662 1633 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $37129 m0 *1 738.76,127.84
X$37129 29 1692 1729 1730 1636 1634 1635 48 48 29 sky130_fd_sc_hd__o311a_4
* cell instance $37131 m0 *1 747.04,127.84
X$37131 48 1318 1593 1584 29 48 1630 29 sky130_fd_sc_hd__and3_2
* cell instance $37135 m0 *1 752.1,127.84
X$37135 29 1734 1637 1438 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $37136 m0 *1 762.22,127.84
X$37136 48 1693 1735 1639 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $37138 m0 *1 765.9,127.84
X$37138 29 1483 1415 1555 1031 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $37141 m0 *1 774.64,127.84
X$37141 48 1674 1483 1738 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $37142 m0 *1 777.86,127.84
X$37142 29 29 1647 48 1291 1694 48 sky130_fd_sc_hd__nor2_2
* cell instance $37144 m0 *1 781.08,127.84
X$37144 48 1400 1312 48 1640 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $37145 m0 *1 784.3,127.84
X$37145 48 1287 1640 1599 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $37146 m0 *1 786.6,127.84
X$37146 29 1677 1696 1737 1739 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $37147 m0 *1 788.9,127.84
X$37147 48 1642 1417 1599 1678 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $37148 m0 *1 791.2,127.84
X$37148 48 1398 1597 1598 1543 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $37149 m0 *1 793.04,127.84
X$37149 29 1733 1585 1642 1484 1792 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $37153 m0 *1 802.24,127.84
X$37153 29 1701 1732 1673 1540 1700 48 48 29 sky130_fd_sc_hd__a22oi_2
* cell instance $37155 m0 *1 807.3,127.84
X$37155 29 1514 1541 1702 1731 1645 1600 48 48 29 sky130_fd_sc_hd__o2111ai_4
* cell instance $37156 m0 *1 816.96,127.84
X$37156 48 1450 1704 1706 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37158 m0 *1 819.26,127.84
X$37158 29 1707 1580 1450 1706 1702 1604 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $37159 m0 *1 822.48,127.84
X$37159 48 1537 1672 1727 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37161 m0 *1 824.32,127.84
X$37161 29 1707 1782 1487 1671 1325 1305 48 48 29 sky130_fd_sc_hd__o32ai_1
* cell instance $37162 m0 *1 827.54,127.84
X$37162 48 1605 1450 1606 48 29 1709 29 sky130_fd_sc_hd__o21ai_1
* cell instance $37166 m0 *1 831.68,127.84
X$37166 29 1649 1668 1646 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $37170 m0 *1 840.88,127.84
X$37170 29 1724 1664 1572 1518 1571 1422 48 48 29 sky130_fd_sc_hd__o41ai_2
* cell instance $37174 m0 *1 850.08,127.84
X$37174 48 1649 1608 1722 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $37175 m0 *1 852.38,127.84
X$37175 48 1453 1608 1659 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37181 m0 *1 857.44,127.84
X$37181 48 1659 1649 48 1562 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $37184 m0 *1 863.42,127.84
X$37184 29 1427 1610 1650 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $37185 m0 *1 869.4,127.84
X$37185 48 1427 1458 1715 1719 29 48 29 sky130_fd_sc_hd__nor3b_1
* cell instance $37186 m0 *1 872.16,127.84
X$37186 29 1522 1716 1387 1864 1428 1651 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $37187 m0 *1 875.84,127.84
X$37187 29 1716 1653 1654 1717 1718 48 48 29 sky130_fd_sc_hd__a2bb2oi_1
* cell instance $37188 m0 *1 879.06,127.84
X$37188 48 1458 1427 1654 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37845 r0 *1 684.48,127.84
X$37845 29 1682 1928 1768 1740 1583 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $37846 r0 *1 692.3,127.84
X$37846 48 931 1128 1460 48 29 1628 29 sky130_fd_sc_hd__o21ai_1
* cell instance $37850 r0 *1 694.14,127.84
X$37850 29 1691 1683 1583 1657 1681 48 48 29 sky130_fd_sc_hd__a211o_4
* cell instance $37851 r0 *1 700.58,127.84
X$37851 29 1683 937 1741 1574 1684 1742 48 48 29 sky130_fd_sc_hd__o221a_1
* cell instance $37854 r0 *1 705.64,127.84
X$37854 48 1619 1546 1684 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37855 r0 *1 707.02,127.84
X$37855 48 1660 1685 1686 29 48 1743 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37856 r0 *1 708.86,127.84
X$37856 29 1742 1591 1530 1577 1548 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $37858 r0 *1 714.38,127.84
X$37858 29 1687 1591 1552 1632 1631 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $37859 r0 *1 718.98,127.84
X$37859 48 1630 1552 1775 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37863 r0 *1 720.36,127.84
X$37863 29 1570 1726 1689 1688 1633 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $37864 r0 *1 727.72,127.84
X$37864 29 29 1551 1689 1630 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $37867 r0 *1 731.4,127.84
X$37867 48 1745 1690 1956 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37869 r0 *1 733.24,127.84
X$37869 29 1570 1779 1661 1688 1444 48 48 29 sky130_fd_sc_hd__o22ai_2
* cell instance $37870 r0 *1 737.84,127.84
X$37870 48 1830 1551 941 1916 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $37871 r0 *1 739.68,127.84
X$37871 48 1594 1691 1666 1690 48 1729 29 29 sky130_fd_sc_hd__nand4b_1
* cell instance $37872 r0 *1 742.9,127.84
X$37872 48 1626 1594 1636 1690 1730 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $37873 r0 *1 746.12,127.84
X$37873 29 1746 1692 1694 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $37877 r0 *1 756.24,127.84
X$37877 48 1670 1262 1785 48 1693 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $37880 r0 *1 760.84,127.84
X$37880 29 1693 1669 1483 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $37881 r0 *1 770.96,127.84
X$37881 29 1807 1675 1736 1031 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $37885 r0 *1 775.1,127.84
X$37885 29 1790 1287 1789 1792 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $37886 r0 *1 781.08,127.84
X$37886 48 1695 1748 1791 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37888 r0 *1 783.38,127.84
X$37888 29 1515 1739 1398 1640 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $37891 r0 *1 788.44,127.84
X$37891 48 1793 1696 1750 1697 1749 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $37892 r0 *1 790.74,127.84
X$37892 48 1795 1698 1749 29 48 1796 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37893 r0 *1 792.58,127.84
X$37893 48 1375 29 1751 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $37894 r0 *1 795.34,127.84
X$37894 48 1752 1699 1678 48 29 1812 29 sky130_fd_sc_hd__or3_2
* cell instance $37896 r0 *1 799.94,127.84
X$37896 48 1262 1642 1794 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37897 r0 *1 801.32,127.84
X$37897 48 1416 1585 1700 48 29 1755 29 sky130_fd_sc_hd__o21ai_1
* cell instance $37901 r0 *1 803.16,127.84
X$37901 48 1416 1585 1700 1603 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $37902 r0 *1 805,127.84
X$37902 48 1540 1118 1544 29 48 1602 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37903 r0 *1 806.84,127.84
X$37903 48 1118 1540 1544 1705 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $37904 r0 *1 808.68,127.84
X$37904 48 1703 1705 1755 1645 29 48 1787 29 sky130_fd_sc_hd__and4_1
* cell instance $37906 r0 *1 812.36,127.84
X$37906 48 1540 1700 1676 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37907 r0 *1 813.74,127.84
X$37907 48 1703 1755 1705 29 48 1756 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37909 r0 *1 816.04,127.84
X$37909 48 1645 1703 1786 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37910 r0 *1 817.42,127.84
X$37910 48 1704 1755 1705 29 48 1580 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37911 r0 *1 819.26,127.84
X$37911 48 1580 1604 1487 29 48 1757 29 sky130_fd_sc_hd__a21oi_1
* cell instance $37913 r0 *1 821.56,127.84
X$37913 48 1727 1352 1558 1325 1759 48 29 29 sky130_fd_sc_hd__a31o_2
* cell instance $37914 r0 *1 824.78,127.84
X$37914 29 1704 1708 1352 1487 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $37916 r0 *1 827.54,127.84
X$37916 48 1780 1708 1710 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $37921 r0 *1 830.76,127.84
X$37921 48 1489 1709 1711 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37922 r0 *1 832.14,127.84
X$37922 29 1710 1711 1648 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $37926 r0 *1 845.48,127.84
X$37926 29 1648 1764 1566 1712 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $37928 r0 *1 848.24,127.84
X$37928 48 1649 1648 1713 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37930 r0 *1 850.54,127.84
X$37930 48 1649 1608 1774 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $37931 r0 *1 851.92,127.84
X$37931 29 1453 1713 1764 48 1765 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $37936 r0 *1 857.44,127.84
X$37936 29 1384 1721 1525 1773 1714 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $37937 r0 *1 862.04,127.84
X$37937 48 1519 1298 1771 48 1772 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $37938 r0 *1 863.88,127.84
X$37938 48 1298 1519 1565 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $37942 r0 *1 871.24,127.84
X$37942 48 1656 1770 1386 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $37944 r0 *1 873.08,127.84
X$37944 48 1656 1719 1653 1767 1385 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $37946 r0 *1 876.3,127.84
X$37946 48 1564 1654 1717 1651 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $38587 m0 *1 683.56,133.28
X$38587 48 1612 1545 1574 29 48 1769 29 sky130_fd_sc_hd__a21oi_1
* cell instance $38589 m0 *1 685.86,133.28
X$38589 48 1583 29 48 941 29 sky130_fd_sc_hd__inv_4
* cell instance $38590 m0 *1 688.16,133.28
X$38590 48 1688 1687 1570 29 48 1583 29 sky130_fd_sc_hd__o21a_2
* cell instance $38593 m0 *1 692.3,133.28
X$38593 29 1740 1612 1527 1588 1587 1460 48 48 29 sky130_fd_sc_hd__o311a_1
* cell instance $38595 m0 *1 696.9,133.28
X$38595 48 1683 1681 1657 29 48 1797 29 sky130_fd_sc_hd__a21oi_1
* cell instance $38597 m0 *1 699.2,133.28
X$38597 48 1741 1574 1684 1742 1823 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $38599 m0 *1 702.42,133.28
X$38599 48 1616 1548 1741 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $38601 m0 *1 705.18,133.28
X$38601 48 1685 1686 1826 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $38604 m0 *1 708.86,133.28
X$38604 48 1589 1743 1798 29 48 1666 29 sky130_fd_sc_hd__and3_2
* cell instance $38607 m0 *1 713,133.28
X$38607 48 1742 1691 1666 1827 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $38610 m0 *1 717.6,133.28
X$38610 48 1689 1577 1799 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $38612 m0 *1 719.44,133.28
X$38612 29 1744 1632 1912 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $38614 m0 *1 730.02,133.28
X$38614 29 1666 1691 1781 1778 1665 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $38616 m0 *1 738.3,133.28
X$38616 29 1232 1801 1553 1784 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $38618 m0 *1 747.04,133.28
X$38618 29 1634 1784 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $38619 m0 *1 751.18,133.28
X$38619 29 1692 1746 1637 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $38620 m0 *1 757.16,133.28
X$38620 48 1804 1090 1803 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $38621 m0 *1 758.54,133.28
X$38621 29 1734 1324 1735 1670 1785 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $38622 m0 *1 763.14,133.28
X$38622 29 1977 1535 1586 1674 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $38623 m0 *1 767.28,133.28
X$38623 29 1833 1555 1483 1747 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $38625 m0 *1 772.34,133.28
X$38625 48 1810 1806 1439 1790 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $38627 m0 *1 774.64,133.28
X$38627 48 1262 1738 1232 29 1748 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $38628 m0 *1 777.86,133.28
X$38628 29 1417 1811 1848 1748 48 48 29 sky130_fd_sc_hd__o21a_4
* cell instance $38629 m0 *1 783.38,133.28
X$38629 29 1642 1792 1677 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $38630 m0 *1 789.36,133.28
X$38630 48 1699 1417 1750 48 29 1517 29 sky130_fd_sc_hd__o21ai_1
* cell instance $38631 m0 *1 791.2,133.28
X$38631 48 1960 1796 1751 29 1753 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $38632 m0 *1 794.42,133.28
X$38632 29 1699 1752 1484 48 48 29 sky130_fd_sc_hd__nor2_8
* cell instance $38634 m0 *1 802.24,133.28
X$38634 48 1416 1751 1704 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $38635 m0 *1 805.46,133.28
X$38635 48 1416 1753 1754 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $38636 m0 *1 806.84,133.28
X$38636 29 1643 1815 1754 1788 1540 48 48 29 sky130_fd_sc_hd__a22oi_4
* cell instance $38637 m0 *1 814.66,133.28
X$38637 29 1831 1622 1352 1787 1756 1786 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $38638 m0 *1 817.88,133.28
X$38638 48 1602 1603 1758 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $38641 m0 *1 820.64,133.28
X$38641 48 1758 29 1352 48 29 sky130_fd_sc_hd__buf_2
* cell instance $38643 m0 *1 823.4,133.28
X$38643 48 1450 1757 1783 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $38645 m0 *1 825.7,133.28
X$38645 29 1761 1505 1783 1782 1817 1759 48 48 29 sky130_fd_sc_hd__a2111oi_1
* cell instance $38648 m0 *1 830.3,133.28
X$38648 48 1759 1505 1776 1709 1760 29 48 29 sky130_fd_sc_hd__nor4bb_1
* cell instance $38651 m0 *1 835.36,133.28
X$38651 48 1240 1760 1761 48 1762 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $38652 m0 *1 838.12,133.28
X$38652 48 1761 1240 1760 48 29 1828 29 sky130_fd_sc_hd__o21ai_1
* cell instance $38653 m0 *1 839.96,133.28
X$38653 29 1763 1518 1724 1820 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $38654 m0 *1 845.94,133.28
X$38654 48 1608 1649 1712 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $38655 m0 *1 849.16,133.28
X$38655 29 1765 1613 1566 1877 1648 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $38659 m0 *1 858.82,133.28
X$38659 29 1873 1721 1714 1766 1825 1519 48 48 29 sky130_fd_sc_hd__a41oi_2
* cell instance $38660 m0 *1 864.8,133.28
X$38660 48 1613 1565 1824 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $38663 m0 *1 868.94,133.28
X$38663 48 1822 1719 1866 48 1770 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $38664 m0 *1 870.78,133.28
X$38664 48 1767 1715 1564 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $38668 m0 *1 877.22,133.28
X$38668 48 1564 1717 1718 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $39295 r0 *1 684.48,133.28
X$39295 48 931 1460 941 48 1865 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $39296 r0 *1 686.32,133.28
X$39296 48 1128 1652 1835 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $39298 r0 *1 688.16,133.28
X$39298 29 1682 1570 1688 1835 1687 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $39303 r0 *1 693.68,133.28
X$39303 29 1868 1570 1687 1460 1688 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $39305 r0 *1 699.2,133.28
X$39305 48 941 1868 1720 48 1870 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $39308 r0 *1 703.8,133.28
X$39308 48 1619 48 29 1837 29 sky130_fd_sc_hd__inv_1
* cell instance $39311 r0 *1 706.1,133.28
X$39311 48 1797 937 1838 48 29 1871 29 sky130_fd_sc_hd__o21ai_1
* cell instance $39313 r0 *1 708.86,133.28
X$39313 48 1589 1743 1838 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $39315 r0 *1 710.7,133.28
X$39315 48 1784 29 960 48 29 sky130_fd_sc_hd__clkinv_4
* cell instance $39318 r0 *1 715.3,133.28
X$39318 29 1779 1689 1775 48 1876 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $39322 r0 *1 720.36,133.28
X$39322 29 1777 1551 1797 1838 1745 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $39323 r0 *1 723.58,133.28
X$39323 48 1139 1570 1688 48 1829 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $39324 r0 *1 725.42,133.28
X$39324 48 1799 1829 1800 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $39325 r0 *1 726.8,133.28
X$39325 48 1139 1570 1582 1878 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $39327 r0 *1 729.56,133.28
X$39327 48 1779 1551 1778 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $39329 r0 *1 733.24,133.28
X$39329 29 1935 1663 1582 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $39330 r0 *1 739.22,133.28
X$39330 29 1841 1777 1842 1830 1318 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $39331 r0 *1 742.44,133.28
X$39331 48 1515 1594 1830 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $39332 r0 *1 743.82,133.28
X$39332 48 1880 1376 1041 1843 29 1802 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $39333 r0 *1 746.58,133.28
X$39333 29 1832 1444 1669 1670 1785 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $39337 r0 *1 751.18,133.28
X$39337 29 1882 1917 1845 48 1805 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $39338 r0 *1 757.62,133.28
X$39338 48 1802 1803 1669 48 29 29 sky130_fd_sc_hd__or2_2
* cell instance $39341 r0 *1 760.84,133.28
X$39341 48 1785 1694 1670 1669 48 1845 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $39342 r0 *1 763.14,133.28
X$39342 48 1287 1438 1893 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $39343 r0 *1 764.52,133.28
X$39343 29 29 1846 1834 1847 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $39344 r0 *1 766.82,133.28
X$39344 48 1810 1806 2046 29 1886 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $39345 r0 *1 770.04,133.28
X$39345 48 1807 1808 1809 29 48 1789 29 sky130_fd_sc_hd__a21oi_1
* cell instance $39346 r0 *1 771.88,133.28
X$39346 29 1811 1808 1809 1415 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $39350 r0 *1 775.56,133.28
X$39350 29 1748 1811 1695 1398 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $39351 r0 *1 781.54,133.28
X$39351 48 1415 1791 1596 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $39352 r0 *1 784.76,133.28
X$39352 48 1737 1677 1739 29 48 1793 29 sky130_fd_sc_hd__a21oi_1
* cell instance $39356 r0 *1 788.44,133.28
X$39356 29 1699 1750 1739 1677 48 1850 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $39357 r0 *1 796.26,133.28
X$39357 29 1813 1751 1812 1850 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $39358 r0 *1 799.94,133.28
X$39358 48 1597 1598 1852 1851 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $39362 r0 *1 801.78,133.28
X$39362 48 1679 1642 1792 48 29 1733 29 sky130_fd_sc_hd__o21ai_1
* cell instance $39363 r0 *1 803.62,133.28
X$39363 29 1814 1645 1753 1644 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $39364 r0 *1 811.9,133.28
X$39364 48 1644 1814 1815 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $39369 r0 *1 816.96,133.28
X$39369 48 1794 1558 1855 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $39372 r0 *1 819.72,133.28
X$39372 29 1881 1558 1758 1450 1856 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $39374 r0 *1 823.4,133.28
X$39374 48 1704 1352 1487 29 48 1780 29 sky130_fd_sc_hd__a21oi_1
* cell instance $39376 r0 *1 826.16,133.28
X$39376 48 1780 1708 1857 1816 1776 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $39377 r0 *1 828.46,133.28
X$39377 48 1857 1816 1817 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $39382 r0 *1 831.68,133.28
X$39382 48 1489 1759 1505 29 48 1858 29 sky130_fd_sc_hd__a21oi_1
* cell instance $39383 r0 *1 833.52,133.28
X$39383 48 1858 1817 1820 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $39384 r0 *1 836.74,133.28
X$39384 48 1879 1710 1859 1819 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $39386 r0 *1 839.04,133.28
X$39386 29 1860 1566 1818 1324 1819 1762 48 48 29 sky130_fd_sc_hd__o221a_1
* cell instance $39388 r0 *1 843.64,133.28
X$39388 48 1762 1819 1566 29 1986 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $39389 r0 *1 846.86,133.28
X$39389 48 1860 29 1518 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $39392 r0 *1 851,133.28
X$39392 48 1774 1453 1722 29 48 1877 29 sky130_fd_sc_hd__a21oi_1
* cell instance $39394 r0 *1 853.3,133.28
X$39394 29 1721 1566 1877 1648 1765 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $39399 r0 *1 856.98,133.28
X$39399 29 1915 1519 1298 1874 1821 1561 48 48 29 sky130_fd_sc_hd__o32a_1
* cell instance $39400 r0 *1 860.66,133.28
X$39400 29 29 1821 1500 1613 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $39402 r0 *1 863.42,133.28
X$39402 48 1613 1298 1519 48 1862 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $39404 r0 *1 866.64,133.28
X$39404 48 1763 1862 1869 29 48 1717 29 sky130_fd_sc_hd__a21o_1
* cell instance $40052 m0 *1 684.94,138.72
X$40052 48 1865 1128 2002 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40058 m0 *1 692.3,138.72
X$40058 48 1128 1688 1652 1460 890 48 1798 29 29 sky130_fd_sc_hd__o2111ai_1
* cell instance $40059 m0 *1 695.52,138.72
X$40059 48 890 48 29 1836 29 sky130_fd_sc_hd__buf_4
* cell instance $40060 m0 *1 698.28,138.72
X$40060 29 1929 1836 1868 1823 941 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $40062 m0 *1 703.34,138.72
X$40062 48 1619 1512 1888 29 48 1909 29 sky130_fd_sc_hd__a21o_1
* cell instance $40063 m0 *1 706.1,138.72
X$40063 48 1837 1688 1910 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40065 m0 *1 708.4,138.72
X$40065 48 1512 1742 1889 1691 48 1872 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $40066 m0 *1 711.62,138.72
X$40066 48 1512 1889 1691 29 48 1839 29 sky130_fd_sc_hd__a21oi_1
* cell instance $40067 m0 *1 713.46,138.72
X$40067 48 1836 1872 1827 29 48 1911 29 sky130_fd_sc_hd__a21oi_1
* cell instance $40068 m0 *1 715.3,138.72
X$40068 48 1013 1548 1890 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40069 m0 *1 716.68,138.72
X$40069 48 1836 960 1875 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $40072 m0 *1 719.44,138.72
X$40072 29 1892 1839 1552 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $40073 m0 *1 725.42,138.72
X$40073 29 1688 1878 1529 1570 1799 1970 48 48 29 sky130_fd_sc_hd__o221a_2
* cell instance $40075 m0 *1 730.02,138.72
X$40075 48 1552 1512 1745 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $40077 m0 *1 731.86,138.72
X$40077 29 1728 1840 1841 48 2010 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $40078 m0 *1 738.3,138.72
X$40078 29 1777 1842 1830 1318 48 1840 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $40079 m0 *1 742.9,138.72
X$40079 48 1801 1376 1842 1892 1804 48 29 29 sky130_fd_sc_hd__a31o_2
* cell instance $40082 m0 *1 747.04,138.72
X$40082 29 1324 1746 1804 1843 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $40083 m0 *1 753.02,138.72
X$40083 48 1883 1976 1844 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40084 m0 *1 756.24,138.72
X$40084 29 29 1735 48 1802 1803 48 sky130_fd_sc_hd__nor2_2
* cell instance $40085 m0 *1 758.54,138.72
X$40085 29 1844 1287 1747 1805 48 1846 48 29 sky130_fd_sc_hd__nand4_4
* cell instance $40086 m0 *1 766.36,138.72
X$40086 48 1224 1807 1895 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40087 m0 *1 767.74,138.72
X$40087 29 1806 1848 1810 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $40089 m0 *1 772.34,138.72
X$40089 48 1810 1415 1806 48 29 1400 29 sky130_fd_sc_hd__o21ai_1
* cell instance $40091 m0 *1 774.64,138.72
X$40091 29 1886 1834 1642 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $40092 m0 *1 784.76,138.72
X$40092 48 1848 48 29 1695 29 sky130_fd_sc_hd__buf_4
* cell instance $40094 m0 *1 787.98,138.72
X$40094 48 1848 29 1160 48 29 sky130_fd_sc_hd__clkinv_4
* cell instance $40096 m0 *1 791.66,138.72
X$40096 29 1812 1850 1897 1849 1851 1898 48 48 29 sky130_fd_sc_hd__a32oi_4
* cell instance $40098 m0 *1 802.24,138.72
X$40098 48 1751 1795 1853 48 1925 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $40100 m0 *1 804.54,138.72
X$40100 48 1638 1896 1924 1923 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $40102 m0 *1 806.84,138.72
X$40102 48 1638 1701 1957 1854 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $40104 m0 *1 809.14,138.72
X$40104 48 1854 1794 1815 48 29 1901 29 sky130_fd_sc_hd__o21ai_1
* cell instance $40106 m0 *1 811.44,138.72
X$40106 48 1644 1813 1900 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $40107 m0 *1 813.74,138.72
X$40107 48 1601 1673 1855 29 48 1922 29 sky130_fd_sc_hd__a21o_1
* cell instance $40108 m0 *1 816.5,138.72
X$40108 48 1855 1601 1673 29 48 1885 29 sky130_fd_sc_hd__a21oi_1
* cell instance $40109 m0 *1 818.34,138.72
X$40109 29 1884 1703 1885 1856 1901 1831 48 48 29 sky130_fd_sc_hd__o32a_1
* cell instance $40110 m0 *1 822.02,138.72
X$40110 48 1856 1885 1293 29 48 1816 29 sky130_fd_sc_hd__a21oi_1
* cell instance $40112 m0 *1 824.32,138.72
X$40112 48 1922 1902 1537 1857 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $40114 m0 *1 828,138.72
X$40114 48 1816 1857 1879 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40119 m0 *1 833.06,138.72
X$40119 48 1709 1505 1759 1383 29 48 1859 29 sky130_fd_sc_hd__a31oi_1
* cell instance $40120 m0 *1 835.36,138.72
X$40120 29 2203 1422 1818 1504 1828 1919 48 48 29 sky130_fd_sc_hd__a2111oi_4
* cell instance $40121 m0 *1 845.48,138.72
X$40121 48 1422 1571 1860 1572 1861 48 29 29 sky130_fd_sc_hd__or4_1
* cell instance $40123 m0 *1 848.7,138.72
X$40123 48 1861 48 29 1453 29 sky130_fd_sc_hd__buf_4
* cell instance $40126 m0 *1 853.76,138.72
X$40126 48 1763 48 29 1825 29 sky130_fd_sc_hd__inv_1
* cell instance $40127 m0 *1 855.14,138.72
X$40127 48 1766 1763 1771 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40130 m0 *1 857.44,138.72
X$40130 29 1915 1715 1873 1914 1500 1772 48 48 29 sky130_fd_sc_hd__o221ai_2
* cell instance $40131 m0 *1 862.96,138.72
X$40131 29 1191 1561 1821 1613 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $40132 m0 *1 868.94,138.72
X$40132 29 1767 1191 1867 1862 1863 1908 48 48 29 sky130_fd_sc_hd__o311a_1
* cell instance $40710 r0 *1 687.24,138.72
X$40710 29 1652 1944 1769 941 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $40711 r0 *1 689.54,138.72
X$40711 48 1769 1652 941 48 1927 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $40715 r0 *1 695.52,138.72
X$40715 48 1691 1798 1945 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $40716 r0 *1 697.82,138.72
X$40716 29 1887 1889 1826 1660 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $40717 r0 *1 701.5,138.72
X$40717 48 1742 1512 1888 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40719 r0 *1 703.34,138.72
X$40719 48 1836 960 1946 1947 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $40721 r0 *1 705.64,138.72
X$40721 29 1871 1910 960 1930 937 1909 48 48 29 sky130_fd_sc_hd__a32oi_4
* cell instance $40722 r0 *1 715.76,138.72
X$40722 48 1890 1912 1876 1728 29 48 1913 29 sky130_fd_sc_hd__and4_1
* cell instance $40723 r0 *1 718.98,138.72
X$40723 29 1891 1911 1953 1836 1784 1512 48 48 29 sky130_fd_sc_hd__a221oi_4
* cell instance $40726 r0 *1 729.56,138.72
X$40726 48 1916 1318 1933 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40728 r0 *1 733.24,138.72
X$40728 48 1956 960 1880 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40729 r0 *1 736.46,138.72
X$40729 29 2013 1892 1842 1140 1801 1692 48 48 29 sky130_fd_sc_hd__a311o_2
* cell instance $40730 r0 *1 740.6,138.72
X$40730 29 1892 1692 1842 1376 1937 1801 48 48 29 sky130_fd_sc_hd__a311oi_4
* cell instance $40732 r0 *1 750.26,138.72
X$40732 48 1804 1843 1959 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $40733 r0 *1 751.64,138.72
X$40733 48 1918 1376 1694 1735 48 1917 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $40734 r0 *1 753.94,138.72
X$40734 48 1959 1920 1962 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40735 r0 *1 757.16,138.72
X$40735 29 1847 1747 1805 1287 1844 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $40737 r0 *1 760.84,138.72
X$40737 29 1939 1893 1833 1847 1846 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $40738 r0 *1 765.44,138.72
X$40738 48 1894 1939 1895 48 1964 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $40739 r0 *1 767.28,138.72
X$40739 29 1939 1895 1965 1894 1810 1806 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $40742 r0 *1 777.86,138.72
X$40742 29 1695 1042 1896 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $40744 r0 *1 788.44,138.72
X$40744 48 1737 1896 1963 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $40745 r0 *1 789.82,138.72
X$40745 29 1737 1750 1897 1795 1853 1697 48 48 29 sky130_fd_sc_hd__o2111ai_4
* cell instance $40746 r0 *1 799.48,138.72
X$40746 29 1926 1924 1899 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $40748 r0 *1 809.6,138.72
X$40748 48 1701 1644 48 29 29 sky130_fd_sc_hd__clkinv_2
* cell instance $40750 r0 *1 812.36,138.72
X$40750 48 1900 1899 48 1856 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $40752 r0 *1 816.04,138.72
X$40752 48 1601 1673 1901 29 48 1955 29 sky130_fd_sc_hd__a21o_1
* cell instance $40754 r0 *1 820.64,138.72
X$40754 29 1884 1921 1537 1621 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $40755 r0 *1 824.32,138.72
X$40755 29 1903 1325 1902 1703 1952 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $40758 r0 *1 830.76,138.72
X$40758 29 1950 1903 1505 1759 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $40761 r0 *1 838.12,138.72
X$40761 48 1879 1710 1859 1919 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $40767 r0 *1 849.16,138.72
X$40767 48 1518 1948 1263 1905 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $40768 r0 *1 851.46,138.72
X$40768 48 1905 1904 1908 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $40770 r0 *1 855.6,138.72
X$40770 48 1766 1763 1906 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $40773 r0 *1 858.36,138.72
X$40773 48 1613 1773 1906 1914 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $40774 r0 *1 860.2,138.72
X$40774 48 1906 1500 1991 29 48 1907 29 sky130_fd_sc_hd__a21oi_1
* cell instance $40775 r0 *1 862.04,138.72
X$40775 48 1500 1766 1824 1907 48 29 1990 29 sky130_fd_sc_hd__o31ai_1
* cell instance $40776 r0 *1 864.8,138.72
X$40776 48 1771 48 29 1867 29 sky130_fd_sc_hd__inv_1
* cell instance $40777 r0 *1 866.18,138.72
X$40777 48 1763 1191 1862 1869 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $40778 r0 *1 868.02,138.72
X$40778 48 1191 1867 1862 1908 48 29 1822 29 sky130_fd_sc_hd__o31ai_1
* cell instance $41416 m0 *1 692.3,144.16
X$41416 29 1989 1928 1927 1944 1929 1889 48 48 29 sky130_fd_sc_hd__a2111oi_1
* cell instance $41420 m0 *1 696.44,144.16
X$41420 48 1826 1887 2003 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $41422 m0 *1 699.2,144.16
X$41422 48 1929 2030 1993 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $41424 m0 *1 701.5,144.16
X$41424 48 1888 1619 1946 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $41426 m0 *1 705.64,144.16
X$41426 48 1512 1619 1994 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $41427 m0 *1 708.86,144.16
X$41427 29 1891 1839 1512 1913 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $41428 m0 *1 713,144.16
X$41428 48 980 1931 1932 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $41429 m0 *1 714.38,144.16
X$41429 29 1890 1912 1876 1728 48 1949 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $41431 m0 *1 719.44,144.16
X$41431 29 29 1876 1954 1728 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $41434 m0 *1 721.74,144.16
X$41434 48 1784 1912 2034 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $41435 m0 *1 723.12,144.16
X$41435 29 1800 1548 1934 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $41436 m0 *1 733.24,144.16
X$41436 29 1971 1933 1934 1185 48 2126 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $41437 m0 *1 737.84,144.16
X$41437 29 1781 1935 1997 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $41438 m0 *1 743.82,144.16
X$41438 29 29 1666 1842 1512 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $41441 m0 *1 747.04,144.16
X$41441 48 1880 1376 1041 1692 29 2014 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $41444 m0 *1 749.8,144.16
X$41444 48 1973 1938 2127 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $41445 m0 *1 751.18,144.16
X$41445 29 1832 1998 1694 1936 48 1961 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $41446 m0 *1 759,144.16
X$41446 29 29 1975 48 1139 1976 48 sky130_fd_sc_hd__nor2_2
* cell instance $41447 m0 *1 761.3,144.16
X$41447 29 29 1936 48 1224 1976 48 sky130_fd_sc_hd__nor2_2
* cell instance $41449 m0 *1 764.06,144.16
X$41449 29 1894 1893 1833 1846 1847 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $41450 m0 *1 767.74,144.16
X$41450 29 1978 1847 1846 1977 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $41452 m0 *1 772.34,144.16
X$41452 48 1940 1638 1979 29 48 1966 29 sky130_fd_sc_hd__a21oi_1
* cell instance $41456 m0 *1 774.64,144.16
X$41456 29 1941 1980 2001 1999 1965 1964 48 48 29 sky130_fd_sc_hd__a32o_2
* cell instance $41457 m0 *1 778.78,144.16
X$41457 29 2001 1980 1795 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $41458 m0 *1 788.9,144.16
X$41458 48 1638 1852 2000 1940 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $41459 m0 *1 790.74,144.16
X$41459 29 1698 1960 1795 1749 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $41461 m0 *1 793.96,144.16
X$41461 48 1697 1750 1982 29 1898 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $41462 m0 *1 797.18,144.16
X$41462 48 1697 1750 1737 29 1926 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $41468 m0 *1 802.24,144.16
X$41468 48 1119 1925 1923 29 48 1958 29 sky130_fd_sc_hd__a21oi_1
* cell instance $41470 m0 *1 804.54,144.16
X$41470 48 1899 1813 1957 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $41471 m0 *1 807.76,144.16
X$41471 48 1638 1899 1814 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $41472 m0 *1 809.14,144.16
X$41472 48 1644 48 29 1118 29 sky130_fd_sc_hd__buf_4
* cell instance $41474 m0 *1 812.82,144.16
X$41474 29 1902 1900 1899 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $41476 m0 *1 819.72,144.16
X$41476 48 1902 1922 1942 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $41477 m0 *1 822.94,144.16
X$41477 48 1996 1995 1942 29 48 1951 29 sky130_fd_sc_hd__a21oi_1
* cell instance $41479 m0 *1 825.24,144.16
X$41479 48 1325 1621 1995 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $41480 m0 *1 826.62,144.16
X$41480 48 1884 1325 1952 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $41488 m0 *1 832.6,144.16
X$41488 48 1383 29 1489 48 29 sky130_fd_sc_hd__buf_2
* cell instance $41493 m0 *1 845.94,144.16
X$41493 48 1571 1422 1987 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $41496 m0 *1 853.76,144.16
X$41496 48 1763 1943 1766 1988 29 1773 48 29 sky130_fd_sc_hd__nor4b_1
* cell instance $41500 m0 *1 857.44,144.16
X$41500 48 1763 1766 1874 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $41501 m0 *1 859.74,144.16
X$41501 48 1992 29 1561 48 29 sky130_fd_sc_hd__buf_2
* cell instance $41504 m0 *1 863.88,144.16
X$41504 48 1863 2143 1990 1864 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $42146 r0 *1 689.08,144.16
X$42146 29 1944 1968 1927 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $42149 r0 *1 693.68,144.16
X$42149 29 2029 1967 2028 1913 48 48 29 sky130_fd_sc_hd__mux2i_1
* cell instance $42150 r0 *1 697.36,144.16
X$42150 48 1836 1969 1967 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $42151 r0 *1 698.74,144.16
X$42151 29 29 1969 48 1887 1826 48 sky130_fd_sc_hd__nor2_2
* cell instance $42153 r0 *1 701.96,144.16
X$42153 48 1870 1913 2032 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $42156 r0 *1 705.64,144.16
X$42156 48 1994 1949 2004 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $42157 r0 *1 708.86,144.16
X$42157 29 1953 1619 2300 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $42158 r0 *1 718.98,144.16
X$42158 48 1912 48 29 1931 29 sky130_fd_sc_hd__inv_1
* cell instance $42160 r0 *1 720.36,144.16
X$42160 29 2109 1875 1836 2034 2036 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $42161 r0 *1 727.72,144.16
X$42161 48 980 1934 2037 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $42163 r0 *1 730.48,144.16
X$42163 48 1468 1970 2012 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $42165 r0 *1 733.24,144.16
X$42165 29 1971 1935 1781 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $42166 r0 *1 739.22,144.16
X$42166 29 29 1840 1976 1841 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $42167 r0 *1 741.52,144.16
X$42167 29 1938 696 1624 1974 1969 2016 48 48 29 sky130_fd_sc_hd__a41oi_4
* cell instance $42169 r0 *1 751.64,144.16
X$42169 48 1843 1090 48 29 29 sky130_fd_sc_hd__inv_6
* cell instance $42170 r0 *1 754.86,144.16
X$42170 48 1515 1692 1962 1883 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42171 r0 *1 756.7,144.16
X$42171 48 1735 1670 1785 29 48 1920 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42172 r0 *1 758.54,144.16
X$42172 48 1108 1976 2044 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42175 r0 *1 760.84,144.16
X$42175 29 1747 1031 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $42176 r0 *1 764.98,144.16
X$42176 48 1893 1833 2046 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42178 r0 *1 766.82,144.16
X$42178 29 1846 2078 1847 1977 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $42179 r0 *1 769.12,144.16
X$42179 29 2001 1978 1809 1808 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $42181 r0 *1 775.1,144.16
X$42181 48 1980 2053 1999 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42184 r0 *1 777.86,144.16
X$42184 29 2001 2017 1924 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $42186 r0 *1 788.44,144.16
X$42186 29 2077 1981 2047 2019 1679 1398 48 48 29 sky130_fd_sc_hd__o311ai_1
* cell instance $42187 r0 *1 791.66,144.16
X$42187 48 1896 1795 1852 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42189 r0 *1 793.5,144.16
X$42189 48 1966 1484 1896 29 48 2020 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42190 r0 *1 795.34,144.16
X$42190 48 1737 1853 1795 1982 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42191 r0 *1 797.18,144.16
X$42191 48 1851 1897 1898 1983 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $42193 r0 *1 799.94,144.16
X$42193 48 1679 1737 1751 1896 29 2042 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $42195 r0 *1 802.24,144.16
X$42195 48 2020 2042 2040 1958 29 2041 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $42198 r0 *1 805.92,144.16
X$42198 48 1701 29 1416 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $42200 r0 *1 809.6,144.16
X$42200 48 2088 1813 1983 29 48 2039 29 sky130_fd_sc_hd__a21boi_0
* cell instance $42201 r0 *1 812.36,144.16
X$42201 48 1416 1813 1983 29 48 2184 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42208 r0 *1 822.02,144.16
X$42208 48 1158 1881 1996 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42209 r0 *1 823.4,144.16
X$42209 48 1881 1703 2038 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $42211 r0 *1 827.54,144.16
X$42211 48 1537 29 1325 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $42214 r0 *1 831.22,144.16
X$42214 48 1951 2035 2059 48 1985 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $42217 r0 *1 835.82,144.16
X$42217 48 2021 1489 1950 48 29 2023 29 sky130_fd_sc_hd__o21bai_1
* cell instance $42218 r0 *1 838.58,144.16
X$42218 48 1984 2060 1904 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42219 r0 *1 839.96,144.16
X$42219 48 2021 2022 1984 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42220 r0 *1 841.34,144.16
X$42220 48 1489 1950 2022 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42223 r0 *1 843.64,144.16
X$42223 48 1985 1986 2024 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $42224 r0 *1 846.86,144.16
X$42224 48 2024 1572 1987 29 48 1766 29 sky130_fd_sc_hd__o21a_2
* cell instance $42225 r0 *1 850.08,144.16
X$42225 48 1518 1948 2061 2026 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42226 r0 *1 851.92,144.16
X$42226 48 2033 1453 2026 29 48 1988 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42228 r0 *1 854.68,144.16
X$42228 48 2031 1988 2025 1766 29 48 2027 29 sky130_fd_sc_hd__a31oi_1
* cell instance $42230 r0 *1 856.98,144.16
X$42230 29 1988 1992 1763 1766 48 48 1943 29 sky130_fd_sc_hd__or4b_1
* cell instance $42232 r0 *1 861.12,144.16
X$42232 48 1763 2027 1991 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42869 m0 *1 686.78,149.6
X$42869 48 1928 2098 2029 48 29 2048 29 sky130_fd_sc_hd__o21bai_1
* cell instance $42870 m0 *1 689.54,149.6
X$42870 48 2003 1928 1870 2062 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42872 m0 *1 691.84,149.6
X$42872 48 1989 1945 2002 48 29 2063 29 sky130_fd_sc_hd__o21ai_1
* cell instance $42875 m0 *1 693.68,149.6
X$42875 48 1836 2003 1870 2028 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $42876 m0 *1 695.52,149.6
X$42876 48 1929 1889 1928 29 48 2099 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42878 m0 *1 697.82,149.6
X$42878 48 1928 1660 1969 29 48 2030 29 sky130_fd_sc_hd__a21boi_0
* cell instance $42879 m0 *1 700.58,149.6
X$42879 48 937 1928 2065 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42881 m0 *1 702.42,149.6
X$42881 29 2004 960 1836 2049 1947 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $42883 m0 *1 710.7,149.6
X$42883 29 29 1969 1972 1660 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $42885 m0 *1 713.46,149.6
X$42885 29 29 1912 2005 980 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $42887 m0 *1 716.68,149.6
X$42887 48 1934 1954 1784 2005 29 2080 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $42889 m0 *1 719.44,149.6
X$42889 29 2006 2005 1932 48 2007 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $42892 m0 *1 724.5,149.6
X$42892 29 2008 2006 1912 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $42893 m0 *1 730.48,149.6
X$42893 48 2009 2036 2066 2011 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $42894 m0 *1 732.32,149.6
X$42894 48 1692 2010 1804 2007 29 48 2068 29 sky130_fd_sc_hd__or4b_2
* cell instance $42895 m0 *1 736,149.6
X$42895 48 2010 2013 2008 2179 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $42896 m0 *1 738.3,149.6
X$42896 29 2072 1108 1976 1997 2014 48 48 29 sky130_fd_sc_hd__nor4b_2
* cell instance $42897 m0 *1 743.82,149.6
X$42897 48 1529 2043 2016 2052 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $42900 m0 *1 747.04,149.6
X$42900 48 1972 48 29 1973 29 sky130_fd_sc_hd__inv_1
* cell instance $42904 m0 *1 748.88,149.6
X$42904 48 2015 2050 2051 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42905 m0 *1 750.26,149.6
X$42905 48 2073 1918 1735 1998 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42906 m0 *1 752.1,149.6
X$42906 48 1785 2051 2075 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $42907 m0 *1 753.48,149.6
X$42907 29 1970 2076 2045 1974 2043 2212 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $42908 m0 *1 763.14,149.6
X$42908 48 1674 29 1747 48 29 sky130_fd_sc_hd__clkinv_4
* cell instance $42910 m0 *1 768.2,149.6
X$42910 48 2078 29 2053 48 29 sky130_fd_sc_hd__buf_2
* cell instance $42912 m0 *1 770.96,149.6
X$42912 48 1848 1978 2017 48 2018 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $42920 m0 *1 776.02,149.6
X$42920 48 1980 2053 2122 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $42922 m0 *1 778.32,149.6
X$42922 29 1848 2054 1853 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $42923 m0 *1 788.44,149.6
X$42923 48 1324 2118 2077 29 48 1516 29 sky130_fd_sc_hd__a21oi_1
* cell instance $42924 m0 *1 790.28,149.6
X$42924 48 1853 1924 2000 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $42926 m0 *1 792.12,149.6
X$42926 48 1853 1737 2055 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $42927 m0 *1 794.42,149.6
X$42927 48 1598 1597 1751 1795 29 48 2074 29 sky130_fd_sc_hd__a31oi_1
* cell instance $42928 m0 *1 796.72,149.6
X$42928 48 1697 1924 1750 48 29 2057 29 sky130_fd_sc_hd__o21ai_1
* cell instance $42929 m0 *1 798.56,149.6
X$42929 48 2057 1853 2058 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $42933 m0 *1 802.24,149.6
X$42933 48 1751 1896 1795 2071 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42936 m0 *1 806.84,149.6
X$42936 29 2070 1703 2058 1118 48 48 29 sky130_fd_sc_hd__o21bai_4
* cell instance $42937 m0 *1 813.74,149.6
X$42937 29 1813 2069 2040 1983 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $42938 m0 *1 816.04,149.6
X$42938 48 1955 29 2067 48 29 sky130_fd_sc_hd__buf_2
* cell instance $42941 m0 *1 823.4,149.6
X$42941 48 1293 29 1158 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $42942 m0 *1 826.16,149.6
X$42942 48 2097 1703 2059 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $42948 m0 *1 832.6,149.6
X$42948 48 1383 1951 2059 2035 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $42950 m0 *1 836.28,149.6
X$42950 48 1950 1383 2021 2060 29 48 29 sky130_fd_sc_hd__nor3b_1
* cell instance $42951 m0 *1 839.04,149.6
X$42951 29 2023 1572 2060 1985 2025 48 48 29 sky130_fd_sc_hd__nand4b_4
* cell instance $42952 m0 *1 847.78,149.6
X$42952 48 1985 48 29 1948 29 sky130_fd_sc_hd__inv_1
* cell instance $42953 m0 *1 849.16,149.6
X$42953 48 2061 1948 1518 48 2033 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $42954 m0 *1 851.92,149.6
X$42954 48 1518 1986 2064 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $42955 m0 *1 854.22,149.6
X$42955 48 2025 2031 1943 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $43656 r0 *1 689.54,149.6
X$43656 48 2003 1870 2098 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43658 r0 *1 691.38,149.6
X$43658 48 1945 2002 1989 48 2101 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $43663 r0 *1 694.6,149.6
X$43663 48 2099 1870 1913 48 29 2100 29 sky130_fd_sc_hd__a21bo_2
* cell instance $43664 r0 *1 698.28,149.6
X$43664 29 2217 1949 1929 2030 2062 2065 48 48 29 sky130_fd_sc_hd__a2111o_1
* cell instance $43666 r0 *1 702.88,149.6
X$43666 29 29 2081 48 1945 2032 48 sky130_fd_sc_hd__nor2_2
* cell instance $43668 r0 *1 705.64,149.6
X$43668 48 1468 2048 1993 48 29 2102 29 sky130_fd_sc_hd__a21boi_1
* cell instance $43669 r0 *1 708.4,149.6
X$43669 29 1784 937 2249 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $43670 r0 *1 718.52,149.6
X$43670 48 2080 2106 2079 2107 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $43674 r0 *1 720.82,149.6
X$43674 29 29 2006 48 1784 1954 48 sky130_fd_sc_hd__nor2_2
* cell instance $43676 r0 *1 723.58,149.6
X$43676 29 1784 2125 1954 2005 48 48 29 sky130_fd_sc_hd__nor3_4
* cell instance $43677 r0 *1 729.56,149.6
X$43677 48 1931 1954 2109 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $43679 r0 *1 733.24,149.6
X$43679 48 2006 1931 2112 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $43680 r0 *1 736.46,149.6
X$43680 29 29 2009 48 2010 2013 48 sky130_fd_sc_hd__nor2_2
* cell instance $43681 r0 *1 738.76,149.6
X$43681 48 2010 2013 2008 48 2114 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $43682 r0 *1 740.6,149.6
X$43682 48 1936 1937 2115 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $43684 r0 *1 742.9,149.6
X$43684 48 2012 2081 2016 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $43685 r0 *1 745.2,149.6
X$43685 48 2015 2052 2082 2116 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $43686 r0 *1 747.04,149.6
X$43686 48 2015 2082 2150 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43690 r0 *1 748.42,149.6
X$43690 48 1973 2043 1146 2156 2150 2083 29 48 29 sky130_fd_sc_hd__a311o_1
* cell instance $43692 r0 *1 752.56,149.6
X$43692 29 2081 2085 640 2043 1970 48 48 29 sky130_fd_sc_hd__nor4_4
* cell instance $43694 r0 *1 760.84,149.6
X$43694 48 1936 2014 2119 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $43696 r0 *1 763.14,149.6
X$43696 48 2151 2075 2120 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $43697 r0 *1 765.44,149.6
X$43697 29 29 2094 48 2052 2045 48 sky130_fd_sc_hd__nor2_2
* cell instance $43699 r0 *1 768.66,149.6
X$43699 48 1445 48 29 2054 29 sky130_fd_sc_hd__buf_4
* cell instance $43700 r0 *1 771.42,149.6
X$43700 48 1695 2121 2131 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43701 r0 *1 772.8,149.6
X$43701 48 1848 2122 2134 2123 48 2084 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $43706 r0 *1 776.48,149.6
X$43706 48 1695 2122 1941 29 48 2124 29 sky130_fd_sc_hd__a21oi_1
* cell instance $43708 r0 *1 778.78,149.6
X$43708 29 2047 2018 2084 1642 1417 48 48 29 sky130_fd_sc_hd__a211o_2
* cell instance $43710 r0 *1 782.92,149.6
X$43710 48 1981 2047 2055 1963 48 29 1979 29 sky130_fd_sc_hd__o31ai_1
* cell instance $43712 r0 *1 786.6,149.6
X$43712 48 1981 2047 2086 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43714 r0 *1 788.44,149.6
X$43714 29 2118 1417 1750 2117 2019 2086 48 48 29 sky130_fd_sc_hd__o41ai_1
* cell instance $43717 r0 *1 793.04,149.6
X$43717 48 1751 2087 2055 29 48 2056 29 sky130_fd_sc_hd__a21oi_1
* cell instance $43719 r0 *1 795.34,149.6
X$43719 48 1982 1941 1853 29 48 2113 29 sky130_fd_sc_hd__a21oi_1
* cell instance $43720 r0 *1 797.18,149.6
X$43720 29 2111 2074 2057 1896 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $43721 r0 *1 801.32,149.6
X$43721 48 2110 2088 2111 2056 48 2070 29 29 sky130_fd_sc_hd__o2bb2ai_1
* cell instance $43726 r0 *1 805,149.6
X$43726 29 2108 2162 2040 1701 2088 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $43727 r0 *1 812.82,149.6
X$43727 48 2105 29 1731 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $43732 r0 *1 819.26,149.6
X$43732 48 2140 2104 2103 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43735 r0 *1 823.4,149.6
X$43735 48 1537 29 48 1293 29 sky130_fd_sc_hd__inv_2
* cell instance $43736 r0 *1 824.78,149.6
X$43736 29 1703 2096 2067 1293 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $43737 r0 *1 827.08,149.6
X$43737 48 1788 1158 2097 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $43738 r0 *1 828.46,149.6
X$43738 48 1325 2038 2089 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $43744 r0 *1 832.6,149.6
X$43744 29 2089 1240 2095 1921 2021 48 48 29 sky130_fd_sc_hd__and4b_1
* cell instance $43747 r0 *1 839.04,149.6
X$43747 48 2022 2021 2061 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $43751 r0 *1 845.48,149.6
X$43751 48 1518 1572 2093 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $43752 r0 *1 846.86,149.6
X$43752 48 1904 1985 1986 2025 29 48 2174 29 sky130_fd_sc_hd__a31oi_1
* cell instance $43753 r0 *1 849.16,149.6
X$43753 48 1572 48 29 2092 29 sky130_fd_sc_hd__inv_1
* cell instance $43754 r0 *1 850.54,149.6
X$43754 48 1987 2092 2064 2091 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $43755 r0 *1 852.38,149.6
X$43755 48 1986 1518 2031 2090 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $44413 m0 *1 695.52,155.04
X$44413 29 2100 1968 2144 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $44414 m0 *1 705.64,155.04
X$44414 48 1784 1836 2079 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $44415 m0 *1 708.86,155.04
X$44415 48 1784 1954 1931 48 2155 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $44417 m0 *1 711.16,155.04
X$44417 29 2101 2102 1972 2204 48 2082 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $44419 m0 *1 719.44,155.04
X$44419 48 2080 2049 2106 48 29 2176 29 sky130_fd_sc_hd__or3_2
* cell instance $44420 m0 *1 722.2,155.04
X$44420 29 1934 2125 2145 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $44421 m0 *1 728.18,155.04
X$44421 29 2010 2013 2037 2036 48 2220 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $44422 m0 *1 736,155.04
X$44422 48 2037 2036 2013 2010 48 29 2148 29 sky130_fd_sc_hd__o211a_2
* cell instance $44423 m0 *1 739.68,155.04
X$44423 48 2179 2189 2114 2072 48 2243 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $44424 m0 *1 741.98,155.04
X$44424 29 2050 1529 2043 2016 2082 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $44426 m0 *1 747.04,155.04
X$44426 29 2050 2073 2015 48 48 29 sky130_fd_sc_hd__nand2b_4
* cell instance $44428 m0 *1 753.02,155.04
X$44428 48 2075 2127 640 48 2129 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $44429 m0 *1 755.78,155.04
X$44429 48 640 2127 2151 29 48 2152 29 sky130_fd_sc_hd__a21oi_1
* cell instance $44431 m0 *1 758.08,155.04
X$44431 29 1674 2128 2129 2130 48 2153 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $44432 m0 *1 765.9,155.04
X$44432 48 2130 1160 2132 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $44434 m0 *1 768.2,155.04
X$44434 29 2133 2120 2158 2085 2132 2121 48 48 29 sky130_fd_sc_hd__o2111a_1
* cell instance $44435 m0 *1 772.34,155.04
X$44435 48 2134 2131 2135 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $44438 m0 *1 774.64,155.04
X$44438 48 1808 1809 2053 2159 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $44440 m0 *1 776.94,155.04
X$44440 29 2187 1695 2054 2124 1941 48 48 29 sky130_fd_sc_hd__a2bb2oi_1
* cell instance $44442 m0 *1 780.62,155.04
X$44442 29 1981 2047 2133 2136 48 1699 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $44444 m0 *1 788.9,155.04
X$44444 48 2133 2136 2047 1981 48 29 1597 29 sky130_fd_sc_hd__o211a_2
* cell instance $44446 m0 *1 793.04,155.04
X$44446 48 1697 1750 1941 48 2087 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $44449 m0 *1 796.26,155.04
X$44449 48 1751 2113 2137 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $44450 m0 *1 797.64,155.04
X$44450 29 2110 2071 2137 1484 48 48 29 sky130_fd_sc_hd__mux2_1
* cell instance $44452 m0 *1 802.24,155.04
X$44452 29 2137 2108 2071 1484 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $44453 m0 *1 810.52,155.04
X$44453 29 2039 2070 2105 2154 2041 2069 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $44454 m0 *1 814.2,155.04
X$44454 29 29 2138 2140 2139 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $44455 m0 *1 816.5,155.04
X$44455 29 2139 2067 2182 2104 2138 1703 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $44457 m0 *1 823.86,155.04
X$44457 48 2140 1788 48 2149 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $44461 m0 *1 829.84,155.04
X$44461 29 2021 2096 2104 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $44462 m0 *1 835.82,155.04
X$44462 48 2147 2141 2095 48 2025 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $44463 m0 *1 838.58,155.04
X$44463 48 2178 2146 1866 2273 48 2142 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $44465 m0 *1 841.8,155.04
X$44465 29 2143 2142 2085 2172 1987 2093 48 48 29 sky130_fd_sc_hd__a41oi_2
* cell instance $44467 m0 *1 849.62,155.04
X$44467 48 2031 2091 2090 2092 1987 2169 29 48 29 sky130_fd_sc_hd__a32oi_1
* cell instance $45109 r0 *1 695.06,155.04
X$45109 29 1968 2100 2219 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $45111 r0 *1 705.64,155.04
X$45111 29 1546 1930 2218 48 48 29 sky130_fd_sc_hd__xor2_2
* cell instance $45112 r0 *1 711.62,155.04
X$45112 48 2171 2188 2144 48 2170 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $45113 r0 *1 714.84,155.04
X$45113 48 1934 980 2155 48 29 2106 29 sky130_fd_sc_hd__a21boi_1
* cell instance $45115 r0 *1 718.06,155.04
X$45115 29 2125 1934 2066 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $45120 r0 *1 728.64,155.04
X$45120 29 2206 2191 2126 2008 2013 1013 48 48 29 sky130_fd_sc_hd__o41a_1
* cell instance $45122 r0 *1 733.24,155.04
X$45122 29 2126 2043 2148 2176 2207 48 48 29 sky130_fd_sc_hd__nor4_4
* cell instance $45123 r0 *1 741.06,155.04
X$45123 29 1090 2115 2119 48 2208 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $45124 r0 *1 746.12,155.04
X$45124 48 2183 2209 2156 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $45128 r0 *1 748.42,155.04
X$45128 29 1938 2150 2156 1146 2043 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $45129 r0 *1 751.64,155.04
X$45129 29 2157 2183 1918 1670 2052 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $45130 r0 *1 754.86,155.04
X$45130 48 2076 2157 29 48 1307 29 sky130_fd_sc_hd__nor2b_2
* cell instance $45131 r0 *1 758.08,155.04
X$45131 48 1031 2128 2151 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $45133 r0 *1 760.84,155.04
X$45133 29 2085 2132 2117 2120 2158 2121 48 48 29 sky130_fd_sc_hd__o2111ai_4
* cell instance $45134 r0 *1 770.5,155.04
X$45134 48 2120 2132 2121 48 2194 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $45135 r0 *1 773.26,155.04
X$45135 29 2215 2186 1965 2159 2228 2214 48 48 29 sky130_fd_sc_hd__a221oi_2
* cell instance $45139 r0 *1 778.78,155.04
X$45139 48 2159 1965 2213 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $45142 r0 *1 783.38,155.04
X$45142 29 1981 2185 2160 1310 2230 48 48 29 sky130_fd_sc_hd__a211o_2
* cell instance $45146 r0 *1 789.36,155.04
X$45146 29 2195 2196 1679 2019 2117 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $45148 r0 *1 797.64,155.04
X$45148 29 2147 2086 2136 1679 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $45154 r0 *1 804.08,155.04
X$45154 29 2161 2154 2162 2058 2088 2108 48 48 29 sky130_fd_sc_hd__a2111oi_0
* cell instance $45156 r0 *1 807.76,155.04
X$45156 48 2161 2162 2110 48 29 2138 29 sky130_fd_sc_hd__o21ai_1
* cell instance $45157 r0 *1 809.6,155.04
X$45157 29 2104 2184 2161 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $45159 r0 *1 816.04,155.04
X$45159 48 1702 2163 2198 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $45161 r0 *1 817.88,155.04
X$45161 48 2163 2067 1731 48 29 1487 29 sky130_fd_sc_hd__a21bo_2
* cell instance $45162 r0 *1 821.56,155.04
X$45162 48 2180 1293 2164 2182 2181 48 29 29 sky130_fd_sc_hd__a31o_2
* cell instance $45163 r0 *1 824.78,155.04
X$45163 48 2067 1731 2149 2164 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $45169 r0 *1 832.14,155.04
X$45169 48 2165 2140 48 2141 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $45170 r0 *1 835.36,155.04
X$45170 48 2140 2165 1866 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $45172 r0 *1 837.66,155.04
X$45172 48 2166 2168 2167 2201 29 2177 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $45174 r0 *1 840.42,155.04
X$45174 48 2181 1950 2241 2202 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $45177 r0 *1 843.64,155.04
X$45177 48 2175 48 29 2172 29 sky130_fd_sc_hd__inv_1
* cell instance $45179 r0 *1 845.48,155.04
X$45179 29 1863 2173 2168 2174 2169 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $45841 m0 *1 697.82,160.48
X$45841 29 29 2217 2188 2063 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $45842 m0 *1 700.12,160.48
X$45842 48 2063 2217 48 2191 29 29 sky130_fd_sc_hd__and2_2
* cell instance $45844 m0 *1 703.8,160.48
X$45844 29 1930 1546 2171 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $45845 m0 *1 713.92,160.48
X$45845 29 2049 2248 2080 2106 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $45846 m0 *1 717.6,160.48
X$45846 48 2066 2079 2189 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $45848 m0 *1 719.44,160.48
X$45848 29 2144 2204 2171 2101 2145 2049 48 48 29 sky130_fd_sc_hd__o2111ai_2
* cell instance $45850 m0 *1 725.42,160.48
X$45850 29 2190 2148 2144 2171 2176 48 48 29 sky130_fd_sc_hd__o211ai_2
* cell instance $45851 m0 *1 730.02,160.48
X$45851 29 2190 2191 2222 2115 1971 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $45852 m0 *1 737.38,160.48
X$45852 29 2011 2183 2243 1090 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $45855 m0 *1 747.04,160.48
X$45855 29 2223 2192 2051 2244 2015 2245 48 48 29 sky130_fd_sc_hd__o32a_1
* cell instance $45856 m0 *1 750.72,160.48
X$45856 48 2192 2051 2183 1785 2245 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $45859 m0 *1 755.32,160.48
X$45859 48 1670 2211 2224 2305 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $45860 m0 *1 757.16,160.48
X$45860 29 2212 2131 2120 2130 2152 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $45862 m0 *1 762.68,160.48
X$45862 48 2012 2153 2134 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $45863 m0 *1 764.06,160.48
X$45863 48 2130 2153 2246 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $45864 m0 *1 765.44,160.48
X$45864 29 2158 2130 2246 2226 48 48 29 sky130_fd_sc_hd__mux2_2
* cell instance $45866 m0 *1 770.5,160.48
X$45866 48 2017 2216 1978 48 29 2214 29 sky130_fd_sc_hd__o21ai_1
* cell instance $45868 m0 *1 772.8,160.48
X$45868 48 2153 48 29 2227 29 sky130_fd_sc_hd__inv_1
* cell instance $45871 m0 *1 775.1,160.48
X$45871 48 2193 1980 2053 2228 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $45872 m0 *1 776.94,160.48
X$45872 29 29 2231 48 2216 2187 48 sky130_fd_sc_hd__nor2_2
* cell instance $45873 m0 *1 779.24,160.48
X$45873 48 2213 29 1737 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $45874 m0 *1 782,160.48
X$45874 29 2017 1737 2196 2186 2229 48 48 29 sky130_fd_sc_hd__o2bb2ai_2
* cell instance $45875 m0 *1 787.52,160.48
X$45875 48 1737 2160 2185 29 48 2247 29 sky130_fd_sc_hd__a21oi_1
* cell instance $45877 m0 *1 789.82,160.48
X$45877 29 29 2195 1598 2196 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $45878 m0 *1 792.12,160.48
X$45878 48 2195 2196 2210 2019 29 2234 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $45880 m0 *1 795.34,160.48
X$45880 29 2197 2086 1679 2234 2194 48 48 29 sky130_fd_sc_hd__a2bb2oi_2
* cell instance $45884 m0 *1 804.08,160.48
X$45884 29 2147 2236 1307 2135 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $45887 m0 *1 807.76,160.48
X$45887 48 1751 2162 2280 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $45888 m0 *1 809.14,160.48
X$45888 48 2108 2040 2260 2088 48 2139 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $45890 m0 *1 815.12,160.48
X$45890 48 2237 2173 2045 2178 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $45891 m0 *1 816.96,160.48
X$45891 48 1731 2067 2103 2198 29 2180 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $45892 m0 *1 819.72,160.48
X$45892 29 1537 2198 1731 2067 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $45894 m0 *1 826.16,160.48
X$45894 48 2205 1921 2199 2089 29 2238 48 29 sky130_fd_sc_hd__nor4b_1
* cell instance $45897 m0 *1 831.68,160.48
X$45897 48 2173 2240 2200 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $45898 m0 *1 833.06,160.48
X$45898 29 2181 1950 2242 2203 2200 48 48 29 sky130_fd_sc_hd__o31ai_2
* cell instance $45899 m0 *1 837.66,160.48
X$45899 29 2094 1571 2175 2146 2200 48 48 29 sky130_fd_sc_hd__nand4b_4
* cell instance $45900 m0 *1 846.4,160.48
X$45900 48 2202 2201 2031 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $46544 r0 *1 699.2,160.48
X$46544 29 2219 2191 2218 2251 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $46547 r0 *1 706.56,160.48
X$46547 48 2188 2219 2271 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $46549 r0 *1 708.4,160.48
X$46549 29 2066 2270 2007 2079 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $46551 r0 *1 711.16,160.48
X$46551 48 2218 2220 2248 29 48 2272 29 sky130_fd_sc_hd__a21oi_1
* cell instance $46553 r0 *1 713.46,160.48
X$46553 29 2188 2148 2049 2066 2251 48 2274 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $46558 r0 *1 723.58,160.48
X$46558 29 2206 2248 2220 2170 1843 48 48 29 sky130_fd_sc_hd__a31o_4
* cell instance $46560 r0 *1 730.48,160.48
X$46560 48 1937 2171 2144 2007 48 2207 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $46562 r0 *1 733.24,160.48
X$46562 29 1997 1936 2251 2221 1937 2250 48 48 29 sky130_fd_sc_hd__a41oi_4
* cell instance $46563 r0 *1 743.36,160.48
X$46563 29 29 2276 48 2222 2221 48 sky130_fd_sc_hd__nor2_2
* cell instance $46564 r0 *1 745.66,160.48
X$46564 48 2116 29 1670 48 29 sky130_fd_sc_hd__clkbuf_4
* cell instance $46568 r0 *1 748.42,160.48
X$46568 29 2223 2277 2083 2157 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $46569 r0 *1 752.1,160.48
X$46569 29 2279 2252 2223 2083 2130 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $46572 r0 *1 760.84,160.48
X$46572 48 2211 2224 2244 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $46573 r0 *1 762.22,160.48
X$46573 48 2211 2183 2281 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $46575 r0 *1 764.06,160.48
X$46575 48 2225 2254 2253 48 2123 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $46577 r0 *1 766.36,160.48
X$46577 48 1810 2225 2226 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $46579 r0 *1 768.2,160.48
X$46579 48 2054 1980 2053 29 48 2282 29 sky130_fd_sc_hd__a21oi_1
* cell instance $46580 r0 *1 770.04,160.48
X$46580 48 2017 1978 2255 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $46581 r0 *1 771.42,160.48
X$46581 29 2216 2226 2227 2054 48 2160 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $46585 r0 *1 776.02,160.48
X$46585 29 2227 2226 2229 2054 2216 48 48 29 sky130_fd_sc_hd__and4_2
* cell instance $46586 r0 *1 779.7,160.48
X$46586 29 2257 2213 2017 2229 2186 48 48 29 sky130_fd_sc_hd__a2bb2oi_2
* cell instance $46587 r0 *1 785.22,160.48
X$46587 48 2230 2258 1941 2284 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $46592 r0 *1 792.58,160.48
X$46592 29 2283 2233 2231 2161 2232 1697 48 48 29 sky130_fd_sc_hd__o32ai_4
* cell instance $46596 r0 *1 802.7,160.48
X$46596 48 2040 1849 2235 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $46597 r0 *1 804.08,160.48
X$46597 29 2259 2235 2280 2327 2236 48 2237 48 29 sky130_fd_sc_hd__o311ai_4
* cell instance $46598 r0 *1 813.74,160.48
X$46598 48 2147 2135 2278 2240 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $46601 r0 *1 816.96,160.48
X$46601 48 1702 2237 29 48 2265 29 sky130_fd_sc_hd__nor2b_2
* cell instance $46604 r0 *1 824.78,160.48
X$46604 29 2038 2302 2239 2205 1537 2275 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $46605 r0 *1 828.46,160.48
X$46605 29 2181 1383 2199 1921 2239 48 48 29 sky130_fd_sc_hd__nor4_4
* cell instance $46609 r0 *1 836.28,160.48
X$46609 48 2167 2238 2241 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $46610 r0 *1 838.58,160.48
X$46610 48 2181 1950 2241 2177 48 29 2175 29 sky130_fd_sc_hd__o31ai_1
* cell instance $47278 m0 *1 705.64,165.92
X$47278 29 2219 2015 2271 2272 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $47279 m0 *1 713.92,165.92
X$47279 29 2250 2220 2248 2206 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $47280 m0 *1 717.6,165.92
X$47280 48 2066 2249 2286 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $47282 m0 *1 719.44,165.92
X$47282 29 2301 1013 2211 2250 2286 1843 48 48 29 sky130_fd_sc_hd__a221oi_4
* cell instance $47284 m0 *1 729.56,165.92
X$47284 29 2066 2206 2248 2220 48 2336 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $47285 m0 *1 734.16,165.92
X$47285 29 2009 2287 2072 1090 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $47286 m0 *1 742.44,165.92
X$47286 48 2209 48 29 1785 29 sky130_fd_sc_hd__buf_4
* cell instance $47287 m0 *1 745.2,165.92
X$47287 48 2288 2252 2304 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $47289 m0 *1 747.04,165.92
X$47289 29 2289 2208 2209 2116 48 48 29 sky130_fd_sc_hd__a21boi_4
* cell instance $47290 m0 *1 753.94,165.92
X$47290 29 2128 2223 2372 2315 48 48 29 sky130_fd_sc_hd__o21bai_2
* cell instance $47291 m0 *1 758.08,165.92
X$47291 29 2291 2290 2017 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $47292 m0 *1 768.2,165.92
X$47292 48 2253 2282 2254 2225 2121 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $47294 m0 *1 772.34,165.92
X$47294 48 2054 2255 1941 29 48 2307 29 sky130_fd_sc_hd__a21oi_1
* cell instance $47296 m0 *1 774.64,165.92
X$47296 48 2214 2228 2215 29 48 2185 29 sky130_fd_sc_hd__a21o_1
* cell instance $47297 m0 *1 777.4,165.92
X$47297 29 2193 2258 2215 2334 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $47298 m0 *1 781.08,165.92
X$47298 48 1042 1695 2193 2309 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $47299 m0 *1 782.92,165.92
X$47299 48 2384 2333 2284 2257 2256 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $47300 m0 *1 785.22,165.92
X$47300 29 2233 1941 2185 2160 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $47301 m0 *1 791.2,165.92
X$47301 29 29 2195 48 2230 2258 48 sky130_fd_sc_hd__nor2_2
* cell instance $47302 m0 *1 793.5,165.92
X$47302 29 2231 2233 2232 2283 1697 2040 48 48 29 sky130_fd_sc_hd__o32a_4
* cell instance $47305 m0 *1 802.7,165.92
X$47305 48 2040 1849 2293 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $47307 m0 *1 805.46,165.92
X$47307 48 2197 2259 2306 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $47308 m0 *1 806.84,165.92
X$47308 48 1638 2260 2259 2261 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $47309 m0 *1 808.68,165.92
X$47309 29 2306 2293 2262 2308 2292 2261 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $47310 m0 *1 812.36,165.92
X$47310 48 2293 2085 2197 2261 48 2278 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $47311 m0 *1 814.66,165.92
X$47311 48 2237 2262 2264 2263 29 2163 48 29 sky130_fd_sc_hd__nor4b_1
* cell instance $47312 m0 *1 817.88,165.92
X$47312 48 2067 2265 2267 2266 48 29 2302 29 sky130_fd_sc_hd__o31ai_1
* cell instance $47313 m0 *1 820.64,165.92
X$47313 29 2173 2265 2267 2303 48 48 29 sky130_fd_sc_hd__nor3b_2
* cell instance $47315 m0 *1 826.16,165.92
X$47315 29 2201 1158 2263 2268 2205 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $47317 m0 *1 829.84,165.92
X$47317 48 2297 2263 2269 2275 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $47318 m0 *1 831.68,165.92
X$47318 48 1158 2269 2165 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $47319 m0 *1 833.06,165.92
X$47319 48 2238 2167 2242 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $47320 m0 *1 835.36,165.92
X$47320 48 2181 1950 2242 2146 48 29 29 sky130_fd_sc_hd__or3_1
* cell instance $47321 m0 *1 837.66,165.92
X$47321 48 2181 1950 2167 48 2273 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $47973 r0 *1 707.94,165.92
X$47973 29 2285 2049 2145 2188 2218 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $47974 r0 *1 711.62,165.92
X$47974 48 2220 2248 2285 2299 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $47975 r0 *1 713.46,165.92
X$47975 29 2310 2300 2224 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $47980 r0 *1 724.5,165.92
X$47980 29 2170 2301 2009 2270 2068 2189 48 48 29 sky130_fd_sc_hd__a221oi_2
* cell instance $47981 r0 *1 730.02,165.92
X$47981 48 2009 1090 2112 29 48 2323 29 sky130_fd_sc_hd__a21o_1
* cell instance $47983 r0 *1 733.24,165.92
X$47983 29 2192 2312 1090 2171 2413 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $47984 r0 *1 737.84,165.92
X$47984 29 2388 2287 1785 1670 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $47985 r0 *1 743.82,165.92
X$47985 48 2222 2221 1445 48 2425 29 29 sky130_fd_sc_hd__o21ai_0
* cell instance $47986 r0 *1 745.66,165.92
X$47986 29 2351 2326 2352 2289 48 48 29 sky130_fd_sc_hd__mux2i_4
* cell instance $47990 r0 *1 753.94,165.92
X$47990 48 2192 2305 1785 29 2252 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $47991 r0 *1 757.16,165.92
X$47991 48 1961 2277 2329 48 29 2290 29 sky130_fd_sc_hd__a21o_2
* cell instance $47993 r0 *1 760.84,165.92
X$47993 29 2290 2291 1980 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $47994 r0 *1 770.96,165.92
X$47994 48 2363 2317 2331 1445 2332 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $47996 r0 *1 773.72,165.92
X$47996 48 1806 2254 1042 29 2215 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $48000 r0 *1 776.94,165.92
X$48000 29 1699 2232 1695 2193 2307 48 48 29 sky130_fd_sc_hd__o31ai_4
* cell instance $48001 r0 *1 784.76,165.92
X$48001 48 2255 2216 1160 2284 2257 48 2367 29 29 sky130_fd_sc_hd__o2111ai_1
* cell instance $48003 r0 *1 788.44,165.92
X$48003 48 1752 48 29 1750 29 sky130_fd_sc_hd__buf_4
* cell instance $48006 r0 *1 795.34,165.92
X$48006 48 1699 48 29 1697 29 sky130_fd_sc_hd__buf_4
* cell instance $48007 r0 *1 798.1,165.92
X$48007 29 2308 1598 1697 2136 2347 48 48 29 sky130_fd_sc_hd__a31o_1
* cell instance $48012 r0 *1 802.24,165.92
X$48012 48 1849 2318 48 2328 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $48014 r0 *1 805.92,165.92
X$48014 48 2197 2381 2327 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $48016 r0 *1 808.68,165.92
X$48016 29 2266 2306 2293 2308 2292 2261 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $48017 r0 *1 811.9,165.92
X$48017 48 2293 2261 2294 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $48019 r0 *1 813.74,165.92
X$48019 48 2076 2294 2327 2166 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $48021 r0 *1 816.04,165.92
X$48021 48 2264 2263 2295 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $48022 r0 *1 817.42,165.92
X$48022 48 2262 2067 1731 29 48 2303 29 sky130_fd_sc_hd__a21oi_1
* cell instance $48023 r0 *1 819.26,165.92
X$48023 29 2322 2296 2324 2067 1731 48 48 29 sky130_fd_sc_hd__o211a_1
* cell instance $48024 r0 *1 822.94,165.92
X$48024 48 2297 1788 2296 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $48025 r0 *1 825.24,165.92
X$48025 48 2264 2263 2320 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $48026 r0 *1 826.62,165.92
X$48026 48 2302 2275 2167 48 29 29 sky130_fd_sc_hd__and2_0
* cell instance $48030 r0 *1 828.92,165.92
X$48030 48 2269 1158 2263 2264 29 48 2298 29 sky130_fd_sc_hd__a31oi_1
* cell instance $48031 r0 *1 831.22,165.92
X$48031 48 2269 1158 2263 2264 29 48 2319 29 sky130_fd_sc_hd__and4_1
* cell instance $48033 r0 *1 835.36,165.92
X$48033 48 2298 2147 2319 48 29 2168 29 sky130_fd_sc_hd__o21ai_1
* cell instance $48990 r0 *1 711.62,171.36
X$48990 48 2299 2349 2348 2370 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $48991 m0 *1 711.62,171.36
X$48991 48 2171 2170 2300 2348 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $48992 m0 *1 713.46,171.36
X$48992 29 2310 2170 2148 2107 2250 48 48 29 sky130_fd_sc_hd__nor4b_2
* cell instance $48993 r0 *1 713.46,171.36
X$48993 48 2148 2107 2285 2300 2349 48 29 29 sky130_fd_sc_hd__o211ai_1
* cell instance $48995 r0 *1 716.68,171.36
X$48995 48 2066 2049 2312 29 48 29 sky130_fd_sc_hd__nand2b_1
* cell instance $48996 r0 *1 718.98,171.36
X$48996 29 2369 2251 2145 2068 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $48998 m0 *1 719.44,171.36
X$48998 29 2274 2249 2321 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $49000 r0 *1 722.66,171.36
X$49000 48 2251 2068 2145 29 48 2335 29 sky130_fd_sc_hd__a21o_1
* cell instance $49001 r0 *1 725.42,171.36
X$49001 29 2380 2369 2335 2336 1013 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $49002 m0 *1 729.56,171.36
X$49002 29 2338 2337 1042 2313 2314 2311 48 48 29 sky130_fd_sc_hd__o32ai_4
* cell instance $49004 r0 *1 730.48,171.36
X$49004 29 29 2338 48 2008 2287 48 sky130_fd_sc_hd__nor2_2
* cell instance $49006 r0 *1 733.24,171.36
X$49006 29 2350 2009 2112 1090 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $49007 r0 *1 736.92,171.36
X$49007 29 2287 2311 2350 2323 48 48 29 sky130_fd_sc_hd__a21boi_2
* cell instance $49008 m0 *1 739.68,171.36
X$49008 48 2208 2221 2222 48 2337 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $49010 r0 *1 741.98,171.36
X$49010 29 2313 2353 2325 2288 2339 48 48 29 sky130_fd_sc_hd__a22oi_4
* cell instance $49012 m0 *1 743.36,171.36
X$49012 48 1670 980 1785 48 2325 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $49014 m0 *1 747.04,171.36
X$49014 29 2289 2276 2291 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $49017 r0 *1 750.26,171.36
X$49017 29 2390 2326 2357 2359 1805 1975 48 48 29 sky130_fd_sc_hd__a41oi_4
* cell instance $49018 m0 *1 757.16,171.36
X$49018 48 2359 2304 2315 29 48 2329 29 sky130_fd_sc_hd__a21o_1
* cell instance $49021 m0 *1 760.38,171.36
X$49021 29 2316 2044 1805 2291 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $49022 r0 *1 760.84,171.36
X$49022 29 2376 2291 1805 2044 2317 48 48 29 sky130_fd_sc_hd__a31oi_2
* cell instance $49023 m0 *1 764.06,171.36
X$49023 48 1747 2316 48 2363 29 29 sky130_fd_sc_hd__and2_2
* cell instance $49024 r0 *1 765.44,171.36
X$49024 29 2363 2375 2216 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $49025 m0 *1 766.82,171.36
X$49025 29 2193 2363 2317 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $49030 m0 *1 774.64,171.36
X$49030 48 2053 1980 2334 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $49031 r0 *1 775.56,171.36
X$49031 29 2364 2385 1160 2230 2366 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $49032 m0 *1 777.86,171.36
X$49032 29 2340 2054 1160 2216 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $49033 m0 *1 781.54,171.36
X$49033 48 2054 2216 2255 2333 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $49034 m0 *1 783.38,171.36
X$49034 29 2309 2340 2367 2256 48 2283 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $49035 r0 *1 783.38,171.36
X$49035 29 2342 2230 2258 2229 1980 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $49038 r0 *1 788.44,171.36
X$49038 48 2258 2230 2395 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $49039 m0 *1 788.9,171.36
X$49039 48 2258 2230 2229 1980 48 2345 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $49040 r0 *1 790.74,171.36
X$49040 48 2341 1699 2368 2383 29 2343 48 29 sky130_fd_sc_hd__a211oi_1
* cell instance $49041 m0 *1 792.12,171.36
X$49041 48 2258 2229 1980 29 48 2330 29 sky130_fd_sc_hd__a21oi_1
* cell instance $49042 r0 *1 793.5,171.36
X$49042 48 2019 2210 2342 2344 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $49043 m0 *1 793.96,171.36
X$49043 48 2158 2136 2345 29 48 2365 29 sky130_fd_sc_hd__a21oi_1
* cell instance $49044 r0 *1 795.34,171.36
X$49044 48 2365 1697 2344 29 48 2381 29 sky130_fd_sc_hd__a21oi_1
* cell instance $49045 m0 *1 795.8,171.36
X$49045 48 1750 2343 2318 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $49048 r0 *1 797.64,171.36
X$49048 29 2362 1699 1752 2346 2347 48 48 29 sky130_fd_sc_hd__nor4_2
* cell instance $49053 r0 *1 802.24,171.36
X$49053 48 2361 2360 2260 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $49054 m0 *1 802.7,171.36
X$49054 48 2318 2088 2358 29 48 29 sky130_fd_sc_hd__nor2b_1
* cell instance $49056 r0 *1 805.46,171.36
X$49056 29 2292 2356 2162 2263 2358 2328 48 48 29 sky130_fd_sc_hd__o32ai_4
* cell instance $49057 m0 *1 805.46,171.36
X$49057 29 2292 2040 2162 2108 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $49059 m0 *1 810.06,171.36
X$49059 29 2108 2356 2040 2318 48 48 29 sky130_fd_sc_hd__and3_1
* cell instance $49061 m0 *1 812.82,171.36
X$49061 29 2355 2205 2327 2354 48 48 29 sky130_fd_sc_hd__a21boi_2
* cell instance $49066 m0 *1 818.34,171.36
X$49066 48 1788 2295 2324 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $49067 m0 *1 819.72,171.36
X$49067 29 2265 2322 2303 2297 2199 2320 48 48 29 sky130_fd_sc_hd__a311oi_4
* cell instance $49070 r0 *1 821.1,171.36
X$49070 48 2297 2263 2267 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $49073 r0 *1 825.24,171.36
X$49073 48 2067 1731 2268 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $49074 r0 *1 826.62,171.36
X$49074 48 1731 1788 2269 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $49075 r0 *1 828,171.36
X$49075 48 2264 48 29 2297 29 sky130_fd_sc_hd__inv_1
* cell instance $50061 m0 *1 719.9,176.8
X$50061 48 2218 1843 2312 2387 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $50064 m0 *1 721.74,176.8
X$50064 48 2211 2370 2387 2398 48 29 29 sky130_fd_sc_hd__o21ba_1
* cell instance $50065 m0 *1 725.42,176.8
X$50065 29 2369 2335 2336 48 2406 48 29 sky130_fd_sc_hd__nand3_4
* cell instance $50066 m0 *1 731.86,176.8
X$50066 29 2209 2211 2370 2387 48 48 29 sky130_fd_sc_hd__o21bai_2
* cell instance $50067 m0 *1 736,176.8
X$50067 29 2350 2371 2323 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $50068 m0 *1 740.14,176.8
X$50068 48 2222 2221 2208 2314 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $50070 m0 *1 742.9,176.8
X$50070 48 2222 2371 2221 48 29 2351 29 sky130_fd_sc_hd__o21ai_1
* cell instance $50071 m0 *1 744.74,176.8
X$50071 48 2315 2277 2389 48 29 2386 29 sky130_fd_sc_hd__o21ai_1
* cell instance $50073 m0 *1 747.04,176.8
X$50073 29 29 2353 48 2073 1918 48 sky130_fd_sc_hd__nor2_2
* cell instance $50076 m0 *1 749.34,176.8
X$50076 29 2326 2390 1961 1445 2372 2288 48 48 29 sky130_fd_sc_hd__a311oi_4
* cell instance $50077 m0 *1 759,176.8
X$50077 48 1805 2326 2357 1975 48 2389 29 29 sky130_fd_sc_hd__nand4_1
* cell instance $50078 m0 *1 761.3,176.8
X$50078 48 2375 2374 2373 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $50079 m0 *1 762.68,176.8
X$50079 29 2401 2400 2316 2377 2376 48 48 29 sky130_fd_sc_hd__a2bb2oi_1
* cell instance $50080 m0 *1 765.9,176.8
X$50080 48 2317 2374 2377 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $50082 m0 *1 768.2,176.8
X$50082 48 2375 1674 2331 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $50084 m0 *1 770.5,176.8
X$50084 48 2374 2402 2316 2379 2331 2385 29 48 29 sky130_fd_sc_hd__a311o_1
* cell instance $50088 m0 *1 774.64,176.8
X$50088 29 2404 2374 2378 1042 2017 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $50089 m0 *1 779.24,176.8
X$50089 48 1160 2216 2384 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $50090 m0 *1 780.62,176.8
X$50090 29 2340 2392 2360 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $50091 m0 *1 790.74,176.8
X$50091 29 2395 1752 2257 48 48 29 sky130_fd_sc_hd__nor2_4
* cell instance $50093 m0 *1 795.34,176.8
X$50093 48 2396 2347 2403 48 2397 29 29 sky130_fd_sc_hd__a21oi_2
* cell instance $50094 m0 *1 798.56,176.8
X$50094 48 2397 2362 2382 29 2259 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $50098 m0 *1 802.24,176.8
X$50098 29 2360 2361 2162 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $50099 m0 *1 812.36,176.8
X$50099 48 2108 2162 2040 2318 29 48 2355 29 sky130_fd_sc_hd__a31oi_1
* cell instance $50778 r0 *1 724.5,176.8
X$50778 29 2398 1918 48 48 29 sky130_fd_sc_hd__buf_6
* cell instance $50781 r0 *1 730.94,176.8
X$50781 48 2171 1090 2312 29 48 2413 29 sky130_fd_sc_hd__a21oi_1
* cell instance $50784 r0 *1 733.7,176.8
X$50784 29 2338 980 2073 1918 2416 48 48 29 sky130_fd_sc_hd__o22ai_4
* cell instance $50785 r0 *1 741.06,176.8
X$50785 29 2371 2388 2375 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $50787 r0 *1 751.18,176.8
X$50787 48 2399 2325 2400 29 48 29 sky130_fd_sc_hd__or2_1
* cell instance $50789 r0 *1 754.4,176.8
X$50789 29 2391 2390 2386 2408 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $50791 r0 *1 760.84,176.8
X$50791 29 1747 2317 2376 48 2378 48 29 sky130_fd_sc_hd__mux2i_2
* cell instance $50792 r0 *1 765.9,176.8
X$50792 48 2317 1031 2415 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $50793 r0 *1 767.28,176.8
X$50793 48 2419 2378 1042 2391 29 2402 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $50795 r0 *1 770.04,176.8
X$50795 29 2392 2331 2374 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $50797 r0 *1 776.02,176.8
X$50797 48 2392 1806 1810 2379 29 2366 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $50799 r0 *1 780.16,176.8
X$50799 29 2423 2393 2405 2410 48 2019 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $50801 r0 *1 788.44,176.8
X$50801 29 2382 1597 2342 2394 2411 2414 48 48 29 sky130_fd_sc_hd__o311a_1
* cell instance $50802 r0 *1 792.12,176.8
X$50802 48 2233 2360 2341 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $50803 r0 *1 793.5,176.8
X$50803 29 1752 2330 1699 2361 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $50804 r0 *1 799.48,176.8
X$50804 29 2397 2362 2197 2382 48 2088 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $50806 r0 *1 807.3,176.8
X$50806 48 2362 2397 2354 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $50809 r0 *1 812.36,176.8
X$50809 48 2355 2412 2076 29 2264 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $51485 m0 *1 727.72,182.24
X$51485 48 2406 2338 48 2407 29 29 sky130_fd_sc_hd__xor2_1
* cell instance $51486 m0 *1 730.94,182.24
X$51486 29 2407 2353 2357 2325 2380 48 48 29 sky130_fd_sc_hd__a22o_2
* cell instance $51487 m0 *1 734.62,182.24
X$51487 29 2388 2371 2317 48 48 29 sky130_fd_sc_hd__xnor2_4
* cell instance $51488 m0 *1 744.74,182.24
X$51488 48 2338 2276 2311 48 29 2352 29 sky130_fd_sc_hd__o21ai_1
* cell instance $51490 m0 *1 747.04,182.24
X$51490 29 29 2374 48 2325 2399 48 sky130_fd_sc_hd__nor2_2
* cell instance $51493 m0 *1 749.34,182.24
X$51493 29 2326 1961 1445 2408 2288 48 48 29 sky130_fd_sc_hd__a31oi_4
* cell instance $51494 m0 *1 757.16,182.24
X$51494 48 2426 48 29 1674 29 sky130_fd_sc_hd__buf_4
* cell instance $51495 m0 *1 759.92,182.24
X$51495 48 2315 2389 2418 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $51496 m0 *1 761.3,182.24
X$51496 29 2417 2418 2408 2076 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $51497 m0 *1 767.28,182.24
X$51497 29 2316 2409 2400 2415 48 48 29 sky130_fd_sc_hd__nor3_2
* cell instance $51498 m0 *1 770.96,182.24
X$51498 48 2420 2400 2379 2332 48 2364 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $51502 m0 *1 774.64,182.24
X$51502 48 2225 2254 2393 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $51503 m0 *1 776.02,182.24
X$51503 29 2404 2437 2410 2409 2054 2053 48 48 29 sky130_fd_sc_hd__o221ai_4
* cell instance $51504 m0 *1 785.68,182.24
X$51504 29 2394 2158 2233 2360 2136 48 48 29 sky130_fd_sc_hd__a2bb2oi_1
* cell instance $51505 m0 *1 788.9,182.24
X$51505 48 2368 2383 2395 2257 2411 29 48 29 sky130_fd_sc_hd__o22ai_1
* cell instance $51506 m0 *1 791.2,182.24
X$51506 29 2414 2210 2342 2383 2368 2019 48 48 29 sky130_fd_sc_hd__o41ai_1
* cell instance $51507 m0 *1 794.42,182.24
X$51507 48 2158 48 29 2210 29 sky130_fd_sc_hd__inv_1
* cell instance $51508 m0 *1 795.8,182.24
X$51508 48 1597 2342 2424 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $51510 m0 *1 798.1,182.24
X$51510 48 2346 2424 2412 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $52199 r0 *1 729.56,182.24
X$52199 48 2073 1918 2380 29 2428 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $52201 r0 *1 733.24,182.24
X$52201 29 2406 2416 2390 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $52202 r0 *1 743.36,182.24
X$52202 48 1013 2371 2425 29 48 2339 29 sky130_fd_sc_hd__a21oi_1
* cell instance $52203 r0 *1 745.2,182.24
X$52203 48 1013 2073 1918 2399 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $52204 r0 *1 747.04,182.24
X$52204 29 1918 2281 2073 2430 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $52207 r0 *1 753.94,182.24
X$52207 29 2359 2277 2315 2431 48 48 29 sky130_fd_sc_hd__o21ai_4
* cell instance $52210 r0 *1 760.84,182.24
X$52210 29 2426 2277 2359 2315 2417 2408 48 48 29 sky130_fd_sc_hd__o221a_1
* cell instance $52211 r0 *1 764.98,182.24
X$52211 48 2427 2315 2277 29 48 2419 29 sky130_fd_sc_hd__a21oi_1
* cell instance $52212 r0 *1 766.82,182.24
X$52212 48 2415 2391 2316 2419 29 2420 48 29 sky130_fd_sc_hd__nor4_1
* cell instance $52213 r0 *1 769.12,182.24
X$52213 48 2419 2391 2379 29 48 29 sky130_fd_sc_hd__or2_0
* cell instance $52214 r0 *1 771.42,182.24
X$52214 48 2391 2419 2422 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $52215 r0 *1 772.8,182.24
X$52215 48 2153 2438 2421 48 29 1809 29 sky130_fd_sc_hd__o21ba_2
* cell instance $52217 r0 *1 776.48,182.24
X$52217 48 2409 2404 2053 2054 2423 29 48 29 sky130_fd_sc_hd__o22a_1
* cell instance $52218 r0 *1 779.7,182.24
X$52218 48 2422 2423 1695 48 2368 29 29 sky130_fd_sc_hd__o21a_1
* cell instance $52219 r0 *1 782.46,182.24
X$52219 48 1695 2422 2423 2383 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $52220 r0 *1 784.3,182.24
X$52220 48 2405 2410 2393 2423 48 29 2136 29 sky130_fd_sc_hd__o211a_2
* cell instance $52224 r0 *1 791.2,182.24
X$52224 48 2346 2345 2136 2247 48 2396 29 29 sky130_fd_sc_hd__a211o_1
* cell instance $52225 r0 *1 794.42,182.24
X$52225 48 2019 2345 2346 2403 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $53200 m0 *1 732.32,187.68
X$53200 48 2428 2321 2435 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $53204 r0 *1 734.16,187.68
X$53204 29 2443 2416 2406 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $53205 m0 *1 735.54,187.68
X$53205 29 2321 2428 2429 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $53206 r0 *1 740.14,187.68
X$53206 29 2224 2430 2441 48 48 29 sky130_fd_sc_hd__xor2_4
* cell instance $53213 m0 *1 747.96,187.68
X$53213 29 2252 2443 2441 2429 48 2417 48 29 sky130_fd_sc_hd__nand4_2
* cell instance $53214 r0 *1 750.26,187.68
X$53214 48 2353 29 48 1146 29 sky130_fd_sc_hd__inv_2
* cell instance $53215 r0 *1 751.64,187.68
X$53215 29 2279 2450 2435 2357 2317 48 48 29 sky130_fd_sc_hd__a211oi_2
* cell instance $53216 m0 *1 752.56,187.68
X$53216 29 2373 1445 2439 2431 2443 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $53217 r0 *1 756.24,187.68
X$53217 29 2431 2442 2372 2401 1042 2433 48 48 29 sky130_fd_sc_hd__o221a_2
* cell instance $53218 m0 *1 759.92,187.68
X$53218 48 2408 2390 2427 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $53221 m0 *1 761.3,187.68
X$53221 29 2449 2431 2254 2391 2461 48 48 29 sky130_fd_sc_hd__a211oi_4
* cell instance $53222 r0 *1 761.3,187.68
X$53222 29 2253 1674 2401 2453 2448 48 48 29 sky130_fd_sc_hd__o31a_1
* cell instance $53223 r0 *1 764.52,187.68
X$53223 48 2427 2455 2449 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $53225 r0 *1 766.36,187.68
X$53225 29 2444 2429 2452 1747 48 48 29 sky130_fd_sc_hd__nand3_2
* cell instance $53227 m0 *1 769.12,187.68
X$53227 48 2445 2444 2432 48 29 29 sky130_fd_sc_hd__and2_1
* cell instance $53228 r0 *1 770.04,187.68
X$53228 29 2433 2439 2444 2445 48 1808 48 29 sky130_fd_sc_hd__o211ai_4
* cell instance $53230 m0 *1 772.34,187.68
X$53230 48 2434 2440 2446 48 29 2437 29 sky130_fd_sc_hd__o21ai_1
* cell instance $53235 m0 *1 774.64,187.68
X$53235 29 2432 2436 2225 2422 2433 2439 48 48 29 sky130_fd_sc_hd__o221ai_2
* cell instance $53237 r0 *1 778.32,187.68
X$53237 48 2434 2438 2421 2440 48 29 2459 29 sky130_fd_sc_hd__o31ai_1
* cell instance $53239 m0 *1 780.62,187.68
X$53239 48 2432 2434 2447 29 48 2346 29 sky130_fd_sc_hd__a21o_1
* cell instance $53240 r0 *1 781.08,187.68
X$53240 29 1810 2445 2444 2433 2439 48 48 29 sky130_fd_sc_hd__o211a_4
* cell instance $53242 m0 *1 783.84,187.68
X$53242 29 29 2347 48 1810 2440 48 sky130_fd_sc_hd__nor2_2
* cell instance $54636 m0 *1 747.04,193.12
X$54636 29 2450 2430 2224 48 48 29 sky130_fd_sc_hd__xnor2_2
* cell instance $54640 r0 *1 747.96,193.12
X$54640 29 2441 2315 2429 48 48 29 sky130_fd_sc_hd__nand2_4
* cell instance $54642 r0 *1 752.56,193.12
X$54642 29 29 2451 48 2435 2372 48 sky130_fd_sc_hd__nor2_2
* cell instance $54644 m0 *1 753.48,193.12
X$54644 48 2451 2450 2453 48 29 29 sky130_fd_sc_hd__xnor2_1
* cell instance $54646 r0 *1 755.32,193.12
X$54646 48 2429 2372 2460 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $54647 r0 *1 756.7,193.12
X$54647 48 2408 2443 2442 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $54650 m0 *1 758.08,193.12
X$54650 29 2315 2454 2357 1674 2451 2317 48 48 29 sky130_fd_sc_hd__a2111oi_0
* cell instance $54652 r0 *1 758.54,193.12
X$54652 48 2450 1674 2373 2448 48 29 29 sky130_fd_sc_hd__nand3_1
* cell instance $54654 r0 *1 760.84,193.12
X$54654 48 2429 2441 2452 2315 48 29 2462 29 sky130_fd_sc_hd__o31ai_1
* cell instance $54655 m0 *1 761.3,193.12
X$54655 29 2446 2456 2429 2454 2458 2457 48 48 29 sky130_fd_sc_hd__a221oi_1
* cell instance $54656 r0 *1 763.6,193.12
X$54656 48 2441 1031 2457 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $54657 m0 *1 764.52,193.12
X$54657 48 2429 2452 2455 48 29 29 sky130_fd_sc_hd__nand2_1
* cell instance $54658 r0 *1 764.98,193.12
X$54658 48 2429 2452 1031 29 48 2461 29 sky130_fd_sc_hd__a21oi_1
* cell instance $54659 m0 *1 765.9,193.12
X$54659 29 2438 2441 1747 2451 48 48 29 sky130_fd_sc_hd__a21oi_4
* cell instance $54660 r0 *1 766.82,193.12
X$54660 48 2452 1747 2429 29 48 2445 29 sky130_fd_sc_hd__a21o_1
* cell instance $54661 r0 *1 769.58,193.12
X$54661 48 2441 2451 1747 29 48 2421 29 sky130_fd_sc_hd__and3_2
* cell instance $54663 m0 *1 772.34,193.12
X$54663 48 2438 2153 2421 48 29 2440 29 sky130_fd_sc_hd__o21ai_1
* cell instance $54664 r0 *1 772.34,193.12
X$54664 29 29 2225 48 2438 2421 48 sky130_fd_sc_hd__nor2_2
* cell instance $54670 m0 *1 774.64,193.12
X$54670 29 2153 1806 2421 2438 48 48 29 sky130_fd_sc_hd__o21bai_4
* cell instance $54672 r0 *1 778.78,193.12
X$54672 48 2433 2439 2434 29 48 29 sky130_fd_sc_hd__nor2_1
* cell instance $54673 r0 *1 780.16,193.12
X$54673 48 2432 2434 1809 2447 29 48 29 sky130_fd_sc_hd__nor3_1
* cell instance $54674 m0 *1 781.54,193.12
X$54674 48 2432 2459 2436 29 2405 48 29 sky130_fd_sc_hd__o21ai_2
* cell instance $56079 m0 *1 755.32,198.56
X$56079 29 1031 2357 2456 2441 2460 2317 48 48 29 sky130_fd_sc_hd__a221o_1
* cell instance $56081 m0 *1 759,198.56
X$56081 29 29 2317 2452 2357 48 48 sky130_fd_sc_hd__nand2_2
* cell instance $56086 m0 *1 761.3,198.56
X$56086 48 1031 2452 2441 2462 29 48 2458 29 sky130_fd_sc_hd__a31oi_1
* cell instance $223842 r0 *1 4.14,840.48
X$223842 29 2463 206 48 48 29 sky130_fd_sc_hd__buf_16
* cell instance $225268 m0 *1 5.98,845.92
X$225268 29 2464 178 48 48 29 sky130_fd_sc_hd__buf_16
.ENDS parameterized_freq_divider

* cell sky130_fd_sc_hd__a222oi_1
* pin VGND
* pin Y
* pin C1
* pin C2
* pin B2
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a222oi_1 1 2 3 4 5 6 7 8 14 15 16
* net 1 VGND
* net 2 Y
* net 3 C1
* net 4 C2
* net 5 B2
* net 6 B1
* net 7 A1
* net 8 A2
* net 14 VPWR
* net 15 VPB
* device instance $1 r0 *1 1.89,1.985 pfet_01v8_hvt
M$1 12 5 13 15 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.31,1.985 pfet_01v8_hvt
M$2 13 6 12 15 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 2.73,1.985 pfet_01v8_hvt
M$3 14 7 13 15 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $4 r0 *1 3.21,1.985 pfet_01v8_hvt
M$4 13 8 14 15 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=260000000000P PS=1330000U PD=2520000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 12 3 2 15 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $6 r0 *1 0.89,1.985 pfet_01v8_hvt
M$6 2 4 12 15 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $7 r0 *1 0.47,0.555 nfet_01v8
M$7 9 3 2 16 nfet_01v8 L=150000U W=640000U AS=166400000000P AD=67200000000P
+ PS=1800000U PD=850000U
* device instance $8 r0 *1 0.83,0.555 nfet_01v8
M$8 1 4 9 16 nfet_01v8 L=150000U W=640000U AS=67200000000P AD=291200000000P
+ PS=850000U PD=1550000U
* device instance $9 r0 *1 1.89,0.555 nfet_01v8
M$9 11 5 1 16 nfet_01v8 L=150000U W=640000U AS=291200000000P AD=67200000000P
+ PS=1550000U PD=850000U
* device instance $10 r0 *1 2.25,0.555 nfet_01v8
M$10 2 6 11 16 nfet_01v8 L=150000U W=640000U AS=67200000000P AD=105600000000P
+ PS=850000U PD=970000U
* device instance $11 r0 *1 2.73,0.555 nfet_01v8
M$11 10 7 2 16 nfet_01v8 L=150000U W=640000U AS=105600000000P AD=105600000000P
+ PS=970000U PD=970000U
* device instance $12 r0 *1 3.21,0.555 nfet_01v8
M$12 1 8 10 16 nfet_01v8 L=150000U W=640000U AS=105600000000P AD=166400000000P
+ PS=970000U PD=1800000U
.ENDS sky130_fd_sc_hd__a222oi_1

* cell sky130_fd_sc_hd__dlymetal6s2s_1
* pin VGND
* pin X
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 1 3 8 9 10 11
* net 1 VGND
* net 3 X
* net 8 A
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 3.655,2.275 pfet_01v8_hvt
M$1 6 5 9 10 pfet_01v8_hvt L=150000U W=420000U AS=140750000000P
+ AD=109200000000P PS=1325000U PD=1360000U
* device instance $2 r0 *1 4.13,1.985 pfet_01v8_hvt
M$2 7 6 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $3 r0 *1 2.24,2.275 pfet_01v8_hvt
M$3 4 3 9 10 pfet_01v8_hvt L=150000U W=420000U AS=140750000000P
+ AD=109200000000P PS=1325000U PD=1360000U
* device instance $4 r0 *1 2.715,1.985 pfet_01v8_hvt
M$4 5 4 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $5 r0 *1 0.645,2.275 pfet_01v8_hvt
M$5 2 8 9 10 pfet_01v8_hvt L=150000U W=420000U AS=140750000000P
+ AD=109200000000P PS=1325000U PD=1360000U
* device instance $6 r0 *1 1.12,1.985 pfet_01v8_hvt
M$6 3 2 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $7 r0 *1 3.655,0.445 nfet_01v8
M$7 1 5 6 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $8 r0 *1 4.13,0.56 nfet_01v8
M$8 7 6 1 11 nfet_01v8 L=150000U W=650000U AS=97000000000P AD=169000000000P
+ PS=975000U PD=1820000U
* device instance $9 r0 *1 0.645,0.445 nfet_01v8
M$9 1 8 2 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $10 r0 *1 1.12,0.56 nfet_01v8
M$10 3 2 1 11 nfet_01v8 L=150000U W=650000U AS=97000000000P AD=169000000000P
+ PS=975000U PD=1820000U
* device instance $11 r0 *1 2.24,0.445 nfet_01v8
M$11 1 3 4 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $12 r0 *1 2.715,0.56 nfet_01v8
M$12 5 4 1 11 nfet_01v8 L=150000U W=650000U AS=97000000000P AD=169000000000P
+ PS=975000U PD=1820000U
.ENDS sky130_fd_sc_hd__dlymetal6s2s_1

* cell sky130_fd_sc_hd__clkbuf_2
* pin VPB
* pin A
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_2 1 2 3 4 6 7
* net 1 VPB
* net 2 A
* net 3 VPWR
* net 4 VGND
* net 6 X
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 3 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=162500000000P PS=2530000U PD=1325000U
* device instance $2 r0 *1 0.95,1.985 pfet_01v8_hvt
M$2 6 5 3 1 pfet_01v8_hvt L=150000U W=2000000U AS=297500000000P
+ AD=395000000000P PS=2595000U PD=3790000U
* device instance $4 r0 *1 0.475,0.445 nfet_01v8
M$4 4 2 5 7 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=68250000000P
+ PS=1370000U PD=745000U
* device instance $5 r0 *1 0.95,0.445 nfet_01v8
M$5 6 5 4 7 nfet_01v8 L=150000U W=840000U AS=124950000000P AD=165900000000P
+ PS=1435000U PD=2050000U
.ENDS sky130_fd_sc_hd__clkbuf_2

* cell sky130_fd_sc_hd__o41ai_4
* pin VGND
* pin B1
* pin A4
* pin A3
* pin A1
* pin Y
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o41ai_4 1 2 3 4 5 7 8 9 13 14
* net 1 VGND
* net 2 B1
* net 3 A4
* net 4 A3
* net 5 A1
* net 7 Y
* net 8 A2
* net 9 VPWR
* net 13 VPB
* device instance $1 r0 *1 6.55,1.985 pfet_01v8_hvt
M$1 11 8 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 8.23,1.985 pfet_01v8_hvt
M$5 9 5 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=685000000000P PS=5080000U PD=6370000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 7 2 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=665000000000P PS=6330000U PD=6330000U
* device instance $13 r0 *1 2.67,1.985 pfet_01v8_hvt
M$13 7 3 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $17 r0 *1 4.35,1.985 pfet_01v8_hvt
M$17 11 4 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 6.55,0.56 nfet_01v8
M$21 1 8 6 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $25 r0 *1 8.23,0.56 nfet_01v8
M$25 1 5 6 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=445250000000P
+ PS=3680000U PD=4620000U
* device instance $29 r0 *1 0.47,0.56 nfet_01v8
M$29 7 2 6 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
* device instance $33 r0 *1 2.67,0.56 nfet_01v8
M$33 1 3 6 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $37 r0 *1 4.35,0.56 nfet_01v8
M$37 1 4 6 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__o41ai_4

* cell sky130_fd_sc_hd__and2_4
* pin VPB
* pin A
* pin B
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__and2_4 1 2 3 5 6 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 5 VGND
* net 6 X
* net 7 VPWR
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 4 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 0.905,1.985 pfet_01v8_hvt
M$2 7 3 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=177500000000P PS=1280000U PD=1355000U
* device instance $3 r0 *1 1.41,1.985 pfet_01v8_hvt
M$3 6 4 7 1 pfet_01v8_hvt L=150000U W=4000000U AS=597500000000P
+ AD=705000000000P PS=5195000U PD=6410000U
* device instance $7 r0 *1 0.475,0.56 nfet_01v8
M$7 9 2 4 8 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=68250000000P
+ PS=1830000U PD=860000U
* device instance $8 r0 *1 0.835,0.56 nfet_01v8
M$8 5 3 9 8 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=138125000000P
+ PS=860000U PD=1075000U
* device instance $9 r0 *1 1.41,0.56 nfet_01v8
M$9 6 4 5 8 nfet_01v8 L=150000U W=2600000U AS=411125000000P AD=458250000000P
+ PS=3865000U PD=4660000U
.ENDS sky130_fd_sc_hd__and2_4

* cell sky130_fd_sc_hd__nand4b_2
* pin VGND
* pin Y
* pin A_N
* pin B
* pin C
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand4b_2 1 4 7 8 9 10 11 12 13
* net 1 VGND
* net 4 Y
* net 7 A_N
* net 8 B
* net 9 C
* net 10 D
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 1.41,1.985 pfet_01v8_hvt
M$1 4 2 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 2.25,1.985 pfet_01v8_hvt
M$3 4 8 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=505000000000P PS=2540000U PD=3010000U
* device instance $5 r0 *1 3.56,1.985 pfet_01v8_hvt
M$5 4 9 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=505000000000P
+ AD=315000000000P PS=3010000U PD=2630000U
* device instance $7 r0 *1 4.49,1.985 pfet_01v8_hvt
M$7 4 10 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=315000000000P
+ AD=535000000000P PS=2630000U PD=4070000U
* device instance $9 r0 *1 0.47,2.275 pfet_01v8_hvt
M$9 11 7 2 12 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=109200000000P PS=1360000U PD=1360000U
* device instance $10 r0 *1 3.61,0.56 nfet_01v8
M$10 5 9 6 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=204750000000P
+ PS=2740000U PD=1930000U
* device instance $12 r0 *1 4.54,0.56 nfet_01v8
M$12 1 10 6 13 nfet_01v8 L=150000U W=1300000U AS=204750000000P AD=256750000000P
+ PS=1930000U PD=2740000U
* device instance $14 r0 *1 1.41,0.56 nfet_01v8
M$14 4 2 3 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $16 r0 *1 2.25,0.56 nfet_01v8
M$16 5 8 3 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $18 r0 *1 0.47,0.445 nfet_01v8
M$18 1 7 2 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__nand4b_2

* cell sky130_fd_sc_hd__o41a_2
* pin VGND
* pin X
* pin B1
* pin A4
* pin A3
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o41a_2 1 2 5 6 7 8 9 10 11 15
* net 1 VGND
* net 2 X
* net 5 B1
* net 6 A4
* net 7 A3
* net 8 A2
* net 9 A1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 2 3 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=440000000000P PS=3790000U PD=2880000U
* device instance $3 r0 *1 1.65,1.985 pfet_01v8_hvt
M$3 3 5 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=305000000000P
+ AD=302500000000P PS=1610000U PD=1605000U
* device instance $4 r0 *1 2.405,1.985 pfet_01v8_hvt
M$4 13 6 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=302500000000P
+ AD=177500000000P PS=1605000U PD=1355000U
* device instance $5 r0 *1 2.91,1.985 pfet_01v8_hvt
M$5 14 7 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=177500000000P
+ AD=175000000000P PS=1355000U PD=1350000U
* device instance $6 r0 *1 3.41,1.985 pfet_01v8_hvt
M$6 12 8 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=175000000000P
+ AD=175000000000P PS=1350000U PD=1350000U
* device instance $7 r0 *1 3.91,1.985 pfet_01v8_hvt
M$7 10 9 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=175000000000P
+ AD=410000000000P PS=1350000U PD=2820000U
* device instance $8 r0 *1 1.89,0.56 nfet_01v8
M$8 4 5 3 15 nfet_01v8 L=150000U W=650000U AS=208000000000P AD=118625000000P
+ PS=1940000U PD=1015000U
* device instance $9 r0 *1 2.405,0.56 nfet_01v8
M$9 1 6 4 15 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=115375000000P
+ PS=1015000U PD=1005000U
* device instance $10 r0 *1 2.91,0.56 nfet_01v8
M$10 4 7 1 15 nfet_01v8 L=150000U W=650000U AS=115375000000P AD=113750000000P
+ PS=1005000U PD=1000000U
* device instance $11 r0 *1 3.41,0.56 nfet_01v8
M$11 1 8 4 15 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=113750000000P
+ PS=1000000U PD=1000000U
* device instance $12 r0 *1 3.91,0.56 nfet_01v8
M$12 4 9 1 15 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=266500000000P
+ PS=1000000U PD=2120000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 2 3 1 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
.ENDS sky130_fd_sc_hd__o41a_2

* cell sky130_fd_sc_hd__a22oi_1
* pin VPB
* pin B2
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a22oi_1 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 7 VPWR
* net 8 Y
* net 9 VGND
* device instance $1 r0 *1 1.83,1.985 pfet_01v8_hvt
M$1 6 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.25,1.985 pfet_01v8_hvt
M$2 7 5 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=300000000000P PS=1270000U PD=2600000U
* device instance $3 r0 *1 0.47,1.985 pfet_01v8_hvt
M$3 6 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $4 r0 *1 0.89,1.985 pfet_01v8_hvt
M$4 8 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $5 r0 *1 1.83,0.56 nfet_01v8
M$5 11 4 8 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=68250000000P
+ PS=1820000U PD=860000U
* device instance $6 r0 *1 2.19,0.56 nfet_01v8
M$6 9 5 11 10 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=234000000000P
+ PS=860000U PD=2020000U
* device instance $7 r0 *1 0.47,0.56 nfet_01v8
M$7 12 2 9 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=74750000000P
+ PS=1820000U PD=880000U
* device instance $8 r0 *1 0.85,0.56 nfet_01v8
M$8 8 3 12 10 nfet_01v8 L=150000U W=650000U AS=74750000000P AD=169000000000P
+ PS=880000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22oi_1

* cell sky130_fd_sc_hd__nand3b_4
* pin VGND
* pin B
* pin A_N
* pin Y
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand3b_4 1 2 4 6 8 9 10 11
* net 1 VGND
* net 2 B
* net 4 A_N
* net 6 Y
* net 8 C
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 5.29,1.985 pfet_01v8_hvt
M$1 6 8 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=765000000000P PS=6330000U PD=6530000U
* device instance $5 r0 *1 1.41,1.985 pfet_01v8_hvt
M$5 6 3 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $9 r0 *1 3.09,1.985 pfet_01v8_hvt
M$9 6 2 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $13 r0 *1 0.47,1.985 pfet_01v8_hvt
M$13 9 4 3 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $14 r0 *1 5.29,0.56 nfet_01v8
M$14 7 8 1 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=497250000000P
+ PS=4580000U PD=4780000U
* device instance $18 r0 *1 0.47,0.56 nfet_01v8
M$18 1 4 3 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
* device instance $19 r0 *1 1.41,0.56 nfet_01v8
M$19 6 3 5 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $23 r0 *1 3.09,0.56 nfet_01v8
M$23 7 2 5 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nand3b_4

* cell sky130_fd_sc_hd__ha_4
* pin VGND
* pin SUM
* pin B
* pin COUT
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__ha_4 1 3 5 7 8 11 12 15
* net 1 VGND
* net 3 SUM
* net 5 B
* net 7 COUT
* net 8 A
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 3 2 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=787500000000P PS=6330000U PD=5575000U
* device instance $5 r0 *1 2.645,1.985 pfet_01v8_hvt
M$5 2 6 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=517500000000P
+ AD=282500000000P PS=3035000U PD=2565000U
* device instance $7 r0 *1 3.51,1.985 pfet_01v8_hvt
M$7 13 8 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=147500000000P
+ AD=147500000000P PS=1295000U PD=1295000U
* device instance $8 r0 *1 3.955,1.985 pfet_01v8_hvt
M$8 2 5 13 12 pfet_01v8_hvt L=150000U W=1000000U AS=147500000000P
+ AD=135000000000P PS=1295000U PD=1270000U
* device instance $9 r0 *1 4.375,1.985 pfet_01v8_hvt
M$9 14 5 2 12 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=287500000000P PS=1270000U PD=1575000U
* device instance $10 r0 *1 5.1,1.985 pfet_01v8_hvt
M$10 11 8 14 12 pfet_01v8_hvt L=150000U W=1000000U AS=287500000000P
+ AD=230000000000P PS=1575000U PD=1460000U
* device instance $11 r0 *1 5.71,1.985 pfet_01v8_hvt
M$11 6 8 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=365000000000P
+ AD=310000000000P PS=2730000U PD=2620000U
* device instance $12 r0 *1 6.13,1.985 pfet_01v8_hvt
M$12 11 5 6 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $15 r0 *1 7.47,1.985 pfet_01v8_hvt
M$15 7 6 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=580000000000P
+ AD=665000000000P PS=5160000U PD=6330000U
* device instance $19 r0 *1 5.34,0.56 nfet_01v8
M$19 1 8 4 15 nfet_01v8 L=150000U W=1300000U AS=273000000000P AD=183625000000P
+ PS=2790000U PD=1865000U
* device instance $20 r0 *1 5.76,0.56 nfet_01v8
M$20 10 8 1 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=71500000000P
+ PS=920000U PD=870000U
* device instance $21 r0 *1 6.13,0.56 nfet_01v8
M$21 6 5 10 15 nfet_01v8 L=150000U W=650000U AS=71500000000P AD=87750000000P
+ PS=870000U PD=920000U
* device instance $22 r0 *1 6.55,0.56 nfet_01v8
M$22 9 5 6 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $23 r0 *1 6.97,0.56 nfet_01v8
M$23 1 8 9 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=113750000000P
+ PS=920000U PD=1000000U
* device instance $24 r0 *1 7.47,0.56 nfet_01v8
M$24 7 6 1 15 nfet_01v8 L=150000U W=2600000U AS=377000000000P AD=432250000000P
+ PS=3760000U PD=4580000U
* device instance $28 r0 *1 0.47,0.56 nfet_01v8
M$28 3 2 1 15 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
* device instance $32 r0 *1 2.67,0.56 nfet_01v8
M$32 2 6 4 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $35 r0 *1 3.955,0.56 nfet_01v8
M$35 4 5 1 15 nfet_01v8 L=150000U W=1300000U AS=183625000000P AD=256750000000P
+ PS=1865000U PD=2740000U
.ENDS sky130_fd_sc_hd__ha_4

* cell sky130_fd_sc_hd__a21bo_1
* pin VGND
* pin B1_N
* pin X
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a21bo_1 1 2 5 6 7 9 11 12
* net 1 VGND
* net 2 B1_N
* net 5 X
* net 6 A1
* net 7 A2
* net 9 VPWR
* net 11 VPB
* device instance $1 r0 *1 3.21,1.985 pfet_01v8_hvt
M$1 5 4 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $2 r0 *1 1.415,1.985 pfet_01v8_hvt
M$2 10 3 4 11 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=135000000000P PS=2530000U PD=1270000U
* device instance $3 r0 *1 1.835,1.985 pfet_01v8_hvt
M$3 9 6 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=140000000000P PS=1270000U PD=1280000U
* device instance $4 r0 *1 2.265,1.985 pfet_01v8_hvt
M$4 10 7 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=265000000000P PS=1280000U PD=2530000U
* device instance $5 r0 *1 0.47,2.275 pfet_01v8_hvt
M$5 9 2 3 11 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=109200000000P PS=1360000U PD=1360000U
* device instance $6 r0 *1 0.815,0.445 nfet_01v8
M$6 1 2 3 12 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=135900000000P
+ PS=1370000U PD=1100000U
* device instance $7 r0 *1 1.415,0.56 nfet_01v8
M$7 4 3 1 12 nfet_01v8 L=150000U W=650000U AS=135900000000P AD=87750000000P
+ PS=1100000U PD=920000U
* device instance $8 r0 *1 1.835,0.56 nfet_01v8
M$8 8 6 4 12 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=91000000000P
+ PS=920000U PD=930000U
* device instance $9 r0 *1 2.265,0.56 nfet_01v8
M$9 1 7 8 12 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=258375000000P
+ PS=930000U PD=1445000U
* device instance $10 r0 *1 3.21,0.56 nfet_01v8
M$10 5 4 1 12 nfet_01v8 L=150000U W=650000U AS=258375000000P AD=169000000000P
+ PS=1445000U PD=1820000U
.ENDS sky130_fd_sc_hd__a21bo_1

* cell sky130_fd_sc_hd__fa_2
* pin VGND
* pin COUT
* pin CIN
* pin SUM
* pin A
* pin B
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__fa_2 1 2 6 8 12 13 14 15 21
* net 1 VGND
* net 2 COUT
* net 6 CIN
* net 8 SUM
* net 12 A
* net 13 B
* net 14 VPWR
* net 15 VPB
* device instance $1 r0 *1 4.07,2.165 pfet_01v8_hvt
M$1 17 13 14 15 pfet_01v8_hvt L=150000U W=640000U AS=166400000000P
+ AD=86400000000P PS=1800000U PD=910000U
* device instance $2 r0 *1 4.49,2.165 pfet_01v8_hvt
M$2 14 6 17 15 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=86400000000P PS=910000U PD=910000U
* device instance $3 r0 *1 4.91,2.165 pfet_01v8_hvt
M$3 17 12 14 15 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=94400000000P PS=910000U PD=935000U
* device instance $4 r0 *1 5.355,2.165 pfet_01v8_hvt
M$4 7 3 17 15 pfet_01v8_hvt L=150000U W=640000U AS=94400000000P AD=88000000000P
+ PS=935000U PD=915000U
* device instance $5 r0 *1 5.78,2.165 pfet_01v8_hvt
M$5 19 6 7 15 pfet_01v8_hvt L=150000U W=640000U AS=88000000000P
+ AD=103625000000P PS=915000U PD=965000U
* device instance $6 r0 *1 6.255,2.17 pfet_01v8_hvt
M$6 20 13 19 15 pfet_01v8_hvt L=150000U W=630000U AS=103625000000P
+ AD=122850000000P PS=965000U PD=1020000U
* device instance $7 r0 *1 6.795,2.17 pfet_01v8_hvt
M$7 20 12 14 15 pfet_01v8_hvt L=150000U W=630000U AS=148625000000P
+ AD=122850000000P PS=1325000U PD=1020000U
* device instance $8 r0 *1 7.27,1.985 pfet_01v8_hvt
M$8 8 7 14 15 pfet_01v8_hvt L=150000U W=2000000U AS=283625000000P
+ AD=395000000000P PS=2595000U PD=3790000U
* device instance $10 r0 *1 0.475,1.985 pfet_01v8_hvt
M$10 2 3 14 15 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=283625000000P PS=3790000U PD=2595000U
* device instance $12 r0 *1 1.37,2.17 pfet_01v8_hvt
M$12 18 12 14 15 pfet_01v8_hvt L=150000U W=630000U AS=148625000000P
+ AD=92925000000P PS=1325000U PD=925000U
* device instance $13 r0 *1 1.815,2.17 pfet_01v8_hvt
M$13 3 13 18 15 pfet_01v8_hvt L=150000U W=630000U AS=92925000000P
+ AD=102375000000P PS=925000U PD=955000U
* device instance $14 r0 *1 2.29,2.17 pfet_01v8_hvt
M$14 16 6 3 15 pfet_01v8_hvt L=150000U W=630000U AS=102375000000P
+ AD=85050000000P PS=955000U PD=900000U
* device instance $15 r0 *1 2.71,2.17 pfet_01v8_hvt
M$15 14 12 16 15 pfet_01v8_hvt L=150000U W=630000U AS=85050000000P
+ AD=85050000000P PS=900000U PD=900000U
* device instance $16 r0 *1 3.13,2.17 pfet_01v8_hvt
M$16 16 13 14 15 pfet_01v8_hvt L=150000U W=630000U AS=85050000000P
+ AD=163800000000P PS=900000U PD=1780000U
* device instance $17 r0 *1 1.395,0.445 nfet_01v8
M$17 9 12 1 21 nfet_01v8 L=150000U W=420000U AS=103400000000P AD=68250000000P
+ PS=1000000U PD=745000U
* device instance $18 r0 *1 1.87,0.445 nfet_01v8
M$18 3 13 9 21 nfet_01v8 L=150000U W=420000U AS=68250000000P AD=56700000000P
+ PS=745000U PD=690000U
* device instance $19 r0 *1 2.29,0.445 nfet_01v8
M$19 4 6 3 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $20 r0 *1 2.71,0.445 nfet_01v8
M$20 1 12 4 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $21 r0 *1 3.13,0.445 nfet_01v8
M$21 4 13 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $22 r0 *1 0.475,0.56 nfet_01v8
M$22 2 3 1 21 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=191150000000P
+ PS=2740000U PD=1920000U
* device instance $24 r0 *1 4.07,0.445 nfet_01v8
M$24 5 13 1 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $25 r0 *1 4.49,0.445 nfet_01v8
M$25 1 6 5 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $26 r0 *1 4.91,0.445 nfet_01v8
M$26 5 12 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=61950000000P
+ PS=690000U PD=715000U
* device instance $27 r0 *1 5.355,0.445 nfet_01v8
M$27 7 3 5 21 nfet_01v8 L=150000U W=420000U AS=61950000000P AD=81900000000P
+ PS=715000U PD=810000U
* device instance $28 r0 *1 5.895,0.445 nfet_01v8
M$28 10 6 7 21 nfet_01v8 L=150000U W=420000U AS=81900000000P AD=44100000000P
+ PS=810000U PD=630000U
* device instance $29 r0 *1 6.255,0.445 nfet_01v8
M$29 11 13 10 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $30 r0 *1 6.735,0.445 nfet_01v8
M$30 1 12 11 21 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=102350000000P
+ PS=750000U PD=995000U
* device instance $31 r0 *1 7.23,0.56 nfet_01v8
M$31 8 7 1 21 nfet_01v8 L=150000U W=1300000U AS=229100000000P AD=295750000000P
+ PS=2035000U PD=2860000U
.ENDS sky130_fd_sc_hd__fa_2

* cell sky130_fd_sc_hd__dfrtp_4
* pin VGND
* pin RESET_B
* pin Q
* pin CLK
* pin D
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__dfrtp_4 1 6 9 14 15 17 18 21
* net 1 VGND
* net 6 RESET_B
* net 9 Q
* net 14 CLK
* net 15 D
* net 17 VPB
* net 18 VPWR
* device instance $1 r0 *1 8.63,1.985 pfet_01v8_hvt
M$1 9 8 18 17 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=710000000000P PS=6330000U PD=6420000U
* device instance $5 r0 *1 0.47,2.135 pfet_01v8_hvt
M$5 18 14 2 17 pfet_01v8_hvt L=150000U W=640000U AS=166400000000P
+ AD=86400000000P PS=1800000U PD=910000U
* device instance $6 r0 *1 0.89,2.135 pfet_01v8_hvt
M$6 3 2 18 17 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=166400000000P PS=910000U PD=1800000U
* device instance $7 r0 *1 5.35,2.065 pfet_01v8_hvt
M$7 16 5 18 17 pfet_01v8_hvt L=150000U W=840000U AS=218400000000P
+ AD=129150000000P PS=2200000U PD=1185000U
* device instance $8 r0 *1 5.845,2.275 pfet_01v8_hvt
M$8 7 2 16 17 pfet_01v8_hvt L=150000U W=420000U AS=129150000000P
+ AD=58800000000P PS=1185000U PD=700000U
* device instance $9 r0 *1 6.275,2.275 pfet_01v8_hvt
M$9 20 3 7 17 pfet_01v8_hvt L=150000U W=420000U AS=58800000000P AD=56700000000P
+ PS=700000U PD=690000U
* device instance $10 r0 *1 6.695,2.275 pfet_01v8_hvt
M$10 18 8 20 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=81900000000P PS=690000U PD=810000U
* device instance $11 r0 *1 7.235,2.275 pfet_01v8_hvt
M$11 8 6 18 17 pfet_01v8_hvt L=150000U W=420000U AS=81900000000P
+ AD=56700000000P PS=810000U PD=690000U
* device instance $12 r0 *1 7.655,2.275 pfet_01v8_hvt
M$12 18 7 8 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=113400000000P PS=690000U PD=1380000U
* device instance $13 r0 *1 2.225,2.275 pfet_01v8_hvt
M$13 4 15 18 17 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=65100000000P PS=1360000U PD=730000U
* device instance $14 r0 *1 2.685,2.275 pfet_01v8_hvt
M$14 5 3 4 17 pfet_01v8_hvt L=150000U W=420000U AS=65100000000P AD=72450000000P
+ PS=730000U PD=765000U
* device instance $15 r0 *1 3.18,2.275 pfet_01v8_hvt
M$15 19 2 5 17 pfet_01v8_hvt L=150000U W=420000U AS=72450000000P
+ AD=115500000000P PS=765000U PD=970000U
* device instance $16 r0 *1 3.88,2.275 pfet_01v8_hvt
M$16 18 16 19 17 pfet_01v8_hvt L=150000U W=420000U AS=115500000000P
+ AD=70350000000P PS=970000U PD=755000U
* device instance $17 r0 *1 4.365,2.275 pfet_01v8_hvt
M$17 19 6 18 17 pfet_01v8_hvt L=150000U W=420000U AS=70350000000P
+ AD=109200000000P PS=755000U PD=1360000U
* device instance $18 r0 *1 8.63,0.56 nfet_01v8
M$18 9 8 1 21 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=445250000000P
+ PS=4580000U PD=4620000U
* device instance $22 r0 *1 0.47,0.445 nfet_01v8
M$22 1 14 2 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $23 r0 *1 0.89,0.445 nfet_01v8
M$23 3 2 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $24 r0 *1 2.64,0.415 nfet_01v8
M$24 5 2 4 21 nfet_01v8 L=150000U W=360000U AS=66000000000P AD=59400000000P
+ PS=745000U PD=690000U
* device instance $25 r0 *1 3.12,0.415 nfet_01v8
M$25 10 3 5 21 nfet_01v8 L=150000U W=360000U AS=59400000000P AD=140100000000P
+ PS=690000U PD=1100000U
* device instance $26 r0 *1 5.465,0.415 nfet_01v8
M$26 7 3 16 21 nfet_01v8 L=150000U W=360000U AS=99900000000P AD=71100000000P
+ PS=985000U PD=755000U
* device instance $27 r0 *1 6.01,0.415 nfet_01v8
M$27 13 2 7 21 nfet_01v8 L=150000U W=360000U AS=71100000000P AD=66900000000P
+ PS=755000U PD=750000U
* device instance $28 r0 *1 2.165,0.445 nfet_01v8
M$28 4 15 1 21 nfet_01v8 L=150000U W=420000U AS=220500000000P AD=66000000000P
+ PS=1890000U PD=745000U
* device instance $29 r0 *1 3.95,0.445 nfet_01v8
M$29 11 16 10 21 nfet_01v8 L=150000U W=420000U AS=140100000000P AD=44100000000P
+ PS=1100000U PD=630000U
* device instance $30 r0 *1 4.31,0.445 nfet_01v8
M$30 1 6 11 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=134600000000P
+ PS=630000U PD=1150000U
* device instance $31 r0 *1 6.49,0.445 nfet_01v8
M$31 1 8 13 21 nfet_01v8 L=150000U W=420000U AS=66900000000P AD=124950000000P
+ PS=750000U PD=1015000U
* device instance $32 r0 *1 7.235,0.445 nfet_01v8
M$32 12 6 1 21 nfet_01v8 L=150000U W=420000U AS=124950000000P AD=64050000000P
+ PS=1015000U PD=725000U
* device instance $33 r0 *1 7.69,0.445 nfet_01v8
M$33 8 7 12 21 nfet_01v8 L=150000U W=420000U AS=64050000000P AD=109200000000P
+ PS=725000U PD=1360000U
* device instance $34 r0 *1 4.97,0.555 nfet_01v8
M$34 16 5 1 21 nfet_01v8 L=150000U W=640000U AS=134600000000P AD=99900000000P
+ PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_4

* cell sky130_fd_sc_hd__dfrtp_1
* pin VGND
* pin RESET_B
* pin Q
* pin CLK
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__dfrtp_1 1 6 9 14 15 17 18 21
* net 1 VGND
* net 6 RESET_B
* net 9 Q
* net 14 CLK
* net 15 D
* net 17 VPWR
* net 18 VPB
* device instance $1 r0 *1 8.73,1.985 pfet_01v8_hvt
M$1 9 8 17 18 pfet_01v8_hvt L=150000U W=1000000U AS=301200000000P
+ AD=260000000000P PS=2660000U PD=2520000U
* device instance $2 r0 *1 0.47,2.135 pfet_01v8_hvt
M$2 17 14 2 18 pfet_01v8_hvt L=150000U W=640000U AS=166400000000P
+ AD=86400000000P PS=1800000U PD=910000U
* device instance $3 r0 *1 0.89,2.135 pfet_01v8_hvt
M$3 3 2 17 18 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=166400000000P PS=910000U PD=1800000U
* device instance $4 r0 *1 5.35,2.065 pfet_01v8_hvt
M$4 16 5 17 18 pfet_01v8_hvt L=150000U W=840000U AS=218400000000P
+ AD=129150000000P PS=2200000U PD=1185000U
* device instance $5 r0 *1 5.845,2.275 pfet_01v8_hvt
M$5 7 2 16 18 pfet_01v8_hvt L=150000U W=420000U AS=129150000000P
+ AD=58800000000P PS=1185000U PD=700000U
* device instance $6 r0 *1 6.275,2.275 pfet_01v8_hvt
M$6 20 3 7 18 pfet_01v8_hvt L=150000U W=420000U AS=58800000000P AD=56700000000P
+ PS=700000U PD=690000U
* device instance $7 r0 *1 6.695,2.275 pfet_01v8_hvt
M$7 17 8 20 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=81900000000P PS=690000U PD=810000U
* device instance $8 r0 *1 7.235,2.275 pfet_01v8_hvt
M$8 8 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=81900000000P AD=56700000000P
+ PS=810000U PD=690000U
* device instance $9 r0 *1 7.655,2.275 pfet_01v8_hvt
M$9 17 7 8 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=113400000000P PS=690000U PD=1380000U
* device instance $10 r0 *1 2.225,2.275 pfet_01v8_hvt
M$10 4 15 17 18 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=65100000000P PS=1360000U PD=730000U
* device instance $11 r0 *1 2.685,2.275 pfet_01v8_hvt
M$11 5 3 4 18 pfet_01v8_hvt L=150000U W=420000U AS=65100000000P AD=72450000000P
+ PS=730000U PD=765000U
* device instance $12 r0 *1 3.18,2.275 pfet_01v8_hvt
M$12 19 2 5 18 pfet_01v8_hvt L=150000U W=420000U AS=72450000000P
+ AD=115500000000P PS=765000U PD=970000U
* device instance $13 r0 *1 3.88,2.275 pfet_01v8_hvt
M$13 17 16 19 18 pfet_01v8_hvt L=150000U W=420000U AS=115500000000P
+ AD=70350000000P PS=970000U PD=755000U
* device instance $14 r0 *1 4.365,2.275 pfet_01v8_hvt
M$14 19 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=70350000000P
+ AD=109200000000P PS=755000U PD=1360000U
* device instance $15 r0 *1 8.73,0.56 nfet_01v8
M$15 9 8 1 21 nfet_01v8 L=150000U W=650000U AS=208700000000P AD=169000000000P
+ PS=2020000U PD=1820000U
* device instance $16 r0 *1 0.47,0.445 nfet_01v8
M$16 1 14 2 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $17 r0 *1 0.89,0.445 nfet_01v8
M$17 3 2 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $18 r0 *1 2.64,0.415 nfet_01v8
M$18 5 2 4 21 nfet_01v8 L=150000U W=360000U AS=66000000000P AD=59400000000P
+ PS=745000U PD=690000U
* device instance $19 r0 *1 3.12,0.415 nfet_01v8
M$19 12 3 5 21 nfet_01v8 L=150000U W=360000U AS=59400000000P AD=140100000000P
+ PS=690000U PD=1100000U
* device instance $20 r0 *1 5.465,0.415 nfet_01v8
M$20 7 3 16 21 nfet_01v8 L=150000U W=360000U AS=99900000000P AD=71100000000P
+ PS=985000U PD=755000U
* device instance $21 r0 *1 6.01,0.415 nfet_01v8
M$21 11 2 7 21 nfet_01v8 L=150000U W=360000U AS=71100000000P AD=66900000000P
+ PS=755000U PD=750000U
* device instance $22 r0 *1 2.165,0.445 nfet_01v8
M$22 4 15 1 21 nfet_01v8 L=150000U W=420000U AS=220500000000P AD=66000000000P
+ PS=1890000U PD=745000U
* device instance $23 r0 *1 3.95,0.445 nfet_01v8
M$23 13 16 12 21 nfet_01v8 L=150000U W=420000U AS=140100000000P AD=44100000000P
+ PS=1100000U PD=630000U
* device instance $24 r0 *1 4.31,0.445 nfet_01v8
M$24 1 6 13 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=134600000000P
+ PS=630000U PD=1150000U
* device instance $25 r0 *1 6.49,0.445 nfet_01v8
M$25 1 8 11 21 nfet_01v8 L=150000U W=420000U AS=66900000000P AD=124950000000P
+ PS=750000U PD=1015000U
* device instance $26 r0 *1 7.235,0.445 nfet_01v8
M$26 10 6 1 21 nfet_01v8 L=150000U W=420000U AS=124950000000P AD=64050000000P
+ PS=1015000U PD=725000U
* device instance $27 r0 *1 7.69,0.445 nfet_01v8
M$27 8 7 10 21 nfet_01v8 L=150000U W=420000U AS=64050000000P AD=109200000000P
+ PS=725000U PD=1360000U
* device instance $28 r0 *1 4.97,0.555 nfet_01v8
M$28 16 5 1 21 nfet_01v8 L=150000U W=640000U AS=134600000000P AD=99900000000P
+ PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_1

* cell sky130_fd_sc_hd__clkbuf_1
* pin VPB
* pin A
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_1 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 X
* net 5 VGND
* net 6 VPWR
* device instance $1 r0 *1 0.47,2.09 pfet_01v8_hvt
M$1 6 2 4 1 pfet_01v8_hvt L=150000U W=790000U AS=205400000000P AD=114550000000P
+ PS=2100000U PD=1080000U
* device instance $2 r0 *1 0.91,2.09 pfet_01v8_hvt
M$2 2 3 6 1 pfet_01v8_hvt L=150000U W=790000U AS=114550000000P AD=205400000000P
+ PS=1080000U PD=2100000U
* device instance $3 r0 *1 0.47,0.495 nfet_01v8
M$3 5 2 4 7 nfet_01v8 L=150000U W=520000U AS=135200000000P AD=75400000000P
+ PS=1560000U PD=810000U
* device instance $4 r0 *1 0.91,0.495 nfet_01v8
M$4 2 3 5 7 nfet_01v8 L=150000U W=520000U AS=75400000000P AD=135200000000P
+ PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

* cell sky130_fd_sc_hd__dfrtp_2
* pin VGND
* pin RESET_B
* pin Q
* pin CLK
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__dfrtp_2 1 6 9 14 15 17 18 21
* net 1 VGND
* net 6 RESET_B
* net 9 Q
* net 14 CLK
* net 15 D
* net 17 VPWR
* net 18 VPB
* device instance $1 r0 *1 8.73,1.985 pfet_01v8_hvt
M$1 9 8 17 18 pfet_01v8_hvt L=150000U W=2000000U AS=436200000000P
+ AD=395000000000P PS=3930000U PD=3790000U
* device instance $3 r0 *1 0.47,2.135 pfet_01v8_hvt
M$3 17 14 2 18 pfet_01v8_hvt L=150000U W=640000U AS=166400000000P
+ AD=86400000000P PS=1800000U PD=910000U
* device instance $4 r0 *1 0.89,2.135 pfet_01v8_hvt
M$4 3 2 17 18 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=166400000000P PS=910000U PD=1800000U
* device instance $5 r0 *1 5.35,2.065 pfet_01v8_hvt
M$5 16 5 17 18 pfet_01v8_hvt L=150000U W=840000U AS=218400000000P
+ AD=129150000000P PS=2200000U PD=1185000U
* device instance $6 r0 *1 5.845,2.275 pfet_01v8_hvt
M$6 7 2 16 18 pfet_01v8_hvt L=150000U W=420000U AS=129150000000P
+ AD=58800000000P PS=1185000U PD=700000U
* device instance $7 r0 *1 6.275,2.275 pfet_01v8_hvt
M$7 20 3 7 18 pfet_01v8_hvt L=150000U W=420000U AS=58800000000P AD=56700000000P
+ PS=700000U PD=690000U
* device instance $8 r0 *1 6.695,2.275 pfet_01v8_hvt
M$8 17 8 20 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=81900000000P PS=690000U PD=810000U
* device instance $9 r0 *1 7.235,2.275 pfet_01v8_hvt
M$9 8 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=81900000000P AD=56700000000P
+ PS=810000U PD=690000U
* device instance $10 r0 *1 7.655,2.275 pfet_01v8_hvt
M$10 17 7 8 18 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=113400000000P PS=690000U PD=1380000U
* device instance $11 r0 *1 2.225,2.275 pfet_01v8_hvt
M$11 4 15 17 18 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=65100000000P PS=1360000U PD=730000U
* device instance $12 r0 *1 2.685,2.275 pfet_01v8_hvt
M$12 5 3 4 18 pfet_01v8_hvt L=150000U W=420000U AS=65100000000P AD=72450000000P
+ PS=730000U PD=765000U
* device instance $13 r0 *1 3.18,2.275 pfet_01v8_hvt
M$13 19 2 5 18 pfet_01v8_hvt L=150000U W=420000U AS=72450000000P
+ AD=115500000000P PS=765000U PD=970000U
* device instance $14 r0 *1 3.88,2.275 pfet_01v8_hvt
M$14 17 16 19 18 pfet_01v8_hvt L=150000U W=420000U AS=115500000000P
+ AD=70350000000P PS=970000U PD=755000U
* device instance $15 r0 *1 4.365,2.275 pfet_01v8_hvt
M$15 19 6 17 18 pfet_01v8_hvt L=150000U W=420000U AS=70350000000P
+ AD=109200000000P PS=755000U PD=1360000U
* device instance $16 r0 *1 8.73,0.56 nfet_01v8
M$16 9 8 1 21 nfet_01v8 L=150000U W=1300000U AS=296450000000P AD=256750000000P
+ PS=2940000U PD=2740000U
* device instance $18 r0 *1 0.47,0.445 nfet_01v8
M$18 1 14 2 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $19 r0 *1 0.89,0.445 nfet_01v8
M$19 3 2 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $20 r0 *1 2.64,0.415 nfet_01v8
M$20 5 2 4 21 nfet_01v8 L=150000U W=360000U AS=66000000000P AD=59400000000P
+ PS=745000U PD=690000U
* device instance $21 r0 *1 3.12,0.415 nfet_01v8
M$21 11 3 5 21 nfet_01v8 L=150000U W=360000U AS=59400000000P AD=140100000000P
+ PS=690000U PD=1100000U
* device instance $22 r0 *1 5.465,0.415 nfet_01v8
M$22 7 3 16 21 nfet_01v8 L=150000U W=360000U AS=99900000000P AD=71100000000P
+ PS=985000U PD=755000U
* device instance $23 r0 *1 6.01,0.415 nfet_01v8
M$23 12 2 7 21 nfet_01v8 L=150000U W=360000U AS=71100000000P AD=66900000000P
+ PS=755000U PD=750000U
* device instance $24 r0 *1 2.165,0.445 nfet_01v8
M$24 4 15 1 21 nfet_01v8 L=150000U W=420000U AS=220500000000P AD=66000000000P
+ PS=1890000U PD=745000U
* device instance $25 r0 *1 3.95,0.445 nfet_01v8
M$25 13 16 11 21 nfet_01v8 L=150000U W=420000U AS=140100000000P AD=44100000000P
+ PS=1100000U PD=630000U
* device instance $26 r0 *1 4.31,0.445 nfet_01v8
M$26 1 6 13 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=134600000000P
+ PS=630000U PD=1150000U
* device instance $27 r0 *1 6.49,0.445 nfet_01v8
M$27 1 8 12 21 nfet_01v8 L=150000U W=420000U AS=66900000000P AD=124950000000P
+ PS=750000U PD=1015000U
* device instance $28 r0 *1 7.235,0.445 nfet_01v8
M$28 10 6 1 21 nfet_01v8 L=150000U W=420000U AS=124950000000P AD=64050000000P
+ PS=1015000U PD=725000U
* device instance $29 r0 *1 7.69,0.445 nfet_01v8
M$29 8 7 10 21 nfet_01v8 L=150000U W=420000U AS=64050000000P AD=109200000000P
+ PS=725000U PD=1360000U
* device instance $30 r0 *1 4.97,0.555 nfet_01v8
M$30 16 5 1 21 nfet_01v8 L=150000U W=640000U AS=134600000000P AD=99900000000P
+ PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_2

* cell sky130_fd_sc_hd__ha_2
* pin VGND
* pin SUM
* pin COUT
* pin B
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__ha_2 1 2 6 7 8 10 11 13
* net 1 VGND
* net 2 SUM
* net 6 COUT
* net 7 B
* net 8 A
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 2 3 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=446600000000P PS=3830000U PD=3075000U
* device instance $3 r0 *1 1.845,2.165 pfet_01v8_hvt
M$3 3 5 10 11 pfet_01v8_hvt L=150000U W=640000U AS=291600000000P
+ AD=86400000000P PS=1765000U PD=910000U
* device instance $4 r0 *1 2.265,2.165 pfet_01v8_hvt
M$4 12 7 3 11 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=128000000000P PS=910000U PD=1040000U
* device instance $5 r0 *1 2.815,2.165 pfet_01v8_hvt
M$5 10 8 12 11 pfet_01v8_hvt L=150000U W=640000U AS=128000000000P
+ AD=227200000000P PS=1040000U PD=1350000U
* device instance $6 r0 *1 3.675,2.165 pfet_01v8_hvt
M$6 5 7 10 11 pfet_01v8_hvt L=150000U W=640000U AS=227200000000P
+ AD=92800000000P PS=1350000U PD=930000U
* device instance $7 r0 *1 4.115,2.165 pfet_01v8_hvt
M$7 5 8 10 11 pfet_01v8_hvt L=150000U W=640000U AS=149000000000P
+ AD=92800000000P PS=1325000U PD=930000U
* device instance $8 r0 *1 4.59,1.985 pfet_01v8_hvt
M$8 6 5 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=304000000000P
+ AD=415000000000P PS=2635000U PD=3830000U
* device instance $10 r0 *1 3.755,0.445 nfet_01v8
M$10 9 7 5 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $11 r0 *1 4.115,0.445 nfet_01v8
M$11 1 8 9 13 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=97000000000P
+ PS=630000U PD=975000U
* device instance $12 r0 *1 4.59,0.56 nfet_01v8
M$12 6 5 1 13 nfet_01v8 L=150000U W=1300000U AS=197750000000P AD=269750000000P
+ PS=1935000U PD=2780000U
* device instance $14 r0 *1 0.47,0.56 nfet_01v8
M$14 2 3 1 13 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=269750000000P
+ PS=2780000U PD=2780000U
* device instance $16 r0 *1 1.87,0.445 nfet_01v8
M$16 4 5 3 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $17 r0 *1 2.29,0.445 nfet_01v8
M$17 1 7 4 13 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $18 r0 *1 2.71,0.445 nfet_01v8
M$18 4 8 1 13 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__ha_2

* cell sky130_fd_sc_hd__o311ai_0
* pin VGND
* pin A1
* pin Y
* pin C1
* pin A2
* pin A3
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311ai_0 1 2 4 5 7 8 9 10 11 14
* net 1 VGND
* net 2 A1
* net 4 Y
* net 5 C1
* net 7 A2
* net 8 A3
* net 9 B1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.615,2.165 pfet_01v8_hvt
M$1 12 2 10 11 pfet_01v8_hvt L=150000U W=640000U AS=179200000000P
+ AD=86400000000P PS=1840000U PD=910000U
* device instance $2 r0 *1 1.035,2.165 pfet_01v8_hvt
M$2 13 7 12 11 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=86400000000P PS=910000U PD=910000U
* device instance $3 r0 *1 1.455,2.165 pfet_01v8_hvt
M$3 4 8 13 11 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=144000000000P PS=910000U PD=1090000U
* device instance $4 r0 *1 2.055,2.165 pfet_01v8_hvt
M$4 10 9 4 11 pfet_01v8_hvt L=150000U W=640000U AS=144000000000P
+ AD=118400000000P PS=1090000U PD=1010000U
* device instance $5 r0 *1 2.575,2.165 pfet_01v8_hvt
M$5 4 5 10 11 pfet_01v8_hvt L=150000U W=640000U AS=118400000000P
+ AD=198400000000P PS=1010000U PD=1900000U
* device instance $6 r0 *1 0.615,0.445 nfet_01v8
M$6 3 2 1 14 nfet_01v8 L=150000U W=420000U AS=117600000000P AD=56700000000P
+ PS=1400000U PD=690000U
* device instance $7 r0 *1 1.035,0.445 nfet_01v8
M$7 1 7 3 14 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $8 r0 *1 1.455,0.445 nfet_01v8
M$8 3 8 1 14 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=128100000000P
+ PS=690000U PD=1030000U
* device instance $9 r0 *1 2.215,0.445 nfet_01v8
M$9 6 9 3 14 nfet_01v8 L=150000U W=420000U AS=128100000000P AD=44100000000P
+ PS=1030000U PD=630000U
* device instance $10 r0 *1 2.575,0.445 nfet_01v8
M$10 4 5 6 14 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=117600000000P
+ PS=630000U PD=1400000U
.ENDS sky130_fd_sc_hd__o311ai_0

* cell sky130_fd_sc_hd__o311a_2
* pin VGND
* pin X
* pin A1
* pin A2
* pin A3
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311a_2 1 2 5 6 7 8 9 11 12 15
* net 1 VGND
* net 2 X
* net 5 A1
* net 6 A2
* net 7 A3
* net 8 B1
* net 9 C1
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.53,1.985 pfet_01v8_hvt
M$1 2 4 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=455000000000P
+ AD=447500000000P PS=3910000U PD=2895000U
* device instance $3 r0 *1 1.725,1.985 pfet_01v8_hvt
M$3 13 5 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=312500000000P
+ AD=175000000000P PS=1625000U PD=1350000U
* device instance $4 r0 *1 2.225,1.985 pfet_01v8_hvt
M$4 14 6 13 12 pfet_01v8_hvt L=150000U W=1000000U AS=175000000000P
+ AD=210000000000P PS=1350000U PD=1420000U
* device instance $5 r0 *1 2.795,1.985 pfet_01v8_hvt
M$5 4 7 14 12 pfet_01v8_hvt L=150000U W=1000000U AS=210000000000P
+ AD=137500000000P PS=1420000U PD=1275000U
* device instance $6 r0 *1 3.22,1.985 pfet_01v8_hvt
M$6 11 8 4 12 pfet_01v8_hvt L=150000U W=1000000U AS=137500000000P
+ AD=150000000000P PS=1275000U PD=1300000U
* device instance $7 r0 *1 3.67,1.985 pfet_01v8_hvt
M$7 4 9 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=150000000000P
+ AD=260000000000P PS=1300000U PD=2520000U
* device instance $8 r0 *1 0.53,0.56 nfet_01v8
M$8 2 4 1 15 nfet_01v8 L=150000U W=1300000U AS=295750000000P AD=290875000000P
+ PS=2860000U PD=2195000U
* device instance $10 r0 *1 1.725,0.56 nfet_01v8
M$10 3 5 1 15 nfet_01v8 L=150000U W=650000U AS=203125000000P AD=113750000000P
+ PS=1275000U PD=1000000U
* device instance $11 r0 *1 2.225,0.56 nfet_01v8
M$11 1 6 3 15 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=136500000000P
+ PS=1000000U PD=1070000U
* device instance $12 r0 *1 2.795,0.56 nfet_01v8
M$12 3 7 1 15 nfet_01v8 L=150000U W=650000U AS=136500000000P AD=118625000000P
+ PS=1070000U PD=1015000U
* device instance $13 r0 *1 3.31,0.56 nfet_01v8
M$13 10 8 3 15 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=68250000000P
+ PS=1015000U PD=860000U
* device instance $14 r0 *1 3.67,0.56 nfet_01v8
M$14 4 9 10 15 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=169000000000P
+ PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o311a_2

* cell sky130_fd_sc_hd__a311oi_2
* pin VGND
* pin Y
* pin A3
* pin A2
* pin A1
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a311oi_2 1 4 5 6 7 8 9 10 13 14
* net 1 VGND
* net 4 Y
* net 5 A3
* net 6 A2
* net 7 A1
* net 8 B1
* net 9 C1
* net 10 VPWR
* net 13 VPB
* device instance $1 r0 *1 3.54,1.985 pfet_01v8_hvt
M$1 11 8 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=2790000U
* device instance $3 r0 *1 4.63,1.985 pfet_01v8_hvt
M$3 4 9 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=2790000U PD=3790000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 11 5 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $7 r0 *1 1.31,1.985 pfet_01v8_hvt
M$7 11 6 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=275000000000P
+ AD=285000000000P PS=2550000U PD=2570000U
* device instance $9 r0 *1 2.18,1.985 pfet_01v8_hvt
M$9 11 7 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=395000000000P PS=2560000U PD=3790000U
* device instance $11 r0 *1 2.67,0.56 nfet_01v8
M$11 3 7 4 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=185250000000P
+ PS=2740000U PD=1870000U
* device instance $13 r0 *1 3.54,0.56 nfet_01v8
M$13 1 8 4 14 nfet_01v8 L=150000U W=1300000U AS=185250000000P AD=256750000000P
+ PS=1870000U PD=2090000U
* device instance $15 r0 *1 4.63,0.56 nfet_01v8
M$15 1 9 4 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2090000U PD=2740000U
* device instance $17 r0 *1 0.47,0.56 nfet_01v8
M$17 1 5 2 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $19 r0 *1 1.31,0.56 nfet_01v8
M$19 3 6 2 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__a311oi_2

* cell sky130_fd_sc_hd__or3b_1
* pin VPB
* pin A
* pin B
* pin C_N
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__or3b_1 1 2 3 5 6 7 8 10
* net 1 VPB
* net 2 A
* net 3 B
* net 5 C_N
* net 6 X
* net 7 VPWR
* net 8 VGND
* device instance $1 r0 *1 1.41,1.695 pfet_01v8_hvt
M$1 11 4 9 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 1.77,1.695 pfet_01v8_hvt
M$2 12 3 11 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=68250000000P
+ PS=630000U PD=745000U
* device instance $3 r0 *1 2.245,1.695 pfet_01v8_hvt
M$3 7 2 12 1 pfet_01v8_hvt L=150000U W=420000U AS=68250000000P AD=148250000000P
+ PS=745000U PD=1340000U
* device instance $4 r0 *1 2.735,1.985 pfet_01v8_hvt
M$4 6 9 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=148250000000P
+ AD=275000000000P PS=1340000U PD=2550000U
* device instance $5 r0 *1 0.47,1.695 pfet_01v8_hvt
M$5 4 5 7 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $6 r0 *1 1.41,0.475 nfet_01v8
M$6 8 4 9 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $7 r0 *1 1.83,0.475 nfet_01v8
M$7 9 3 8 10 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $8 r0 *1 2.25,0.475 nfet_01v8
M$8 9 2 8 10 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=56700000000P
+ PS=985000U PD=690000U
* device instance $9 r0 *1 2.735,0.56 nfet_01v8
M$9 6 9 8 10 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=178750000000P
+ PS=985000U PD=1850000U
* device instance $10 r0 *1 0.47,0.675 nfet_01v8
M$10 4 5 8 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__or3b_1

* cell sky130_fd_sc_hd__and3_4
* pin VGND
* pin B
* pin X
* pin A
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__and3_4 1 3 4 5 6 9 10 11
* net 1 VGND
* net 3 B
* net 4 X
* net 5 A
* net 6 C
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.85,1.985 pfet_01v8_hvt
M$1 9 5 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=305000000000P
+ AD=197500000000P PS=2610000U PD=1395000U
* device instance $2 r0 *1 1.395,1.985 pfet_01v8_hvt
M$2 2 3 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=197500000000P
+ AD=140000000000P PS=1395000U PD=1280000U
* device instance $3 r0 *1 1.825,1.985 pfet_01v8_hvt
M$3 9 6 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=177500000000P PS=1280000U PD=1355000U
* device instance $4 r0 *1 2.33,1.985 pfet_01v8_hvt
M$4 4 2 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=597500000000P
+ AD=705000000000P PS=5195000U PD=6410000U
* device instance $8 r0 *1 0.85,0.56 nfet_01v8
M$8 8 5 2 11 nfet_01v8 L=150000U W=650000U AS=198250000000P AD=128375000000P
+ PS=1910000U PD=1045000U
* device instance $9 r0 *1 1.395,0.56 nfet_01v8
M$9 7 3 8 11 nfet_01v8 L=150000U W=650000U AS=128375000000P AD=68250000000P
+ PS=1045000U PD=860000U
* device instance $10 r0 *1 1.755,0.56 nfet_01v8
M$10 1 6 7 11 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=138125000000P
+ PS=860000U PD=1075000U
* device instance $11 r0 *1 2.33,0.56 nfet_01v8
M$11 4 2 1 11 nfet_01v8 L=150000U W=2600000U AS=411125000000P AD=458250000000P
+ PS=3865000U PD=4660000U
.ENDS sky130_fd_sc_hd__and3_4

* cell sky130_fd_sc_hd__o221ai_1
* pin VPB
* pin C1
* pin B1
* pin A2
* pin A1
* pin B2
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o221ai_1 1 2 3 4 5 6 8 10 11 12
* net 1 VPB
* net 2 C1
* net 3 B1
* net 4 A2
* net 5 A1
* net 6 B2
* net 8 Y
* net 10 VPWR
* net 11 VGND
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 10 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=380000000000P PS=2560000U PD=1760000U
* device instance $2 r0 *1 1.4,1.985 pfet_01v8_hvt
M$2 14 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=380000000000P
+ AD=120000000000P PS=1760000U PD=1240000U
* device instance $3 r0 *1 1.79,1.985 pfet_01v8_hvt
M$3 8 6 14 1 pfet_01v8_hvt L=150000U W=1000000U AS=120000000000P
+ AD=225000000000P PS=1240000U PD=1450000U
* device instance $4 r0 *1 2.39,1.985 pfet_01v8_hvt
M$4 13 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=225000000000P
+ AD=105000000000P PS=1450000U PD=1210000U
* device instance $5 r0 *1 2.75,1.985 pfet_01v8_hvt
M$5 10 5 13 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $6 r0 *1 1.4,0.56 nfet_01v8
M$6 9 3 7 12 nfet_01v8 L=150000U W=650000U AS=165200000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 1.82,0.56 nfet_01v8
M$7 7 6 9 12 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=117000000000P
+ PS=920000U PD=1010000U
* device instance $8 r0 *1 2.33,0.56 nfet_01v8
M$8 11 4 7 12 nfet_01v8 L=150000U W=650000U AS=117000000000P AD=87750000000P
+ PS=1010000U PD=920000U
* device instance $9 r0 *1 2.75,0.56 nfet_01v8
M$9 7 5 11 12 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $10 r0 *1 0.47,0.56 nfet_01v8
M$10 9 2 8 12 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=165400000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221ai_1

* cell sky130_fd_sc_hd__a32o_1
* pin VGND
* pin X
* pin A2
* pin A1
* pin B1
* pin A3
* pin B2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a32o_1 1 2 3 4 5 7 8 13 14 15
* net 1 VGND
* net 2 X
* net 3 A2
* net 4 A1
* net 5 B1
* net 7 A3
* net 8 B2
* net 13 VPWR
* net 14 VPB
* device instance $1 r0 *1 0.54,1.985 pfet_01v8_hvt
M$1 13 6 2 14 pfet_01v8_hvt L=150000U W=1000000U AS=330000000000P
+ AD=242500000000P PS=2660000U PD=1485000U
* device instance $2 r0 *1 1.175,1.985 pfet_01v8_hvt
M$2 12 7 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=242500000000P
+ AD=165000000000P PS=1485000U PD=1330000U
* device instance $3 r0 *1 1.655,1.985 pfet_01v8_hvt
M$3 13 3 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=225000000000P PS=1330000U PD=1450000U
* device instance $4 r0 *1 2.255,1.985 pfet_01v8_hvt
M$4 12 4 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=225000000000P
+ AD=185000000000P PS=1450000U PD=1370000U
* device instance $5 r0 *1 2.775,1.985 pfet_01v8_hvt
M$5 6 5 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=185000000000P
+ AD=140000000000P PS=1370000U PD=1280000U
* device instance $6 r0 *1 3.205,1.985 pfet_01v8_hvt
M$6 12 8 6 14 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=265000000000P PS=1280000U PD=2530000U
* device instance $7 r0 *1 0.54,0.56 nfet_01v8
M$7 1 6 2 15 nfet_01v8 L=150000U W=650000U AS=214500000000P AD=167375000000P
+ PS=1960000U PD=1165000U
* device instance $8 r0 *1 1.205,0.56 nfet_01v8
M$8 9 7 1 15 nfet_01v8 L=150000U W=650000U AS=167375000000P AD=97500000000P
+ PS=1165000U PD=950000U
* device instance $9 r0 *1 1.655,0.56 nfet_01v8
M$9 11 3 9 15 nfet_01v8 L=150000U W=650000U AS=97500000000P AD=146250000000P
+ PS=950000U PD=1100000U
* device instance $10 r0 *1 2.255,0.56 nfet_01v8
M$10 6 4 11 15 nfet_01v8 L=150000U W=650000U AS=146250000000P AD=143000000000P
+ PS=1100000U PD=1090000U
* device instance $11 r0 *1 2.845,0.56 nfet_01v8
M$11 10 5 6 15 nfet_01v8 L=150000U W=650000U AS=143000000000P AD=68250000000P
+ PS=1090000U PD=860000U
* device instance $12 r0 *1 3.205,0.56 nfet_01v8
M$12 1 8 10 15 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=172250000000P
+ PS=860000U PD=1830000U
.ENDS sky130_fd_sc_hd__a32o_1

* cell sky130_fd_sc_hd__nand2b_2
* pin VGND
* pin Y
* pin A_N
* pin B
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand2b_2 1 4 5 6 7 8 9
* net 1 VGND
* net 4 Y
* net 5 A_N
* net 6 B
* net 7 VPWR
* net 8 VPB
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 7 5 2 8 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=146800000000P
+ PS=1360000U PD=1340000U
* device instance $2 r0 *1 0.96,1.985 pfet_01v8_hvt
M$2 4 2 7 8 pfet_01v8_hvt L=150000U W=2000000U AS=311800000000P
+ AD=500000000000P PS=2670000U PD=3000000U
* device instance $4 r0 *1 2.26,1.985 pfet_01v8_hvt
M$4 4 6 7 8 pfet_01v8_hvt L=150000U W=2000000U AS=470000000000P
+ AD=410000000000P PS=2940000U PD=3820000U
* device instance $6 r0 *1 1.48,0.56 nfet_01v8
M$6 4 2 3 9 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $8 r0 *1 2.32,0.56 nfet_01v8
M$8 1 6 3 9 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $10 r0 *1 0.47,0.675 nfet_01v8
M$10 2 5 1 9 nfet_01v8 L=150000U W=420000U AS=194000000000P AD=109200000000P
+ PS=1950000U PD=1360000U
.ENDS sky130_fd_sc_hd__nand2b_2

* cell sky130_fd_sc_hd__a311oi_1
* pin VPB
* pin A3
* pin A2
* pin B1
* pin A1
* pin C1
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a311oi_1 1 2 3 4 5 6 7 9 10 11
* net 1 VPB
* net 2 A3
* net 3 A2
* net 4 B1
* net 5 A1
* net 6 C1
* net 7 VPWR
* net 9 Y
* net 10 VGND
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=137500000000P PS=2520000U PD=1275000U
* device instance $2 r0 *1 0.895,1.985 pfet_01v8_hvt
M$2 7 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=137500000000P
+ AD=140000000000P PS=1275000U PD=1280000U
* device instance $3 r0 *1 1.325,1.985 pfet_01v8_hvt
M$3 8 5 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=165000000000P PS=1280000U PD=1330000U
* device instance $4 r0 *1 1.805,1.985 pfet_01v8_hvt
M$4 12 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=172500000000P PS=1330000U PD=1345000U
* device instance $5 r0 *1 2.3,1.985 pfet_01v8_hvt
M$5 9 6 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=172500000000P
+ AD=260000000000P PS=1345000U PD=2520000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 14 2 10 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=89375000000P
+ PS=1820000U PD=925000U
* device instance $7 r0 *1 0.895,0.56 nfet_01v8
M$7 13 3 14 11 nfet_01v8 L=150000U W=650000U AS=89375000000P AD=91000000000P
+ PS=925000U PD=930000U
* device instance $8 r0 *1 1.325,0.56 nfet_01v8
M$8 9 5 13 11 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=115375000000P
+ PS=930000U PD=1005000U
* device instance $9 r0 *1 1.83,0.56 nfet_01v8
M$9 10 4 9 11 nfet_01v8 L=150000U W=650000U AS=115375000000P AD=112125000000P
+ PS=1005000U PD=995000U
* device instance $10 r0 *1 2.325,0.56 nfet_01v8
M$10 9 6 10 11 nfet_01v8 L=150000U W=650000U AS=112125000000P AD=169000000000P
+ PS=995000U PD=1820000U
.ENDS sky130_fd_sc_hd__a311oi_1

* cell sky130_fd_sc_hd__a2bb2oi_4
* pin VGND
* pin B2
* pin B1
* pin Y
* pin A1_N
* pin A2_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a2bb2oi_4 1 2 4 6 7 8 11 12 13
* net 1 VGND
* net 2 B2
* net 4 B1
* net 6 Y
* net 7 A1_N
* net 8 A2_N
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 6.03,1.985 pfet_01v8_hvt
M$1 11 7 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 7.71,1.985 pfet_01v8_hvt
M$5 3 8 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=685000000000P PS=5080000U PD=6370000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 11 4 9 12 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $12 r0 *1 1.73,1.985 pfet_01v8_hvt
M$12 9 2 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $17 r0 *1 3.83,1.985 pfet_01v8_hvt
M$17 6 3 9 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 0.47,0.56 nfet_01v8
M$21 5 4 1 13 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $24 r0 *1 1.73,0.56 nfet_01v8
M$24 6 2 5 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $29 r0 *1 3.83,0.56 nfet_01v8
M$29 6 3 1 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=520000000000P
+ PS=3680000U PD=4200000U
* device instance $33 r0 *1 6.03,0.56 nfet_01v8
M$33 3 7 1 13 nfet_01v8 L=150000U W=2600000U AS=520000000000P AD=351000000000P
+ PS=4200000U PD=3680000U
* device instance $37 r0 *1 7.71,0.56 nfet_01v8
M$37 3 8 1 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__a2bb2oi_4

* cell sky130_fd_sc_hd__nor3b_4
* pin VGND
* pin A
* pin B
* pin Y
* pin C_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor3b_4 1 2 3 4 5 7 10 11
* net 1 VGND
* net 2 A
* net 3 B
* net 4 Y
* net 5 C_N
* net 7 VPWR
* net 10 VPB
* device instance $1 r0 *1 3.11,1.985 pfet_01v8_hvt
M$1 8 3 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 4.79,1.985 pfet_01v8_hvt
M$5 4 6 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $9 r0 *1 0.49,1.985 pfet_01v8_hvt
M$9 7 5 6 10 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=135000000000P PS=2560000U PD=1270000U
* device instance $10 r0 *1 0.91,1.985 pfet_01v8_hvt
M$10 8 2 7 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $14 r0 *1 0.49,0.56 nfet_01v8
M$14 1 5 6 11 nfet_01v8 L=150000U W=650000U AS=182000000000P AD=87750000000P
+ PS=1860000U PD=920000U
* device instance $15 r0 *1 0.91,0.56 nfet_01v8
M$15 4 2 1 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=520000000000P
+ PS=3680000U PD=4200000U
* device instance $19 r0 *1 3.11,0.56 nfet_01v8
M$19 4 3 1 11 nfet_01v8 L=150000U W=2600000U AS=520000000000P AD=351000000000P
+ PS=4200000U PD=3680000U
* device instance $23 r0 *1 4.79,0.56 nfet_01v8
M$23 4 6 1 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nor3b_4

* cell sky130_fd_sc_hd__o22ai_2
* pin VGND
* pin B1
* pin Y
* pin B2
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o22ai_2 1 3 4 5 6 7 9 11 12
* net 1 VGND
* net 3 B1
* net 4 Y
* net 5 B2
* net 6 A2
* net 7 A1
* net 9 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.73,1.985 pfet_01v8_hvt
M$1 4 6 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 3.57,1.985 pfet_01v8_hvt
M$3 9 7 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $5 r0 *1 0.49,1.985 pfet_01v8_hvt
M$5 9 3 8 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $7 r0 *1 1.33,1.985 pfet_01v8_hvt
M$7 4 5 8 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $9 r0 *1 0.49,0.56 nfet_01v8
M$9 4 3 2 12 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $11 r0 *1 1.33,0.56 nfet_01v8
M$11 4 5 2 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=357500000000P
+ PS=1840000U PD=2400000U
* device instance $13 r0 *1 2.73,0.56 nfet_01v8
M$13 1 6 2 12 nfet_01v8 L=150000U W=1300000U AS=357500000000P AD=175500000000P
+ PS=2400000U PD=1840000U
* device instance $15 r0 *1 3.57,0.56 nfet_01v8
M$15 1 7 2 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__o22ai_2

* cell sky130_fd_sc_hd__o311a_4
* pin VGND
* pin X
* pin C1
* pin B1
* pin A3
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311a_4 1 3 6 7 8 9 10 11 14 15
* net 1 VGND
* net 3 X
* net 6 C1
* net 7 B1
* net 8 A3
* net 9 A2
* net 10 A1
* net 11 VPWR
* net 14 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 3 2 11 14 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=710000000000P PS=6330000U PD=5420000U
* device instance $5 r0 *1 2.49,1.985 pfet_01v8_hvt
M$5 2 6 11 14 pfet_01v8_hvt L=150000U W=2000000U AS=440000000000P
+ AD=270000000000P PS=2880000U PD=2540000U
* device instance $7 r0 *1 3.33,1.985 pfet_01v8_hvt
M$7 2 7 11 14 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $9 r0 *1 4.71,1.985 pfet_01v8_hvt
M$9 2 8 12 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $11 r0 *1 6.07,1.985 pfet_01v8_hvt
M$11 12 9 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $13 r0 *1 6.91,1.985 pfet_01v8_hvt
M$13 11 10 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $15 r0 *1 4.88,0.56 nfet_01v8
M$15 1 8 5 15 nfet_01v8 L=150000U W=1300000U AS=370500000000P AD=289250000000P
+ PS=3090000U PD=2190000U
* device instance $17 r0 *1 6.07,0.56 nfet_01v8
M$17 1 9 5 15 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $19 r0 *1 6.91,0.56 nfet_01v8
M$19 1 10 5 15 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $21 r0 *1 0.47,0.56 nfet_01v8
M$21 3 2 1 15 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
* device instance $25 r0 *1 2.67,0.56 nfet_01v8
M$25 2 6 4 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $27 r0 *1 3.51,0.56 nfet_01v8
M$27 5 7 4 15 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__o311a_4

* cell sky130_fd_sc_hd__or4b_1
* pin VGND
* pin D_N
* pin X
* pin C
* pin A
* pin VPWR
* pin VPB
* pin B
* pin 
.SUBCKT sky130_fd_sc_hd__or4b_1 1 2 5 6 7 8 9 10 14
* net 1 VGND
* net 2 D_N
* net 5 X
* net 6 C
* net 7 A
* net 8 VPWR
* net 9 VPB
* net 10 B
* device instance $1 r0 *1 1.41,1.695 pfet_01v8_hvt
M$1 11 3 4 9 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=68250000000P
+ PS=1360000U PD=745000U
* device instance $2 r0 *1 1.885,1.695 pfet_01v8_hvt
M$2 13 6 11 9 pfet_01v8_hvt L=150000U W=420000U AS=68250000000P AD=45150000000P
+ PS=745000U PD=635000U
* device instance $3 r0 *1 2.25,1.695 pfet_01v8_hvt
M$3 12 10 13 9 pfet_01v8_hvt L=150000U W=420000U AS=45150000000P
+ AD=64050000000P PS=635000U PD=725000U
* device instance $4 r0 *1 2.705,1.695 pfet_01v8_hvt
M$4 8 7 12 9 pfet_01v8_hvt L=150000U W=420000U AS=64050000000P AD=148250000000P
+ PS=725000U PD=1340000U
* device instance $5 r0 *1 3.195,1.985 pfet_01v8_hvt
M$5 5 4 8 9 pfet_01v8_hvt L=150000U W=1000000U AS=148250000000P
+ AD=275000000000P PS=1340000U PD=2550000U
* device instance $6 r0 *1 0.47,1.695 pfet_01v8_hvt
M$6 3 2 8 9 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $7 r0 *1 1.41,0.475 nfet_01v8
M$7 4 3 1 14 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=64050000000P
+ PS=1360000U PD=725000U
* device instance $8 r0 *1 1.865,0.475 nfet_01v8
M$8 1 6 4 14 nfet_01v8 L=150000U W=420000U AS=64050000000P AD=56700000000P
+ PS=725000U PD=690000U
* device instance $9 r0 *1 2.285,0.475 nfet_01v8
M$9 4 10 1 14 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $10 r0 *1 2.705,0.475 nfet_01v8
M$10 4 7 1 14 nfet_01v8 L=150000U W=420000U AS=101875000000P AD=56700000000P
+ PS=990000U PD=690000U
* device instance $11 r0 *1 3.195,0.56 nfet_01v8
M$11 5 4 1 14 nfet_01v8 L=150000U W=650000U AS=101875000000P AD=178750000000P
+ PS=990000U PD=1850000U
* device instance $12 r0 *1 0.47,0.475 nfet_01v8
M$12 3 2 1 14 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__or4b_1

* cell sky130_fd_sc_hd__or4_2
* pin VPB
* pin D
* pin C
* pin B
* pin A
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__or4_2 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 D
* net 3 C
* net 4 B
* net 5 A
* net 7 VGND
* net 8 VPWR
* net 9 X
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 13 2 6 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=69300000000P
+ PS=1360000U PD=750000U
* device instance $2 r0 *1 0.95,1.695 pfet_01v8_hvt
M$2 12 3 13 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=44100000000P
+ PS=750000U PD=630000U
* device instance $3 r0 *1 1.31,1.695 pfet_01v8_hvt
M$3 11 4 12 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $4 r0 *1 1.79,1.695 pfet_01v8_hvt
M$4 8 5 11 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=148250000000P
+ PS=750000U PD=1340000U
* device instance $5 r0 *1 2.28,1.985 pfet_01v8_hvt
M$5 9 6 8 1 pfet_01v8_hvt L=150000U W=2000000U AS=283250000000P
+ AD=440000000000P PS=2610000U PD=3880000U
* device instance $7 r0 *1 0.47,0.475 nfet_01v8
M$7 6 2 7 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=69300000000P
+ PS=1360000U PD=750000U
* device instance $8 r0 *1 0.95,0.475 nfet_01v8
M$8 7 3 6 10 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=56700000000P
+ PS=750000U PD=690000U
* device instance $9 r0 *1 1.37,0.475 nfet_01v8
M$9 6 4 7 10 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $10 r0 *1 1.79,0.475 nfet_01v8
M$10 6 5 7 10 nfet_01v8 L=150000U W=420000U AS=101875000000P AD=56700000000P
+ PS=990000U PD=690000U
* device instance $11 r0 *1 2.28,0.56 nfet_01v8
M$11 9 6 7 10 nfet_01v8 L=150000U W=1300000U AS=189625000000P AD=286000000000P
+ PS=1910000U PD=2830000U
.ENDS sky130_fd_sc_hd__or4_2

* cell sky130_fd_sc_hd__nand4b_1
* pin VPB
* pin A_N
* pin B
* pin C
* pin D
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__nand4b_1 1 2 3 4 6 7 8 9 10
* net 1 VPB
* net 2 A_N
* net 3 B
* net 4 C
* net 6 D
* net 7 VPWR
* net 8 Y
* net 9 VGND
* device instance $1 r0 *1 0.6,1.695 pfet_01v8_hvt
M$1 7 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=145750000000P
+ PS=1360000U PD=1335000U
* device instance $2 r0 *1 1.085,1.985 pfet_01v8_hvt
M$2 8 6 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=145750000000P
+ AD=135000000000P PS=1335000U PD=1270000U
* device instance $3 r0 *1 1.505,1.985 pfet_01v8_hvt
M$3 7 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=192500000000P PS=1270000U PD=1385000U
* device instance $4 r0 *1 2.04,1.985 pfet_01v8_hvt
M$4 8 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=192500000000P
+ AD=195000000000P PS=1385000U PD=1390000U
* device instance $5 r0 *1 2.58,1.985 pfet_01v8_hvt
M$5 7 5 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=280000000000P PS=1390000U PD=2560000U
* device instance $6 r0 *1 0.545,0.675 nfet_01v8
M$6 5 2 9 10 nfet_01v8 L=150000U W=420000U AS=118125000000P AD=111300000000P
+ PS=1040000U PD=1370000U
* device instance $7 r0 *1 1.085,0.56 nfet_01v8
M$7 11 6 9 10 nfet_01v8 L=150000U W=650000U AS=118125000000P AD=87750000000P
+ PS=1040000U PD=920000U
* device instance $8 r0 *1 1.505,0.56 nfet_01v8
M$8 13 4 11 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=125125000000P
+ PS=920000U PD=1035000U
* device instance $9 r0 *1 2.04,0.56 nfet_01v8
M$9 12 3 13 10 nfet_01v8 L=150000U W=650000U AS=125125000000P AD=126750000000P
+ PS=1035000U PD=1040000U
* device instance $10 r0 *1 2.58,0.56 nfet_01v8
M$10 8 5 12 10 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=227500000000P
+ PS=1040000U PD=2000000U
.ENDS sky130_fd_sc_hd__nand4b_1

* cell sky130_fd_sc_hd__nand3b_1
* pin VPB
* pin A_N
* pin C
* pin B
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nand3b_1 1 2 3 4 5 7 8 9
* net 1 VPB
* net 2 A_N
* net 3 C
* net 4 B
* net 5 Y
* net 7 VGND
* net 8 VPWR
* device instance $1 r0 *1 0.6,1.695 pfet_01v8_hvt
M$1 8 2 6 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=145750000000P
+ PS=1360000U PD=1335000U
* device instance $2 r0 *1 1.085,1.985 pfet_01v8_hvt
M$2 5 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=145750000000P
+ AD=135000000000P PS=1335000U PD=1270000U
* device instance $3 r0 *1 1.505,1.985 pfet_01v8_hvt
M$3 8 4 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=192500000000P PS=1270000U PD=1385000U
* device instance $4 r0 *1 2.04,1.985 pfet_01v8_hvt
M$4 5 6 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=192500000000P
+ AD=280000000000P PS=1385000U PD=2560000U
* device instance $5 r0 *1 0.6,0.675 nfet_01v8
M$5 6 2 7 9 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
* device instance $6 r0 *1 1.085,0.56 nfet_01v8
M$6 11 3 7 9 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=87750000000P
+ PS=985000U PD=920000U
* device instance $7 r0 *1 1.505,0.56 nfet_01v8
M$7 10 4 11 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=125125000000P
+ PS=920000U PD=1035000U
* device instance $8 r0 *1 2.04,0.56 nfet_01v8
M$8 5 6 10 9 nfet_01v8 L=150000U W=650000U AS=125125000000P AD=182000000000P
+ PS=1035000U PD=1860000U
.ENDS sky130_fd_sc_hd__nand3b_1

* cell sky130_fd_sc_hd__a2111o_1
* pin VGND
* pin X
* pin A1
* pin D1
* pin C1
* pin B1
* pin A2
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a2111o_1 1 2 4 5 6 7 8 11 12 15
* net 1 VGND
* net 2 X
* net 4 A1
* net 5 D1
* net 6 C1
* net 7 B1
* net 8 A2
* net 11 VPB
* net 12 VPWR
* device instance $1 r0 *1 1.595,1.985 pfet_01v8_hvt
M$1 13 5 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=385000000000P
+ AD=125000000000P PS=2770000U PD=1250000U
* device instance $2 r0 *1 1.995,1.985 pfet_01v8_hvt
M$2 14 6 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=125000000000P
+ AD=180000000000P PS=1250000U PD=1360000U
* device instance $3 r0 *1 2.505,1.985 pfet_01v8_hvt
M$3 10 7 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=180000000000P
+ AD=280000000000P PS=1360000U PD=1560000U
* device instance $4 r0 *1 3.215,1.985 pfet_01v8_hvt
M$4 12 4 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=135000000000P PS=1560000U PD=1270000U
* device instance $5 r0 *1 3.635,1.985 pfet_01v8_hvt
M$5 10 8 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=290000000000P PS=1270000U PD=2580000U
* device instance $6 r0 *1 0.5,1.985 pfet_01v8_hvt
M$6 12 3 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=290000000000P
+ AD=265000000000P PS=2580000U PD=2530000U
* device instance $7 r0 *1 0.54,0.56 nfet_01v8
M$7 1 3 2 15 nfet_01v8 L=150000U W=650000U AS=214500000000P AD=274625000000P
+ PS=1960000U PD=1495000U
* device instance $8 r0 *1 1.535,0.56 nfet_01v8
M$8 3 5 1 15 nfet_01v8 L=150000U W=650000U AS=274625000000P AD=100750000000P
+ PS=1495000U PD=960000U
* device instance $9 r0 *1 1.995,0.56 nfet_01v8
M$9 1 6 3 15 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=117000000000P
+ PS=960000U PD=1010000U
* device instance $10 r0 *1 2.505,0.56 nfet_01v8
M$10 3 7 1 15 nfet_01v8 L=150000U W=650000U AS=117000000000P AD=185250000000P
+ PS=1010000U PD=1220000U
* device instance $11 r0 *1 3.225,0.56 nfet_01v8
M$11 9 4 3 15 nfet_01v8 L=150000U W=650000U AS=185250000000P AD=82875000000P
+ PS=1220000U PD=905000U
* device instance $12 r0 *1 3.63,0.56 nfet_01v8
M$12 1 8 9 15 nfet_01v8 L=150000U W=650000U AS=82875000000P AD=188500000000P
+ PS=905000U PD=1880000U
.ENDS sky130_fd_sc_hd__a2111o_1

* cell sky130_fd_sc_hd__or4b_2
* pin VPB
* pin A
* pin C
* pin B
* pin D_N
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__or4b_2 1 2 3 4 5 7 8 9 11
* net 1 VPB
* net 2 A
* net 3 C
* net 4 B
* net 5 D_N
* net 7 VGND
* net 8 VPWR
* net 9 X
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 8 5 10 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=169300000000P PS=1360000U PD=1500000U
* device instance $2 r0 *1 1.86,1.695 pfet_01v8_hvt
M$2 14 2 8 1 pfet_01v8_hvt L=150000U W=420000U AS=168350000000P AD=69300000000P
+ PS=1495000U PD=750000U
* device instance $3 r0 *1 2.34,1.695 pfet_01v8_hvt
M$3 13 4 14 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=44100000000P
+ PS=750000U PD=630000U
* device instance $4 r0 *1 2.7,1.695 pfet_01v8_hvt
M$4 12 3 13 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $5 r0 *1 3.18,1.695 pfet_01v8_hvt
M$5 6 10 12 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P
+ AD=109200000000P PS=750000U PD=1360000U
* device instance $6 r0 *1 0.955,1.985 pfet_01v8_hvt
M$6 9 6 8 1 pfet_01v8_hvt L=150000U W=2000000U AS=304300000000P
+ AD=303350000000P PS=2770000U PD=2765000U
* device instance $8 r0 *1 0.47,0.475 nfet_01v8
M$8 10 5 7 11 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
* device instance $9 r0 *1 1.86,0.475 nfet_01v8
M$9 6 2 7 11 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=69300000000P
+ PS=985000U PD=750000U
* device instance $10 r0 *1 2.34,0.475 nfet_01v8
M$10 7 4 6 11 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=56700000000P
+ PS=750000U PD=690000U
* device instance $11 r0 *1 2.76,0.475 nfet_01v8
M$11 6 3 7 11 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $12 r0 *1 3.18,0.475 nfet_01v8
M$12 7 10 6 11 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $13 r0 *1 0.955,0.56 nfet_01v8
M$13 9 6 7 11 nfet_01v8 L=150000U W=1300000U AS=188000000000P AD=188000000000P
+ PS=1905000U PD=1905000U
.ENDS sky130_fd_sc_hd__or4b_2

* cell sky130_fd_sc_hd__a311o_2
* pin VGND
* pin X
* pin A3
* pin A2
* pin A1
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a311o_2 1 2 6 7 8 9 10 11 13 15
* net 1 VGND
* net 2 X
* net 6 A3
* net 7 A2
* net 8 A1
* net 9 B1
* net 10 C1
* net 11 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 2 3 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=375000000000P PS=3790000U PD=2750000U
* device instance $3 r0 *1 1.52,1.985 pfet_01v8_hvt
M$3 12 6 11 13 pfet_01v8_hvt L=150000U W=1000000U AS=240000000000P
+ AD=170000000000P PS=1480000U PD=1340000U
* device instance $4 r0 *1 2.01,1.985 pfet_01v8_hvt
M$4 11 7 12 13 pfet_01v8_hvt L=150000U W=1000000U AS=170000000000P
+ AD=185000000000P PS=1340000U PD=1370000U
* device instance $5 r0 *1 2.53,1.985 pfet_01v8_hvt
M$5 12 8 11 13 pfet_01v8_hvt L=150000U W=1000000U AS=185000000000P
+ AD=210000000000P PS=1370000U PD=1420000U
* device instance $6 r0 *1 3.1,1.985 pfet_01v8_hvt
M$6 14 9 12 13 pfet_01v8_hvt L=150000U W=1000000U AS=210000000000P
+ AD=210000000000P PS=1420000U PD=1420000U
* device instance $7 r0 *1 3.67,1.985 pfet_01v8_hvt
M$7 3 10 14 13 pfet_01v8_hvt L=150000U W=1000000U AS=210000000000P
+ AD=260000000000P PS=1420000U PD=2520000U
* device instance $8 r0 *1 0.47,0.56 nfet_01v8
M$8 2 3 1 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=243750000000P
+ PS=2740000U PD=2050000U
* device instance $10 r0 *1 1.52,0.56 nfet_01v8
M$10 5 6 1 15 nfet_01v8 L=150000U W=650000U AS=156000000000P AD=110500000000P
+ PS=1130000U PD=990000U
* device instance $11 r0 *1 2.01,0.56 nfet_01v8
M$11 4 7 5 15 nfet_01v8 L=150000U W=650000U AS=110500000000P AD=120250000000P
+ PS=990000U PD=1020000U
* device instance $12 r0 *1 2.53,0.56 nfet_01v8
M$12 3 8 4 15 nfet_01v8 L=150000U W=650000U AS=120250000000P AD=133250000000P
+ PS=1020000U PD=1060000U
* device instance $13 r0 *1 3.09,0.56 nfet_01v8
M$13 1 9 3 15 nfet_01v8 L=150000U W=650000U AS=133250000000P AD=139750000000P
+ PS=1060000U PD=1080000U
* device instance $14 r0 *1 3.67,0.56 nfet_01v8
M$14 3 10 1 15 nfet_01v8 L=150000U W=650000U AS=139750000000P AD=169000000000P
+ PS=1080000U PD=1820000U
.ENDS sky130_fd_sc_hd__a311o_2

* cell sky130_fd_sc_hd__inv_4
* pin VPB
* pin A
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__inv_4 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 VGND
* net 4 VPWR
* net 5 Y
* device instance $1 r0 *1 0.52,1.985 pfet_01v8_hvt
M$1 5 2 4 1 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=665000000000P PS=6330000U PD=6330000U
* device instance $5 r0 *1 0.52,0.56 nfet_01v8
M$5 5 2 3 6 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
.ENDS sky130_fd_sc_hd__inv_4

* cell sky130_fd_sc_hd__a22o_2
* pin VGND
* pin B1
* pin A1
* pin X
* pin B2
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a22o_2 1 3 4 5 8 9 11 12 13
* net 1 VGND
* net 3 B1
* net 4 A1
* net 5 X
* net 8 B2
* net 9 A2
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 1.83,1.985 pfet_01v8_hvt
M$1 10 4 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=165000000000P PS=2520000U PD=1330000U
* device instance $2 r0 *1 2.31,1.985 pfet_01v8_hvt
M$2 11 9 10 12 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=157500000000P PS=1330000U PD=1315000U
* device instance $3 r0 *1 2.775,1.985 pfet_01v8_hvt
M$3 5 2 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=292500000000P
+ AD=405000000000P PS=2585000U PD=3810000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 10 8 2 12 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $6 r0 *1 0.89,1.985 pfet_01v8_hvt
M$6 2 3 10 12 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $7 r0 *1 1.83,0.56 nfet_01v8
M$7 7 4 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $8 r0 *1 2.31,0.56 nfet_01v8
M$8 1 9 7 13 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=102375000000P
+ PS=980000U PD=965000U
* device instance $9 r0 *1 2.775,0.56 nfet_01v8
M$9 5 2 1 13 nfet_01v8 L=150000U W=1300000U AS=190125000000P AD=263250000000P
+ PS=1885000U PD=2760000U
* device instance $11 r0 *1 0.47,0.56 nfet_01v8
M$11 6 8 1 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=74750000000P
+ PS=1820000U PD=880000U
* device instance $12 r0 *1 0.85,0.56 nfet_01v8
M$12 2 3 6 13 nfet_01v8 L=150000U W=650000U AS=74750000000P AD=169000000000P
+ PS=880000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22o_2

* cell sky130_fd_sc_hd__o21ba_1
* pin VPB
* pin B1_N
* pin A2
* pin A1
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o21ba_1 1 2 3 4 8 9 10 11
* net 1 VPB
* net 2 B1_N
* net 3 A2
* net 4 A1
* net 8 X
* net 9 VPWR
* net 10 VGND
* device instance $1 r0 *1 2.165,1.985 pfet_01v8_hvt
M$1 6 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=300000000000P
+ AD=165000000000P PS=2600000U PD=1330000U
* device instance $2 r0 *1 2.645,1.985 pfet_01v8_hvt
M$2 12 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=105000000000P PS=1330000U PD=1210000U
* device instance $3 r0 *1 3.005,1.985 pfet_01v8_hvt
M$3 9 4 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=280000000000P PS=1210000U PD=2560000U
* device instance $4 r0 *1 1.035,1.695 pfet_01v8_hvt
M$4 5 2 9 1 pfet_01v8_hvt L=150000U W=420000U AS=185750000000P AD=117600000000P
+ PS=1415000U PD=1400000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 9 6 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=185750000000P PS=2520000U PD=1415000U
* device instance $6 r0 *1 2.165,0.56 nfet_01v8
M$6 7 5 6 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $7 r0 *1 2.645,0.56 nfet_01v8
M$7 10 3 7 11 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=87750000000P
+ PS=980000U PD=920000U
* device instance $8 r0 *1 3.065,0.56 nfet_01v8
M$8 7 4 10 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=172250000000P
+ PS=920000U PD=1830000U
* device instance $9 r0 *1 0.55,0.56 nfet_01v8
M$9 10 6 8 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=100250000000P
+ PS=1820000U PD=985000U
* device instance $10 r0 *1 1.035,0.675 nfet_01v8
M$10 5 2 10 11 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
.ENDS sky130_fd_sc_hd__o21ba_1

* cell sky130_fd_sc_hd__a221oi_4
* pin VGND
* pin B1
* pin C1
* pin Y
* pin B2
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a221oi_4 1 2 3 4 6 7 9 11 12 14
* net 1 VGND
* net 2 B1
* net 3 C1
* net 4 Y
* net 6 B2
* net 7 A2
* net 9 A1
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 2.69,1.985 pfet_01v8_hvt
M$1 10 6 13 12 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=580000000000P PS=6330000U PD=5160000U
* device instance $4 r0 *1 3.95,1.985 pfet_01v8_hvt
M$4 13 2 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $9 r0 *1 6.13,1.985 pfet_01v8_hvt
M$9 11 7 13 12 pfet_01v8_hvt L=150000U W=4000000U AS=580000000000P
+ AD=700000000000P PS=5160000U PD=6400000U
* device instance $10 r0 *1 6.55,1.985 pfet_01v8_hvt
M$10 13 9 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $17 r0 *1 0.49,1.985 pfet_01v8_hvt
M$17 4 3 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=665000000000P PS=6370000U PD=6330000U
* device instance $21 r0 *1 0.49,0.56 nfet_01v8
M$21 4 3 1 14 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=357500000000P
+ PS=4620000U PD=3700000U
* device instance $25 r0 *1 2.19,0.56 nfet_01v8
M$25 5 6 1 14 nfet_01v8 L=150000U W=2600000U AS=357500000000P AD=539500000000P
+ PS=3700000U PD=4260000U
* device instance $28 r0 *1 3.95,0.56 nfet_01v8
M$28 4 2 5 14 nfet_01v8 L=150000U W=2600000U AS=513500000000P AD=351000000000P
+ PS=4180000U PD=3680000U
* device instance $33 r0 *1 6.13,0.56 nfet_01v8
M$33 8 7 1 14 nfet_01v8 L=150000U W=2600000U AS=377000000000P AD=432250000000P
+ PS=3760000U PD=4580000U
* device instance $34 r0 *1 6.55,0.56 nfet_01v8
M$34 4 9 8 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
.ENDS sky130_fd_sc_hd__a221oi_4

* cell sky130_fd_sc_hd__a31o_4
* pin VGND
* pin A3
* pin A2
* pin A1
* pin B1
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a31o_4 1 2 3 4 5 7 13 14 15
* net 1 VGND
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 B1
* net 7 X
* net 13 VPWR
* net 14 VPB
* device instance $1 r0 *1 4.47,1.985 pfet_01v8_hvt
M$1 7 6 13 14 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=905000000000P PS=6330000U PD=6810000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 13 2 12 14 pfet_01v8_hvt L=150000U W=2000000U AS=425000000000P
+ AD=300000000000P PS=3850000U PD=2600000U
* device instance $6 r0 *1 0.89,1.985 pfet_01v8_hvt
M$6 12 3 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=300000000000P PS=2540000U PD=2600000U
* device instance $7 r0 *1 1.31,1.985 pfet_01v8_hvt
M$7 13 4 12 14 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $11 r0 *1 3.11,1.985 pfet_01v8_hvt
M$11 6 5 12 14 pfet_01v8_hvt L=150000U W=2000000U AS=300000000000P
+ AD=395000000000P PS=2600000U PD=3790000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 8 2 1 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $14 r0 *1 0.89,0.56 nfet_01v8
M$14 9 3 8 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $15 r0 *1 1.31,0.56 nfet_01v8
M$15 6 4 9 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $16 r0 *1 1.73,0.56 nfet_01v8
M$16 11 4 6 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $17 r0 *1 2.15,0.56 nfet_01v8
M$17 10 3 11 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $18 r0 *1 2.63,0.56 nfet_01v8
M$18 1 2 10 15 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=107250000000P
+ PS=980000U PD=980000U
* device instance $19 r0 *1 3.11,0.56 nfet_01v8
M$19 6 5 1 15 nfet_01v8 L=150000U W=1300000U AS=195000000000P AD=344500000000P
+ PS=1900000U PD=2360000U
* device instance $21 r0 *1 4.47,0.56 nfet_01v8
M$21 7 6 1 15 nfet_01v8 L=150000U W=2600000U AS=520000000000P AD=432250000000P
+ PS=4200000U PD=4580000U
.ENDS sky130_fd_sc_hd__a31o_4

* cell sky130_fd_sc_hd__a211o_4
* pin VGND
* pin X
* pin B1
* pin C1
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a211o_4 1 2 4 5 6 7 10 11 15
* net 1 VGND
* net 2 X
* net 4 B1
* net 5 C1
* net 6 A2
* net 7 A1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.7,1.985 pfet_01v8_hvt
M$1 13 4 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=140000000000P PS=2520000U PD=1280000U
* device instance $2 r0 *1 3.13,1.985 pfet_01v8_hvt
M$2 3 5 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $3 r0 *1 3.56,1.985 pfet_01v8_hvt
M$3 14 5 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=160000000000P PS=1280000U PD=1320000U
* device instance $4 r0 *1 4.03,1.985 pfet_01v8_hvt
M$4 12 4 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=160000000000P
+ AD=195000000000P PS=1320000U PD=1390000U
* device instance $5 r0 *1 4.57,1.985 pfet_01v8_hvt
M$5 10 6 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=335000000000P
+ AD=455000000000P PS=2670000U PD=3910000U
* device instance $6 r0 *1 5.11,1.985 pfet_01v8_hvt
M$6 12 7 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=335000000000P
+ AD=280000000000P PS=2670000U PD=2560000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 2 3 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=680000000000P
+ AD=680000000000P PS=6360000U PD=6360000U
* device instance $13 r0 *1 0.865,0.56 nfet_01v8
M$13 2 3 1 15 nfet_01v8 L=150000U W=2600000U AS=450125000000P AD=370500000000P
+ PS=4635000U PD=3740000U
* device instance $17 r0 *1 2.605,0.56 nfet_01v8
M$17 3 4 1 15 nfet_01v8 L=150000U W=1300000U AS=219375000000P AD=243750000000P
+ PS=1975000U PD=2050000U
* device instance $18 r0 *1 3.075,0.56 nfet_01v8
M$18 1 5 3 15 nfet_01v8 L=150000U W=1300000U AS=212875000000P AD=235625000000P
+ PS=1955000U PD=2025000U
* device instance $21 r0 *1 4.68,0.56 nfet_01v8
M$21 8 6 1 15 nfet_01v8 L=150000U W=650000U AS=139750000000P AD=91000000000P
+ PS=1080000U PD=930000U
* device instance $22 r0 *1 5.11,0.56 nfet_01v8
M$22 3 7 8 15 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=91000000000P
+ PS=930000U PD=930000U
* device instance $23 r0 *1 5.54,0.56 nfet_01v8
M$23 9 7 3 15 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=91000000000P
+ PS=930000U PD=930000U
* device instance $24 r0 *1 5.97,0.56 nfet_01v8
M$24 1 6 9 15 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=169000000000P
+ PS=930000U PD=1820000U
.ENDS sky130_fd_sc_hd__a211o_4

* cell sky130_fd_sc_hd__a2111oi_2
* pin VGND
* pin Y
* pin C1
* pin D1
* pin B1
* pin A1
* pin A2
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a2111oi_2 1 2 3 4 5 6 7 10 11 16
* net 1 VGND
* net 2 Y
* net 3 C1
* net 4 D1
* net 5 B1
* net 6 A1
* net 7 A2
* net 10 VPB
* net 11 VPWR
* device instance $1 r0 *1 3.64,1.985 pfet_01v8_hvt
M$1 11 6 13 10 pfet_01v8_hvt L=150000U W=2000000U AS=420000000000P
+ AD=475000000000P PS=3840000U PD=3950000U
* device instance $2 r0 *1 4.07,1.985 pfet_01v8_hvt
M$2 13 7 11 10 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=300000000000P PS=2560000U PD=2600000U
* device instance $5 r0 *1 0.5,1.985 pfet_01v8_hvt
M$5 14 3 12 10 pfet_01v8_hvt L=150000U W=1000000U AS=285000000000P
+ AD=140000000000P PS=2570000U PD=1280000U
* device instance $6 r0 *1 0.93,1.985 pfet_01v8_hvt
M$6 2 4 14 10 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $7 r0 *1 1.36,1.985 pfet_01v8_hvt
M$7 15 4 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $8 r0 *1 1.79,1.985 pfet_01v8_hvt
M$8 12 3 15 10 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=160000000000P PS=1280000U PD=1320000U
* device instance $9 r0 *1 2.26,1.985 pfet_01v8_hvt
M$9 13 5 12 10 pfet_01v8_hvt L=150000U W=2000000U AS=300000000000P
+ AD=400000000000P PS=2600000U PD=3800000U
* device instance $11 r0 *1 0.5,0.56 nfet_01v8
M$11 1 3 2 16 nfet_01v8 L=150000U W=1300000U AS=312000000000P AD=196625000000P
+ PS=2910000U PD=1905000U
* device instance $12 r0 *1 0.93,0.56 nfet_01v8
M$12 2 4 1 16 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=217750000000P
+ PS=1860000U PD=1970000U
* device instance $15 r0 *1 2.375,0.56 nfet_01v8
M$15 1 5 2 16 nfet_01v8 L=150000U W=1300000U AS=232375000000P AD=217750000000P
+ PS=2015000U PD=1970000U
* device instance $17 r0 *1 3.345,0.56 nfet_01v8
M$17 9 6 2 16 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=178750000000P
+ PS=930000U PD=1200000U
* device instance $18 r0 *1 4.045,0.56 nfet_01v8
M$18 1 7 9 16 nfet_01v8 L=150000U W=650000U AS=178750000000P AD=112125000000P
+ PS=1200000U PD=995000U
* device instance $19 r0 *1 4.54,0.56 nfet_01v8
M$19 8 7 1 16 nfet_01v8 L=150000U W=650000U AS=112125000000P AD=91000000000P
+ PS=995000U PD=930000U
* device instance $20 r0 *1 4.97,0.56 nfet_01v8
M$20 2 6 8 16 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=172250000000P
+ PS=930000U PD=1830000U
.ENDS sky130_fd_sc_hd__a2111oi_2

* cell sky130_fd_sc_hd__o41ai_2
* pin VGND
* pin Y
* pin B1
* pin A4
* pin A3
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o41ai_2 1 3 4 5 6 7 8 9 13 14
* net 1 VGND
* net 3 Y
* net 4 B1
* net 5 A4
* net 6 A3
* net 7 A2
* net 8 A1
* net 9 VPWR
* net 13 VPB
* device instance $1 r0 *1 4.07,1.985 pfet_01v8_hvt
M$1 11 7 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 4.91,1.985 pfet_01v8_hvt
M$3 9 8 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $5 r0 *1 1.83,1.985 pfet_01v8_hvt
M$5 3 5 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $7 r0 *1 2.67,1.985 pfet_01v8_hvt
M$7 11 6 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 3 4 9 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $11 r0 *1 4.07,0.56 nfet_01v8
M$11 1 7 2 14 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $13 r0 *1 4.91,0.56 nfet_01v8
M$13 1 8 2 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
* device instance $15 r0 *1 1.83,0.56 nfet_01v8
M$15 2 5 1 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $17 r0 *1 2.67,0.56 nfet_01v8
M$17 2 6 1 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
* device instance $19 r0 *1 0.47,0.56 nfet_01v8
M$19 3 4 2 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
.ENDS sky130_fd_sc_hd__o41ai_2

* cell sky130_fd_sc_hd__nor4bb_1
* pin VPB
* pin C_N
* pin D_N
* pin B
* pin A
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor4bb_1 1 2 3 5 6 8 9 10 11
* net 1 VPB
* net 2 C_N
* net 3 D_N
* net 5 B
* net 6 A
* net 8 Y
* net 9 VGND
* net 10 VPWR
* device instance $1 r0 *1 1.89,1.985 pfet_01v8_hvt
M$1 14 7 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=255900000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.31,1.985 pfet_01v8_hvt
M$2 13 4 14 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $3 r0 *1 2.79,1.985 pfet_01v8_hvt
M$3 12 5 13 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=135000000000P PS=1330000U PD=1270000U
* device instance $4 r0 *1 3.21,1.985 pfet_01v8_hvt
M$4 10 6 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $5 r0 *1 0.955,1.695 pfet_01v8_hvt
M$5 7 3 10 1 pfet_01v8_hvt L=150000U W=420000U AS=122612500000P
+ AD=108500000000P PS=1320000U PD=1360000U
* device instance $6 r0 *1 0.47,2.26 pfet_01v8_hvt
M$6 4 2 10 1 pfet_01v8_hvt L=150000U W=420000U AS=122612500000P
+ AD=109200000000P PS=1320000U PD=1360000U
* device instance $7 r0 *1 1.89,0.56 nfet_01v8
M$7 8 7 9 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 2.31,0.56 nfet_01v8
M$8 9 4 8 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $9 r0 *1 2.79,0.56 nfet_01v8
M$9 8 5 9 11 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=87750000000P
+ PS=980000U PD=920000U
* device instance $10 r0 *1 3.21,0.56 nfet_01v8
M$10 9 6 8 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $11 r0 *1 0.51,0.675 nfet_01v8
M$11 9 2 4 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=60900000000P
+ PS=1360000U PD=710000U
* device instance $12 r0 *1 0.95,0.675 nfet_01v8
M$12 7 3 9 11 nfet_01v8 L=150000U W=420000U AS=60900000000P AD=109200000000P
+ PS=710000U PD=1360000U
.ENDS sky130_fd_sc_hd__nor4bb_1

* cell sky130_fd_sc_hd__a21boi_1
* pin VPB
* pin B1_N
* pin A1
* pin A2
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__a21boi_1 1 2 3 4 6 7 9 10
* net 1 VPB
* net 2 B1_N
* net 3 A1
* net 4 A2
* net 6 VPWR
* net 7 VGND
* net 9 Y
* device instance $1 r0 *1 1.425,1.985 pfet_01v8_hvt
M$1 8 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 1.855,1.985 pfet_01v8_hvt
M$2 6 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $3 r0 *1 2.285,1.985 pfet_01v8_hvt
M$3 8 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=265000000000P PS=1280000U PD=2530000U
* device instance $4 r0 *1 0.475,2.275 pfet_01v8_hvt
M$4 6 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=111300000000P AD=111300000000P
+ PS=1370000U PD=1370000U
* device instance $5 r0 *1 0.765,0.445 nfet_01v8
M$5 7 2 5 10 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=101875000000P
+ PS=1370000U PD=990000U
* device instance $6 r0 *1 1.255,0.56 nfet_01v8
M$6 9 5 7 10 nfet_01v8 L=150000U W=650000U AS=101875000000P AD=143000000000P
+ PS=990000U PD=1090000U
* device instance $7 r0 *1 1.845,0.56 nfet_01v8
M$7 11 3 9 10 nfet_01v8 L=150000U W=650000U AS=143000000000P AD=91000000000P
+ PS=1090000U PD=930000U
* device instance $8 r0 *1 2.275,0.56 nfet_01v8
M$8 7 4 11 10 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=172250000000P
+ PS=930000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21boi_1

* cell sky130_fd_sc_hd__o32ai_1
* pin VGND
* pin B1
* pin Y
* pin B2
* pin A3
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o32ai_1 1 2 4 5 6 7 8 9 10 12
* net 1 VGND
* net 2 B1
* net 4 Y
* net 5 B2
* net 6 A3
* net 7 A2
* net 8 A1
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 11 2 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=105000000000P PS=2520000U PD=1210000U
* device instance $2 r0 *1 0.83,1.985 pfet_01v8_hvt
M$2 4 5 11 10 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=305000000000P PS=1210000U PD=1610000U
* device instance $3 r0 *1 1.59,1.985 pfet_01v8_hvt
M$3 13 6 4 10 pfet_01v8_hvt L=150000U W=1000000U AS=305000000000P
+ AD=245000000000P PS=1610000U PD=1490000U
* device instance $4 r0 *1 2.23,1.985 pfet_01v8_hvt
M$4 14 7 13 10 pfet_01v8_hvt L=150000U W=1000000U AS=245000000000P
+ AD=135000000000P PS=1490000U PD=1270000U
* device instance $5 r0 *1 2.65,1.985 pfet_01v8_hvt
M$5 9 8 14 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=280000000000P PS=1270000U PD=2560000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 4 2 3 12 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=105625000000P
+ PS=1820000U PD=975000U
* device instance $7 r0 *1 0.945,0.56 nfet_01v8
M$7 3 5 4 12 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=100750000000P
+ PS=975000U PD=960000U
* device instance $8 r0 *1 1.405,0.56 nfet_01v8
M$8 1 6 3 12 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=219375000000P
+ PS=960000U PD=1325000U
* device instance $9 r0 *1 2.23,0.56 nfet_01v8
M$9 3 7 1 12 nfet_01v8 L=150000U W=650000U AS=219375000000P AD=87750000000P
+ PS=1325000U PD=920000U
* device instance $10 r0 *1 2.65,0.56 nfet_01v8
M$10 1 8 3 12 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=234000000000P
+ PS=920000U PD=2020000U
.ENDS sky130_fd_sc_hd__o32ai_1

* cell sky130_fd_sc_hd__a31o_2
* pin VPB
* pin B1
* pin A1
* pin A2
* pin A3
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a31o_2 1 2 3 4 5 6 7 8 11
* net 1 VPB
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 A3
* net 6 X
* net 7 VPWR
* net 8 VGND
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 6 10 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 9 5 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $4 r0 *1 1.73,1.985 pfet_01v8_hvt
M$4 7 4 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $5 r0 *1 2.21,1.985 pfet_01v8_hvt
M$5 9 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=165000000000P PS=1330000U PD=1330000U
* device instance $6 r0 *1 2.69,1.985 pfet_01v8_hvt
M$6 10 2 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=320000000000P PS=1330000U PD=2640000U
* device instance $7 r0 *1 0.47,0.56 nfet_01v8
M$7 6 10 8 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $9 r0 *1 1.31,0.56 nfet_01v8
M$9 13 5 8 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $10 r0 *1 1.73,0.56 nfet_01v8
M$10 12 4 13 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $11 r0 *1 2.21,0.56 nfet_01v8
M$11 10 3 12 11 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=126750000000P
+ PS=980000U PD=1040000U
* device instance $12 r0 *1 2.75,0.56 nfet_01v8
M$12 8 2 10 11 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=169000000000P
+ PS=1040000U PD=1820000U
.ENDS sky130_fd_sc_hd__a31o_2

* cell sky130_fd_sc_hd__a21bo_2
* pin VPB
* pin B1_N
* pin A1
* pin A2
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__a21bo_2 1 2 3 4 6 7 8 11
* net 1 VPB
* net 2 B1_N
* net 3 A1
* net 4 A2
* net 6 VPWR
* net 7 VGND
* net 8 X
* device instance $1 r0 *1 2.35,1.985 pfet_01v8_hvt
M$1 5 9 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.77,1.985 pfet_01v8_hvt
M$2 6 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 3.19,1.985 pfet_01v8_hvt
M$3 5 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $4 r0 *1 1.41,1.695 pfet_01v8_hvt
M$4 9 2 6 1 pfet_01v8_hvt L=150000U W=420000U AS=181500000000P AD=109200000000P
+ PS=1510000U PD=1360000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 8 10 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=400000000000P
+ AD=321500000000P PS=3800000U PD=2790000U
* device instance $7 r0 *1 2.35,0.56 nfet_01v8
M$7 10 9 7 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $8 r0 *1 2.83,0.56 nfet_01v8
M$8 12 3 10 11 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=68250000000P
+ PS=980000U PD=860000U
* device instance $9 r0 *1 3.19,0.56 nfet_01v8
M$9 7 4 12 11 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=169000000000P
+ PS=860000U PD=1820000U
* device instance $10 r0 *1 0.47,0.56 nfet_01v8
M$10 8 10 7 11 nfet_01v8 L=150000U W=1300000U AS=260000000000P AD=199375000000P
+ PS=2750000U PD=1940000U
* device instance $12 r0 *1 1.41,0.675 nfet_01v8
M$12 9 2 7 11 nfet_01v8 L=150000U W=420000U AS=108375000000P AD=109200000000P
+ PS=1010000U PD=1360000U
.ENDS sky130_fd_sc_hd__a21bo_2

* cell sky130_fd_sc_hd__a21boi_0
* pin VPB
* pin B1_N
* pin A1
* pin A2
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__a21boi_0 1 2 3 4 6 8 9 10
* net 1 VPB
* net 2 B1_N
* net 3 A1
* net 4 A2
* net 6 VGND
* net 8 VPWR
* net 9 Y
* device instance $1 r0 *1 1.425,2.165 pfet_01v8_hvt
M$1 5 7 9 1 pfet_01v8_hvt L=150000U W=640000U AS=169600000000P AD=89600000000P
+ PS=1810000U PD=920000U
* device instance $2 r0 *1 1.855,2.165 pfet_01v8_hvt
M$2 8 3 5 1 pfet_01v8_hvt L=150000U W=640000U AS=89600000000P AD=89600000000P
+ PS=920000U PD=920000U
* device instance $3 r0 *1 2.285,2.165 pfet_01v8_hvt
M$3 5 4 8 1 pfet_01v8_hvt L=150000U W=640000U AS=89600000000P AD=169600000000P
+ PS=920000U PD=1810000U
* device instance $4 r0 *1 0.475,2.275 pfet_01v8_hvt
M$4 8 2 7 1 pfet_01v8_hvt L=150000U W=420000U AS=111300000000P AD=111300000000P
+ PS=1370000U PD=1370000U
* device instance $5 r0 *1 0.475,0.445 nfet_01v8
M$5 6 2 7 10 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=130200000000P
+ PS=1370000U PD=1040000U
* device instance $6 r0 *1 1.245,0.445 nfet_01v8
M$6 9 7 6 10 nfet_01v8 L=150000U W=420000U AS=130200000000P AD=111300000000P
+ PS=1040000U PD=950000U
* device instance $7 r0 *1 1.925,0.445 nfet_01v8
M$7 11 3 9 10 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=44100000000P
+ PS=950000U PD=630000U
* device instance $8 r0 *1 2.285,0.445 nfet_01v8
M$8 6 4 11 10 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=111300000000P
+ PS=630000U PD=1370000U
.ENDS sky130_fd_sc_hd__a21boi_0

* cell sky130_fd_sc_hd__clkinv_2
* pin VPB
* pin A
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__clkinv_2 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 Y
* net 4 VPWR
* net 5 VGND
* device instance $1 r0 *1 0.495,1.985 pfet_01v8_hvt
M$1 4 2 3 1 pfet_01v8_hvt L=150000U W=3000000U AS=545000000000P
+ AD=545000000000P PS=5090000U PD=5090000U
* device instance $4 r0 *1 0.94,0.445 nfet_01v8
M$4 3 2 5 6 nfet_01v8 L=150000U W=840000U AS=170100000000P AD=168000000000P
+ PS=2070000U PD=2060000U
.ENDS sky130_fd_sc_hd__clkinv_2

* cell sky130_fd_sc_hd__or4_1
* pin VPB
* pin A
* pin B
* pin C
* pin D
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__or4_1 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 A
* net 3 B
* net 4 C
* net 5 D
* net 7 X
* net 8 VPWR
* net 9 VGND
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 13 5 6 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=69300000000P
+ PS=1360000U PD=750000U
* device instance $2 r0 *1 0.95,1.695 pfet_01v8_hvt
M$2 12 4 13 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=44100000000P
+ PS=750000U PD=630000U
* device instance $3 r0 *1 1.31,1.695 pfet_01v8_hvt
M$3 11 3 12 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $4 r0 *1 1.79,1.695 pfet_01v8_hvt
M$4 8 2 11 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=148250000000P
+ PS=750000U PD=1340000U
* device instance $5 r0 *1 2.28,1.985 pfet_01v8_hvt
M$5 7 6 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=148250000000P
+ AD=270000000000P PS=1340000U PD=2540000U
* device instance $6 r0 *1 0.47,0.475 nfet_01v8
M$6 6 5 9 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=69300000000P
+ PS=1360000U PD=750000U
* device instance $7 r0 *1 0.95,0.475 nfet_01v8
M$7 9 4 6 10 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=56700000000P
+ PS=750000U PD=690000U
* device instance $8 r0 *1 1.37,0.475 nfet_01v8
M$8 6 3 9 10 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $9 r0 *1 1.79,0.475 nfet_01v8
M$9 6 2 9 10 nfet_01v8 L=150000U W=420000U AS=101875000000P AD=56700000000P
+ PS=990000U PD=690000U
* device instance $10 r0 *1 2.28,0.56 nfet_01v8
M$10 7 6 9 10 nfet_01v8 L=150000U W=650000U AS=101875000000P AD=175500000000P
+ PS=990000U PD=1840000U
.ENDS sky130_fd_sc_hd__or4_1

* cell sky130_fd_sc_hd__o21bai_1
* pin VPB
* pin B1_N
* pin A1
* pin A2
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__o21bai_1 1 2 4 5 7 8 9 10
* net 1 VPB
* net 2 B1_N
* net 4 A1
* net 5 A2
* net 7 VPWR
* net 8 VGND
* net 9 Y
* device instance $1 r0 *1 0.86,1.97 pfet_01v8_hvt
M$1 3 2 7 1 pfet_01v8_hvt L=150000U W=420000U AS=178250000000P AD=109200000000P
+ PS=1400000U PD=1360000U
* device instance $2 r0 *1 1.41,1.985 pfet_01v8_hvt
M$2 9 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=178250000000P
+ AD=152500000000P PS=1400000U PD=1305000U
* device instance $3 r0 *1 1.865,1.985 pfet_01v8_hvt
M$3 11 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=127500000000P PS=1305000U PD=1255000U
* device instance $4 r0 *1 2.27,1.985 pfet_01v8_hvt
M$4 7 4 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=127500000000P
+ AD=280000000000P PS=1255000U PD=2560000U
* device instance $5 r0 *1 1.41,0.56 nfet_01v8
M$5 6 3 9 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=100750000000P
+ PS=1820000U PD=960000U
* device instance $6 r0 *1 1.87,0.56 nfet_01v8
M$6 8 5 6 10 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=87750000000P
+ PS=960000U PD=920000U
* device instance $7 r0 *1 2.29,0.56 nfet_01v8
M$7 6 4 8 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $8 r0 *1 0.47,0.675 nfet_01v8
M$8 3 2 8 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__o21bai_1

* cell sky130_fd_sc_hd__and4b_1
* pin VGND
* pin B
* pin C
* pin X
* pin A_N
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__and4b_1 1 4 5 6 7 8 12 13 14
* net 1 VGND
* net 4 B
* net 5 C
* net 6 X
* net 7 A_N
* net 8 D
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.47,2.275 pfet_01v8_hvt
M$1 12 7 2 13 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
* device instance $2 r0 *1 0.89,2.275 pfet_01v8_hvt
M$2 3 2 12 13 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P AD=98700000000P
+ PS=690000U PD=890000U
* device instance $3 r0 *1 1.51,2.275 pfet_01v8_hvt
M$3 12 4 3 13 pfet_01v8_hvt L=150000U W=420000U AS=98700000000P
+ AD=128100000000P PS=890000U PD=1030000U
* device instance $4 r0 *1 2.27,2.275 pfet_01v8_hvt
M$4 3 5 12 13 pfet_01v8_hvt L=150000U W=420000U AS=128100000000P
+ AD=66150000000P PS=1030000U PD=735000U
* device instance $5 r0 *1 2.735,2.275 pfet_01v8_hvt
M$5 3 8 12 13 pfet_01v8_hvt L=150000U W=420000U AS=140750000000P
+ AD=66150000000P PS=1325000U PD=735000U
* device instance $6 r0 *1 3.21,1.985 pfet_01v8_hvt
M$6 6 3 12 13 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $7 r0 *1 1.41,0.445 nfet_01v8
M$7 11 2 3 14 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $8 r0 *1 1.77,0.445 nfet_01v8
M$8 10 4 11 14 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=73500000000P
+ PS=630000U PD=770000U
* device instance $9 r0 *1 2.27,0.445 nfet_01v8
M$9 9 5 10 14 nfet_01v8 L=150000U W=420000U AS=73500000000P AD=60900000000P
+ PS=770000U PD=710000U
* device instance $10 r0 *1 2.71,0.445 nfet_01v8
M$10 1 8 9 14 nfet_01v8 L=150000U W=420000U AS=60900000000P AD=103400000000P
+ PS=710000U PD=1000000U
* device instance $11 r0 *1 3.21,0.56 nfet_01v8
M$11 6 3 1 14 nfet_01v8 L=150000U W=650000U AS=103400000000P AD=169000000000P
+ PS=1000000U PD=1820000U
* device instance $12 r0 *1 0.47,0.445 nfet_01v8
M$12 1 7 2 14 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__and4b_1

* cell sky130_fd_sc_hd__a32oi_1
* pin VPB
* pin B2
* pin B1
* pin A3
* pin A2
* pin A1
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a32oi_1 1 2 3 4 5 6 8 9 10 11
* net 1 VPB
* net 2 B2
* net 3 B1
* net 4 A3
* net 5 A2
* net 6 A1
* net 8 Y
* net 9 VGND
* net 10 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 7 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=215000000000P PS=1270000U PD=1430000U
* device instance $3 r0 *1 1.47,1.985 pfet_01v8_hvt
M$3 10 6 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=215000000000P
+ AD=135000000000P PS=1430000U PD=1270000U
* device instance $4 r0 *1 1.89,1.985 pfet_01v8_hvt
M$4 7 5 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=140000000000P PS=1270000U PD=1280000U
* device instance $5 r0 *1 2.32,1.985 pfet_01v8_hvt
M$5 10 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=260000000000P PS=1280000U PD=2520000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 14 2 9 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=74750000000P
+ PS=1820000U PD=880000U
* device instance $7 r0 *1 0.85,0.56 nfet_01v8
M$7 8 3 14 11 nfet_01v8 L=150000U W=650000U AS=74750000000P AD=152750000000P
+ PS=880000U PD=1120000U
* device instance $8 r0 *1 1.47,0.56 nfet_01v8
M$8 12 6 8 11 nfet_01v8 L=150000U W=650000U AS=152750000000P AD=71500000000P
+ PS=1120000U PD=870000U
* device instance $9 r0 *1 1.84,0.56 nfet_01v8
M$9 13 5 12 11 nfet_01v8 L=150000U W=650000U AS=71500000000P AD=107250000000P
+ PS=870000U PD=980000U
* device instance $10 r0 *1 2.32,0.56 nfet_01v8
M$10 9 4 13 11 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=169000000000P
+ PS=980000U PD=1820000U
.ENDS sky130_fd_sc_hd__a32oi_1

* cell sky130_fd_sc_hd__nand4b_4
* pin VGND
* pin D
* pin Y
* pin A_N
* pin B
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand4b_4 1 2 5 8 9 10 11 12 13
* net 1 VGND
* net 2 D
* net 5 Y
* net 8 A_N
* net 9 B
* net 10 C
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 11 8 3 12 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $2 r0 *1 1.41,1.985 pfet_01v8_hvt
M$2 5 3 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $6 r0 *1 3.09,1.985 pfet_01v8_hvt
M$6 5 9 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=800000000000P PS=5080000U PD=5600000U
* device instance $10 r0 *1 5.29,1.985 pfet_01v8_hvt
M$10 5 10 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=800000000000P
+ AD=540000000000P PS=5600000U PD=5080000U
* device instance $14 r0 *1 6.97,1.985 pfet_01v8_hvt
M$14 5 2 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $18 r0 *1 5.29,0.56 nfet_01v8
M$18 6 10 7 13 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $22 r0 *1 6.97,0.56 nfet_01v8
M$22 1 2 7 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $26 r0 *1 0.47,0.56 nfet_01v8
M$26 1 8 3 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
* device instance $27 r0 *1 1.41,0.56 nfet_01v8
M$27 5 3 4 13 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $31 r0 *1 3.09,0.56 nfet_01v8
M$31 6 9 4 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nand4b_4

* cell sky130_fd_sc_hd__a41oi_2
* pin VGND
* pin Y
* pin B1
* pin A1
* pin A2
* pin A3
* pin A4
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a41oi_2 1 2 6 7 8 9 10 12 13 14
* net 1 VGND
* net 2 Y
* net 6 B1
* net 7 A1
* net 8 A2
* net 9 A3
* net 10 A4
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 1.08,1.985 pfet_01v8_hvt
M$1 2 6 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.92,1.985 pfet_01v8_hvt
M$3 12 7 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $5 r0 *1 2.76,1.985 pfet_01v8_hvt
M$5 12 8 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=280000000000P PS=2540000U PD=2560000U
* device instance $7 r0 *1 3.62,1.985 pfet_01v8_hvt
M$7 12 9 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=530000000000P
+ AD=520000000000P PS=3060000U PD=3040000U
* device instance $9 r0 *1 4.96,1.985 pfet_01v8_hvt
M$9 12 10 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $11 r0 *1 4.12,0.56 nfet_01v8
M$11 4 9 5 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $13 r0 *1 4.96,0.56 nfet_01v8
M$13 1 10 5 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $15 r0 *1 1.92,0.56 nfet_01v8
M$15 2 7 3 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $17 r0 *1 2.76,0.56 nfet_01v8
M$17 4 8 3 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $19 r0 *1 0.56,0.56 nfet_01v8
M$19 2 6 1 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
.ENDS sky130_fd_sc_hd__a41oi_2

* cell sky130_fd_sc_hd__a2111oi_4
* pin VGND
* pin D1
* pin Y
* pin C1
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a2111oi_4 1 2 3 4 5 7 8 12 13 14
* net 1 VGND
* net 2 D1
* net 3 Y
* net 4 C1
* net 5 B1
* net 7 A1
* net 8 A2
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 4.44,1.985 pfet_01v8_hvt
M$1 11 5 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=680000000000P
+ AD=565000000000P PS=6360000U PD=5130000U
* device instance $5 r0 *1 6.17,1.985 pfet_01v8_hvt
M$5 12 7 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=575000000000P
+ AD=630000000000P PS=5150000U PD=5260000U
* device instance $9 r0 *1 8.03,1.985 pfet_01v8_hvt
M$9 12 8 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=730000000000P PS=5330000U PD=6460000U
* device instance $13 r0 *1 0.48,1.985 pfet_01v8_hvt
M$13 3 2 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=560000000000P PS=6370000U PD=5120000U
* device instance $17 r0 *1 2.2,1.985 pfet_01v8_hvt
M$17 11 4 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=560000000000P
+ AD=680000000000P PS=5120000U PD=6360000U
* device instance $21 r0 *1 6.38,0.56 nfet_01v8
M$21 3 7 6 14 nfet_01v8 L=150000U W=2600000U AS=455000000000P AD=394875000000P
+ PS=4650000U PD=3815000U
* device instance $25 r0 *1 8.195,0.56 nfet_01v8
M$25 1 8 6 14 nfet_01v8 L=150000U W=2600000U AS=394875000000P AD=445250000000P
+ PS=3815000U PD=4620000U
* device instance $29 r0 *1 0.49,0.56 nfet_01v8
M$29 3 2 1 14 nfet_01v8 L=150000U W=2600000U AS=451750000000P AD=386750000000P
+ PS=4640000U PD=3790000U
* device instance $33 r0 *1 2.28,0.56 nfet_01v8
M$33 3 4 1 14 nfet_01v8 L=150000U W=2600000U AS=390000000000P AD=399750000000P
+ PS=3800000U PD=3830000U
* device instance $37 r0 *1 4.11,0.56 nfet_01v8
M$37 3 5 1 14 nfet_01v8 L=150000U W=2600000U AS=399750000000P AD=455000000000P
+ PS=3830000U PD=4650000U
.ENDS sky130_fd_sc_hd__a2111oi_4

* cell sky130_fd_sc_hd__a2111oi_1
* pin VGND
* pin Y
* pin A2
* pin D1
* pin C1
* pin B1
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a2111oi_1 1 2 3 4 5 6 7 10 11 14
* net 1 VGND
* net 2 Y
* net 3 A2
* net 4 D1
* net 5 C1
* net 6 B1
* net 7 A1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.01,1.985 pfet_01v8_hvt
M$1 12 4 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=755000000000P
+ AD=172500000000P PS=3510000U PD=1345000U
* device instance $2 r0 *1 1.505,1.985 pfet_01v8_hvt
M$2 13 5 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=172500000000P
+ AD=185000000000P PS=1345000U PD=1370000U
* device instance $3 r0 *1 2.025,1.985 pfet_01v8_hvt
M$3 9 6 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=185000000000P
+ AD=290000000000P PS=1370000U PD=1580000U
* device instance $4 r0 *1 2.755,1.985 pfet_01v8_hvt
M$4 10 7 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=290000000000P
+ AD=137500000000P PS=1580000U PD=1275000U
* device instance $5 r0 *1 3.18,1.985 pfet_01v8_hvt
M$5 9 3 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=137500000000P
+ AD=290000000000P PS=1275000U PD=2580000U
* device instance $6 r0 *1 0.97,0.56 nfet_01v8
M$6 2 4 1 14 nfet_01v8 L=150000U W=650000U AS=481000000000P AD=125125000000P
+ PS=2780000U PD=1035000U
* device instance $7 r0 *1 1.505,0.56 nfet_01v8
M$7 1 5 2 14 nfet_01v8 L=150000U W=650000U AS=125125000000P AD=120250000000P
+ PS=1035000U PD=1020000U
* device instance $8 r0 *1 2.025,0.56 nfet_01v8
M$8 2 6 1 14 nfet_01v8 L=150000U W=650000U AS=120250000000P AD=191750000000P
+ PS=1020000U PD=1240000U
* device instance $9 r0 *1 2.765,0.56 nfet_01v8
M$9 8 7 2 14 nfet_01v8 L=150000U W=650000U AS=191750000000P AD=84500000000P
+ PS=1240000U PD=910000U
* device instance $10 r0 *1 3.175,0.56 nfet_01v8
M$10 1 3 8 14 nfet_01v8 L=150000U W=650000U AS=84500000000P AD=191750000000P
+ PS=910000U PD=1890000U
.ENDS sky130_fd_sc_hd__a2111oi_1

* cell sky130_fd_sc_hd__nor3b_1
* pin VPB
* pin B
* pin A
* pin C_N
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor3b_1 1 2 3 4 5 6 7 9
* net 1 VPB
* net 2 B
* net 3 A
* net 4 C_N
* net 5 Y
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 2.055,1.86 pfet_01v8_hvt
M$1 8 4 7 1 pfet_01v8_hvt L=150000U W=420000U AS=145750000000P AD=109200000000P
+ PS=1335000U PD=1360000U
* device instance $2 r0 *1 0.73,1.985 pfet_01v8_hvt
M$2 11 8 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=320000000000P
+ AD=135000000000P PS=2640000U PD=1270000U
* device instance $3 r0 *1 1.15,1.985 pfet_01v8_hvt
M$3 10 2 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $4 r0 *1 1.57,1.985 pfet_01v8_hvt
M$4 7 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=145750000000P PS=1270000U PD=1335000U
* device instance $5 r0 *1 0.73,0.56 nfet_01v8
M$5 6 8 5 9 nfet_01v8 L=150000U W=650000U AS=221000000000P AD=87750000000P
+ PS=1980000U PD=920000U
* device instance $6 r0 *1 1.15,0.56 nfet_01v8
M$6 5 2 6 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $7 r0 *1 1.57,0.56 nfet_01v8
M$7 6 3 5 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=100250000000P
+ PS=920000U PD=985000U
* device instance $8 r0 *1 2.055,0.675 nfet_01v8
M$8 8 4 6 9 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
.ENDS sky130_fd_sc_hd__nor3b_1

* cell sky130_fd_sc_hd__o31ai_2
* pin VGND
* pin A1
* pin A2
* pin A3
* pin Y
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o31ai_2 1 3 4 5 6 7 9 11 12
* net 1 VGND
* net 3 A1
* net 4 A2
* net 5 A3
* net 6 Y
* net 7 B1
* net 9 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.71,1.985 pfet_01v8_hvt
M$1 10 5 6 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 3.55,1.985 pfet_01v8_hvt
M$3 9 7 6 11 pfet_01v8_hvt L=150000U W=2000000U AS=330000000000P
+ AD=455000000000P PS=2660000U PD=3910000U
* device instance $5 r0 *1 0.49,1.985 pfet_01v8_hvt
M$5 9 3 8 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $7 r0 *1 1.33,1.985 pfet_01v8_hvt
M$7 10 4 8 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $9 r0 *1 0.49,0.56 nfet_01v8
M$9 1 3 2 12 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $11 r0 *1 1.33,0.56 nfet_01v8
M$11 1 4 2 12 nfet_01v8 L=150000U W=1300000U AS=286000000000P AD=325000000000P
+ PS=2180000U PD=2300000U
* device instance $13 r0 *1 2.63,0.56 nfet_01v8
M$13 1 5 2 12 nfet_01v8 L=150000U W=1300000U AS=240500000000P AD=201500000000P
+ PS=2040000U PD=1920000U
* device instance $15 r0 *1 3.55,0.56 nfet_01v8
M$15 6 7 2 12 nfet_01v8 L=150000U W=1300000U AS=214500000000P AD=295750000000P
+ PS=1960000U PD=2860000U
.ENDS sky130_fd_sc_hd__o31ai_2

* cell sky130_fd_sc_hd__xnor3_2
* pin VGND
* pin X
* pin C
* pin B
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__xnor3_2 1 2 6 11 12 13 14 15
* net 1 VGND
* net 2 X
* net 6 C
* net 11 B
* net 12 A
* net 13 VPWR
* net 14 VPB
* device instance $1 r0 *1 5.915,1.805 pfet_01v8_hvt
M$1 10 9 8 14 pfet_01v8_hvt L=150000U W=640000U AS=243100000000P
+ AD=246000000000P PS=1445000U PD=1525000U
* device instance $2 r0 *1 6.79,1.965 pfet_01v8_hvt
M$2 3 11 10 14 pfet_01v8_hvt L=150000U W=640000U AS=246000000000P
+ AD=145800000000P PS=1525000U PD=1205000U
* device instance $3 r0 *1 5.16,1.905 pfet_01v8_hvt
M$3 8 11 4 14 pfet_01v8_hvt L=150000U W=840000U AS=352800000000P
+ AD=243100000000P PS=2520000U PD=1445000U
* device instance $4 r0 *1 7.305,2.065 pfet_01v8_hvt
M$4 3 9 4 14 pfet_01v8_hvt L=150000U W=840000U AS=171500000000P
+ AD=145800000000P PS=1355000U PD=1205000U
* device instance $5 r0 *1 7.81,1.985 pfet_01v8_hvt
M$5 13 12 4 14 pfet_01v8_hvt L=150000U W=1000000U AS=171500000000P
+ AD=135000000000P PS=1355000U PD=1270000U
* device instance $6 r0 *1 8.23,1.985 pfet_01v8_hvt
M$6 10 4 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=285000000000P PS=1270000U PD=2570000U
* device instance $7 r0 *1 4.06,1.985 pfet_01v8_hvt
M$7 9 11 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=256550000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $8 r0 *1 1.465,1.805 pfet_01v8_hvt
M$8 7 6 13 14 pfet_01v8_hvt L=150000U W=640000U AS=169000000000P
+ AD=179200000000P PS=1365000U PD=1840000U
* device instance $9 r0 *1 0.53,1.985 pfet_01v8_hvt
M$9 2 5 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=455000000000P
+ AD=304000000000P PS=3910000U PD=2635000U
* device instance $11 r0 *1 3,1.905 pfet_01v8_hvt
M$11 8 7 5 14 pfet_01v8_hvt L=150000U W=840000U AS=152950000000P
+ AD=322350000000P PS=1315000U PD=2450000U
* device instance $12 r0 *1 2.515,2.045 pfet_01v8_hvt
M$12 3 6 5 14 pfet_01v8_hvt L=150000U W=840000U AS=152950000000P
+ AD=273000000000P PS=1315000U PD=2330000U
* device instance $13 r0 *1 5.915,0.455 nfet_01v8
M$13 10 9 3 15 nfet_01v8 L=150000U W=420000U AS=182050000000P AD=192650000000P
+ PS=1245000U PD=1285000U
* device instance $14 r0 *1 7.31,0.535 nfet_01v8
M$14 4 9 8 15 nfet_01v8 L=150000U W=600000U AS=140825000000P AD=110000000000P
+ PS=1100000U PD=990000U
* device instance $15 r0 *1 7.81,0.555 nfet_01v8
M$15 1 12 4 15 nfet_01v8 L=150000U W=640000U AS=110000000000P AD=86400000000P
+ PS=990000U PD=910000U
* device instance $16 r0 *1 8.23,0.555 nfet_01v8
M$16 10 4 1 15 nfet_01v8 L=150000U W=640000U AS=86400000000P AD=182400000000P
+ PS=910000U PD=1850000U
* device instance $17 r0 *1 5.16,0.565 nfet_01v8
M$17 3 11 4 15 nfet_01v8 L=150000U W=640000U AS=162750000000P AD=182050000000P
+ PS=1800000U PD=1245000U
* device instance $18 r0 *1 6.71,0.565 nfet_01v8
M$18 10 11 8 15 nfet_01v8 L=150000U W=640000U AS=140825000000P AD=192650000000P
+ PS=1100000U PD=1285000U
* device instance $19 r0 *1 0.51,0.56 nfet_01v8
M$19 2 5 1 15 nfet_01v8 L=150000U W=1300000U AS=282750000000P AD=204250000000P
+ PS=2820000U PD=1955000U
* device instance $21 r0 *1 1.465,0.675 nfet_01v8
M$21 7 6 1 15 nfet_01v8 L=150000U W=420000U AS=116500000000P AD=178500000000P
+ PS=1035000U PD=1690000U
* device instance $22 r0 *1 4.23,0.56 nfet_01v8
M$22 9 11 1 15 nfet_01v8 L=150000U W=650000U AS=188500000000P AD=165150000000P
+ PS=1880000U PD=1820000U
* device instance $23 r0 *1 2.58,0.565 nfet_01v8
M$23 5 6 8 15 nfet_01v8 L=150000U W=640000U AS=172800000000P AD=92800000000P
+ PS=1820000U PD=930000U
* device instance $24 r0 *1 3.02,0.565 nfet_01v8
M$24 3 7 5 15 nfet_01v8 L=150000U W=640000U AS=92800000000P AD=224000000000P
+ PS=930000U PD=1980000U
.ENDS sky130_fd_sc_hd__xnor3_2

* cell sky130_fd_sc_hd__o21a_4
* pin VGND
* pin X
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o21a_4 1 2 5 6 7 8 9 12
* net 1 VGND
* net 2 X
* net 5 B1
* net 6 A1
* net 7 A2
* net 8 VPWR
* net 9 VPB
* device instance $1 r0 *1 0.795,1.985 pfet_01v8_hvt
M$1 2 3 8 9 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=570000000000P PS=6370000U PD=5140000U
* device instance $5 r0 *1 2.535,1.985 pfet_01v8_hvt
M$5 3 5 8 9 pfet_01v8_hvt L=150000U W=2000000U AS=290000000000P
+ AD=450000000000P PS=2580000U PD=2900000U
* device instance $7 r0 *1 3.735,1.985 pfet_01v8_hvt
M$7 10 6 8 9 pfet_01v8_hvt L=150000U W=1000000U AS=310000000000P
+ AD=140000000000P PS=1620000U PD=1280000U
* device instance $8 r0 *1 4.165,1.985 pfet_01v8_hvt
M$8 3 7 10 9 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $9 r0 *1 4.595,1.985 pfet_01v8_hvt
M$9 11 7 3 9 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $10 r0 *1 5.025,1.985 pfet_01v8_hvt
M$10 8 6 11 9 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=285000000000P PS=1280000U PD=2570000U
* device instance $11 r0 *1 2.715,0.56 nfet_01v8
M$11 3 5 4 12 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=208000000000P
+ PS=2760000U PD=1940000U
* device instance $13 r0 *1 3.655,0.56 nfet_01v8
M$13 1 6 4 12 nfet_01v8 L=150000U W=1300000U AS=208000000000P AD=289250000000P
+ PS=1940000U PD=2840000U
* device instance $14 r0 *1 4.165,0.56 nfet_01v8
M$14 4 7 1 12 nfet_01v8 L=150000U W=1300000U AS=208000000000P AD=182000000000P
+ PS=1940000U PD=1860000U
* device instance $17 r0 *1 0.475,0.56 nfet_01v8
M$17 2 3 1 12 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=445250000000P
+ PS=4620000U PD=4620000U
.ENDS sky130_fd_sc_hd__o21a_4

* cell sky130_fd_sc_hd__o21a_2
* pin VPB
* pin B1
* pin A2
* pin A1
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__o21a_2 1 3 4 5 6 7 8 10
* net 1 VPB
* net 3 B1
* net 4 A2
* net 5 A1
* net 6 VGND
* net 7 VPWR
* net 8 X
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 2 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=397500000000P
+ AD=537500000000P PS=3795000U PD=3075000U
* device instance $3 r0 *1 1.845,1.985 pfet_01v8_hvt
M$3 2 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=400000000000P
+ AD=140000000000P PS=1800000U PD=1280000U
* device instance $4 r0 *1 2.275,1.985 pfet_01v8_hvt
M$4 11 4 2 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=160000000000P PS=1280000U PD=1320000U
* device instance $5 r0 *1 2.745,1.985 pfet_01v8_hvt
M$5 7 5 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=160000000000P
+ AD=265000000000P PS=1320000U PD=2530000U
* device instance $6 r0 *1 1.845,0.56 nfet_01v8
M$6 9 3 2 10 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=91000000000P
+ PS=1830000U PD=930000U
* device instance $7 r0 *1 2.275,0.56 nfet_01v8
M$7 6 4 9 10 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=104000000000P
+ PS=930000U PD=970000U
* device instance $8 r0 *1 2.745,0.56 nfet_01v8
M$8 9 5 6 10 nfet_01v8 L=150000U W=650000U AS=104000000000P AD=172250000000P
+ PS=970000U PD=1830000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 8 2 6 10 nfet_01v8 L=150000U W=1300000U AS=258375000000P AD=261625000000P
+ PS=2745000U PD=2755000U
.ENDS sky130_fd_sc_hd__o21a_2

* cell sky130_fd_sc_hd__or3_2
* pin VPB
* pin B
* pin A
* pin C
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__or3_2 1 2 3 4 5 6 7 9
* net 1 VPB
* net 2 B
* net 3 A
* net 4 C
* net 5 VPWR
* net 6 VGND
* net 7 X
* device instance $1 r0 *1 0.485,1.695 pfet_01v8_hvt
M$1 11 4 8 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 0.845,1.695 pfet_01v8_hvt
M$2 10 2 11 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $3 r0 *1 1.325,1.695 pfet_01v8_hvt
M$3 5 3 10 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=148250000000P
+ PS=750000U PD=1340000U
* device instance $4 r0 *1 1.815,1.985 pfet_01v8_hvt
M$4 7 8 5 1 pfet_01v8_hvt L=150000U W=2000000U AS=283250000000P
+ AD=450000000000P PS=2610000U PD=3900000U
* device instance $6 r0 *1 0.485,0.475 nfet_01v8
M$6 6 4 8 9 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $7 r0 *1 0.905,0.475 nfet_01v8
M$7 8 2 6 9 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $8 r0 *1 1.325,0.475 nfet_01v8
M$8 8 3 6 9 nfet_01v8 L=150000U W=420000U AS=101875000000P AD=56700000000P
+ PS=990000U PD=690000U
* device instance $9 r0 *1 1.815,0.56 nfet_01v8
M$9 7 8 6 9 nfet_01v8 L=150000U W=1300000U AS=189625000000P AD=273000000000P
+ PS=1910000U PD=2790000U
.ENDS sky130_fd_sc_hd__or3_2

* cell sky130_fd_sc_hd__nor2_8
* pin VGND
* pin A
* pin B
* pin Y
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor2_8 1 2 3 4 6 7 8
* net 1 VGND
* net 2 A
* net 3 B
* net 4 Y
* net 6 VPWR
* net 7 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 6 2 5 7 pfet_01v8_hvt L=150000U W=8000000U AS=1.225e+12P AD=1.08e+12P
+ PS=11450000U PD=10160000U
* device instance $9 r0 *1 3.85,1.985 pfet_01v8_hvt
M$9 4 3 5 7 pfet_01v8_hvt L=150000U W=8000000U AS=1.08e+12P AD=1.215e+12P
+ PS=10160000U PD=11430000U
* device instance $17 r0 *1 0.49,0.56 nfet_01v8
M$17 4 2 1 8 nfet_01v8 L=150000U W=5200000U AS=796250000000P AD=702000000000P
+ PS=8300000U PD=7360000U
* device instance $25 r0 *1 3.85,0.56 nfet_01v8
M$25 4 3 1 8 nfet_01v8 L=150000U W=5200000U AS=702000000000P AD=783250000000P
+ PS=7360000U PD=8260000U
.ENDS sky130_fd_sc_hd__nor2_8

* cell sky130_fd_sc_hd__o41a_1
* pin VGND
* pin X
* pin B1
* pin A4
* pin A3
* pin A2
* pin A1
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o41a_1 1 2 5 6 7 8 9 10 11 15
* net 1 VGND
* net 2 X
* net 5 B1
* net 6 A4
* net 7 A3
* net 8 A2
* net 9 A1
* net 10 VPB
* net 11 VPWR
* device instance $1 r0 *1 0.8,1.985 pfet_01v8_hvt
M$1 11 3 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=425000000000P
+ AD=135000000000P PS=2850000U PD=1270000U
* device instance $2 r0 *1 1.22,1.985 pfet_01v8_hvt
M$2 3 5 11 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=1520000U
* device instance $3 r0 *1 1.89,1.985 pfet_01v8_hvt
M$3 12 6 3 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=220000000000P PS=1520000U PD=1440000U
* device instance $4 r0 *1 2.48,1.985 pfet_01v8_hvt
M$4 13 7 12 10 pfet_01v8_hvt L=150000U W=1000000U AS=220000000000P
+ AD=195000000000P PS=1440000U PD=1390000U
* device instance $5 r0 *1 3.02,1.985 pfet_01v8_hvt
M$5 14 8 13 10 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=195000000000P PS=1390000U PD=1390000U
* device instance $6 r0 *1 3.56,1.985 pfet_01v8_hvt
M$6 11 9 14 10 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=280000000000P PS=1390000U PD=2560000U
* device instance $7 r0 *1 1.53,0.56 nfet_01v8
M$7 4 5 3 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 1.95,0.56 nfet_01v8
M$8 1 6 4 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=123500000000P
+ PS=920000U PD=1030000U
* device instance $9 r0 *1 2.48,0.56 nfet_01v8
M$9 4 7 1 15 nfet_01v8 L=150000U W=650000U AS=123500000000P AD=126750000000P
+ PS=1030000U PD=1040000U
* device instance $10 r0 *1 3.02,0.56 nfet_01v8
M$10 1 8 4 15 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=126750000000P
+ PS=1040000U PD=1040000U
* device instance $11 r0 *1 3.56,0.56 nfet_01v8
M$11 4 9 1 15 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=195000000000P
+ PS=1040000U PD=1900000U
* device instance $12 r0 *1 0.59,0.56 nfet_01v8
M$12 1 3 2 15 nfet_01v8 L=150000U W=650000U AS=247000000000P AD=169000000000P
+ PS=2060000U PD=1820000U
.ENDS sky130_fd_sc_hd__o41a_1

* cell sky130_fd_sc_hd__inv_6
* pin VPB
* pin A
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__inv_6 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 Y
* net 4 VPWR
* net 5 VGND
* device instance $1 r0 *1 0.64,1.985 pfet_01v8_hvt
M$1 3 2 4 1 pfet_01v8_hvt L=150000U W=6000000U AS=1.105e+12P AD=945000000000P
+ PS=9210000U PD=8890000U
* device instance $7 r0 *1 0.64,0.56 nfet_01v8
M$7 3 2 5 6 nfet_01v8 L=150000U W=3900000U AS=685750000000P AD=614250000000P
+ PS=6660000U PD=6440000U
.ENDS sky130_fd_sc_hd__inv_6

* cell sky130_fd_sc_hd__mux2_2
* pin VGND
* pin X
* pin A0
* pin A1
* pin S
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2_2 1 2 4 5 6 10 11 14
* net 1 VGND
* net 2 X
* net 4 A0
* net 5 A1
* net 6 S
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 2 3 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=312800000000P PS=3790000U PD=2685000U
* device instance $3 r0 *1 1.455,2.165 pfet_01v8_hvt
M$3 12 9 10 11 pfet_01v8_hvt L=150000U W=640000U AS=177800000000P
+ AD=228800000000P PS=1415000U PD=1355000U
* device instance $4 r0 *1 2.32,2.165 pfet_01v8_hvt
M$4 3 5 12 11 pfet_01v8_hvt L=150000U W=640000U AS=228800000000P
+ AD=131200000000P PS=1355000U PD=1050000U
* device instance $5 r0 *1 2.88,2.165 pfet_01v8_hvt
M$5 13 4 3 11 pfet_01v8_hvt L=150000U W=640000U AS=131200000000P
+ AD=67200000000P PS=1050000U PD=850000U
* device instance $6 r0 *1 3.24,2.165 pfet_01v8_hvt
M$6 10 6 13 11 pfet_01v8_hvt L=150000U W=640000U AS=67200000000P
+ AD=86400000000P PS=850000U PD=910000U
* device instance $7 r0 *1 3.66,2.165 pfet_01v8_hvt
M$7 9 6 10 11 pfet_01v8_hvt L=150000U W=640000U AS=86400000000P
+ AD=172800000000P PS=910000U PD=1820000U
* device instance $8 r0 *1 1.365,0.445 nfet_01v8
M$8 7 9 1 14 nfet_01v8 L=150000U W=420000U AS=97000000000P AD=68250000000P
+ PS=975000U PD=745000U
* device instance $9 r0 *1 1.84,0.445 nfet_01v8
M$9 3 4 7 14 nfet_01v8 L=150000U W=420000U AS=68250000000P AD=173250000000P
+ PS=745000U PD=1245000U
* device instance $10 r0 *1 2.815,0.445 nfet_01v8
M$10 8 5 3 14 nfet_01v8 L=150000U W=420000U AS=173250000000P AD=57750000000P
+ PS=1245000U PD=695000U
* device instance $11 r0 *1 3.24,0.445 nfet_01v8
M$11 1 6 8 14 nfet_01v8 L=150000U W=420000U AS=57750000000P AD=56700000000P
+ PS=695000U PD=690000U
* device instance $12 r0 *1 3.66,0.445 nfet_01v8
M$12 9 6 1 14 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=113400000000P
+ PS=690000U PD=1380000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 2 3 1 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=184750000000P
+ PS=2740000U PD=1895000U
.ENDS sky130_fd_sc_hd__mux2_2

* cell sky130_fd_sc_hd__o311ai_1
* pin VGND
* pin Y
* pin A1
* pin A2
* pin A3
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311ai_1 1 3 4 5 6 7 8 10 11 14
* net 1 VGND
* net 3 Y
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 B1
* net 8 C1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.615,1.985 pfet_01v8_hvt
M$1 12 4 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=135000000000P PS=2560000U PD=1270000U
* device instance $2 r0 *1 1.035,1.985 pfet_01v8_hvt
M$2 13 5 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 1.455,1.985 pfet_01v8_hvt
M$3 3 6 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=225000000000P PS=1270000U PD=1450000U
* device instance $4 r0 *1 2.055,1.985 pfet_01v8_hvt
M$4 10 7 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=225000000000P
+ AD=185000000000P PS=1450000U PD=1370000U
* device instance $5 r0 *1 2.575,1.985 pfet_01v8_hvt
M$5 3 8 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=185000000000P
+ AD=310000000000P PS=1370000U PD=2620000U
* device instance $6 r0 *1 0.615,0.56 nfet_01v8
M$6 2 4 1 14 nfet_01v8 L=150000U W=650000U AS=182000000000P AD=87750000000P
+ PS=1860000U PD=920000U
* device instance $7 r0 *1 1.035,0.56 nfet_01v8
M$7 1 5 2 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $8 r0 *1 1.455,0.56 nfet_01v8
M$8 2 6 1 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=198250000000P
+ PS=920000U PD=1260000U
* device instance $9 r0 *1 2.215,0.56 nfet_01v8
M$9 9 7 2 14 nfet_01v8 L=150000U W=650000U AS=198250000000P AD=68250000000P
+ PS=1260000U PD=860000U
* device instance $10 r0 *1 2.575,0.56 nfet_01v8
M$10 3 8 9 14 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=182000000000P
+ PS=860000U PD=1860000U
.ENDS sky130_fd_sc_hd__o311ai_1

* cell sky130_fd_sc_hd__o2bb2ai_2
* pin VGND
* pin A1_N
* pin A2_N
* pin Y
* pin B1
* pin B2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 1 2 4 7 8 9 10 12 13
* net 1 VGND
* net 2 A1_N
* net 4 A2_N
* net 7 Y
* net 8 B1
* net 9 B2
* net 10 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 5 2 10 12 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=535000000000P PS=3830000U PD=3070000U
* device instance $2 r0 *1 0.91,1.985 pfet_01v8_hvt
M$2 10 4 5 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $5 r0 *1 2.7,1.985 pfet_01v8_hvt
M$5 7 5 10 12 pfet_01v8_hvt L=150000U W=2000000U AS=535000000000P
+ AD=287500000000P PS=3070000U PD=2575000U
* device instance $7 r0 *1 3.575,1.985 pfet_01v8_hvt
M$7 11 8 10 12 pfet_01v8_hvt L=150000U W=2000000U AS=287500000000P
+ AD=420000000000P PS=2575000U PD=3840000U
* device instance $8 r0 *1 3.995,1.985 pfet_01v8_hvt
M$8 7 9 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $11 r0 *1 2.7,0.56 nfet_01v8
M$11 7 5 6 13 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=186875000000P
+ PS=2760000U PD=1875000U
* device instance $13 r0 *1 3.575,0.56 nfet_01v8
M$13 1 8 6 13 nfet_01v8 L=150000U W=1300000U AS=186875000000P AD=256750000000P
+ PS=1875000U PD=2740000U
* device instance $14 r0 *1 3.995,0.56 nfet_01v8
M$14 6 9 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $17 r0 *1 0.49,0.56 nfet_01v8
M$17 3 2 1 13 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=256750000000P
+ PS=2780000U PD=2740000U
* device instance $18 r0 *1 0.91,0.56 nfet_01v8
M$18 5 4 3 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
.ENDS sky130_fd_sc_hd__o2bb2ai_2

* cell sky130_fd_sc_hd__a211o_2
* pin VGND
* pin X
* pin A2
* pin A1
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a211o_2 1 2 5 6 7 8 9 11 12
* net 1 VGND
* net 2 X
* net 5 A2
* net 6 A1
* net 7 B1
* net 8 C1
* net 9 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.83,1.985 pfet_01v8_hvt
M$1 9 5 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=195000000000P PS=2520000U PD=1390000U
* device instance $2 r0 *1 2.37,1.985 pfet_01v8_hvt
M$2 10 6 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=165000000000P PS=1390000U PD=1330000U
* device instance $3 r0 *1 2.85,1.985 pfet_01v8_hvt
M$3 13 7 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=105000000000P PS=1330000U PD=1210000U
* device instance $4 r0 *1 3.21,1.985 pfet_01v8_hvt
M$4 3 8 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 2 3 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $7 r0 *1 0.47,0.56 nfet_01v8
M$7 2 3 1 12 nfet_01v8 L=150000U W=1300000U AS=260000000000P AD=290875000000P
+ PS=2750000U PD=2195000U
* device instance $9 r0 *1 1.665,0.56 nfet_01v8
M$9 4 5 1 12 nfet_01v8 L=150000U W=650000U AS=199875000000P AD=133250000000P
+ PS=1265000U PD=1060000U
* device instance $10 r0 *1 2.225,0.56 nfet_01v8
M$10 3 6 4 12 nfet_01v8 L=150000U W=650000U AS=133250000000P AD=115375000000P
+ PS=1060000U PD=1005000U
* device instance $11 r0 *1 2.73,0.56 nfet_01v8
M$11 1 7 3 12 nfet_01v8 L=150000U W=650000U AS=115375000000P AD=107250000000P
+ PS=1005000U PD=980000U
* device instance $12 r0 *1 3.21,0.56 nfet_01v8
M$12 3 8 1 12 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=169000000000P
+ PS=980000U PD=1820000U
.ENDS sky130_fd_sc_hd__a211o_2

* cell sky130_fd_sc_hd__nand2b_1
* pin VPB
* pin B
* pin A_N
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nand2b_1 1 2 4 5 6 7 8
* net 1 VPB
* net 2 B
* net 4 A_N
* net 5 Y
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 7 4 3 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=145750000000P
+ PS=1360000U PD=1335000U
* device instance $2 r0 *1 0.955,1.985 pfet_01v8_hvt
M$2 5 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=145750000000P
+ AD=135000000000P PS=1335000U PD=1270000U
* device instance $3 r0 *1 1.375,1.985 pfet_01v8_hvt
M$3 7 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=265000000000P PS=1270000U PD=2530000U
* device instance $4 r0 *1 0.47,0.675 nfet_01v8
M$4 3 4 6 8 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
* device instance $5 r0 *1 0.955,0.56 nfet_01v8
M$5 9 2 6 8 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=87750000000P
+ PS=985000U PD=920000U
* device instance $6 r0 *1 1.375,0.56 nfet_01v8
M$6 5 3 9 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2b_1

* cell sky130_fd_sc_hd__clkinv_4
* pin VPB
* pin A
* pin VGND
* pin Y
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__clkinv_4 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 VGND
* net 4 Y
* net 5 VPWR
* device instance $1 r0 *1 0.515,1.985 pfet_01v8_hvt
M$1 4 2 5 1 pfet_01v8_hvt L=150000U W=6000000U AS=1.005e+12P AD=1.045e+12P
+ PS=9010000U PD=9090000U
* device instance $7 r0 *1 0.945,0.445 nfet_01v8
M$7 4 2 3 6 nfet_01v8 L=150000U W=1680000U AS=315000000000P AD=342300000000P
+ PS=3600000U PD=3730000U
.ENDS sky130_fd_sc_hd__clkinv_4

* cell sky130_fd_sc_hd__o2111ai_4
* pin VGND
* pin D1
* pin A2
* pin Y
* pin C1
* pin B1
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o2111ai_4 1 2 3 4 6 9 10 11 13 14
* net 1 VGND
* net 2 D1
* net 3 A2
* net 4 Y
* net 6 C1
* net 9 B1
* net 10 A1
* net 11 VPWR
* net 13 VPB
* device instance $1 r0 *1 7.93,1.985 pfet_01v8_hvt
M$1 12 10 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=657850000000P
+ AD=665000000000P PS=6330000U PD=6330000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 11 2 4 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $9 r0 *1 2.15,1.985 pfet_01v8_hvt
M$9 11 6 4 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=642500000000P PS=5080000U PD=5285000U
* device instance $13 r0 *1 4.035,1.985 pfet_01v8_hvt
M$13 11 9 4 13 pfet_01v8_hvt L=150000U W=4000000U AS=642500000000P
+ AD=552500000000P PS=5285000U PD=5105000U
* device instance $17 r0 *1 5.74,1.985 pfet_01v8_hvt
M$17 12 3 4 13 pfet_01v8_hvt L=150000U W=4000000U AS=552500000000P
+ AD=658350000000P PS=5105000U PD=6330000U
* device instance $21 r0 *1 4.35,0.56 nfet_01v8
M$21 7 9 8 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=359125000000P
+ PS=4580000U PD=3705000U
* device instance $25 r0 *1 6.055,0.56 nfet_01v8
M$25 1 3 8 14 nfet_01v8 L=150000U W=2600000U AS=365625000000P AD=365625000000P
+ PS=3725000U PD=3725000U
* device instance $29 r0 *1 7.78,0.56 nfet_01v8
M$29 1 10 8 14 nfet_01v8 L=150000U W=2600000U AS=359125000000P AD=448500000000P
+ PS=3705000U PD=4630000U
* device instance $33 r0 *1 0.47,0.56 nfet_01v8
M$33 4 2 5 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $37 r0 *1 2.15,0.56 nfet_01v8
M$37 7 6 5 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__o2111ai_4

* cell sky130_fd_sc_hd__a32o_2
* pin VGND
* pin X
* pin A1
* pin A2
* pin B2
* pin B1
* pin A3
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a32o_2 1 2 4 5 6 7 8 13 14 15
* net 1 VGND
* net 2 X
* net 4 A1
* net 5 A2
* net 6 B2
* net 7 B1
* net 8 A3
* net 13 VPWR
* net 14 VPB
* device instance $1 r0 *1 1.83,1.985 pfet_01v8_hvt
M$1 3 6 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 2.25,1.985 pfet_01v8_hvt
M$2 12 7 3 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 2.67,1.985 pfet_01v8_hvt
M$3 13 4 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=215000000000P PS=1270000U PD=1430000U
* device instance $4 r0 *1 3.25,1.985 pfet_01v8_hvt
M$4 12 5 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=215000000000P
+ AD=135000000000P PS=1430000U PD=1270000U
* device instance $5 r0 *1 3.67,1.985 pfet_01v8_hvt
M$5 13 8 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $6 r0 *1 0.47,1.985 pfet_01v8_hvt
M$6 13 3 2 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $8 r0 *1 0.47,0.56 nfet_01v8
M$8 2 3 1 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=297375000000P
+ PS=2740000U PD=2215000U
* device instance $10 r0 *1 1.685,0.56 nfet_01v8
M$10 11 6 1 15 nfet_01v8 L=150000U W=650000U AS=209625000000P AD=115375000000P
+ PS=1295000U PD=1005000U
* device instance $11 r0 *1 2.19,0.56 nfet_01v8
M$11 3 7 11 15 nfet_01v8 L=150000U W=650000U AS=115375000000P AD=107250000000P
+ PS=1005000U PD=980000U
* device instance $12 r0 *1 2.67,0.56 nfet_01v8
M$12 10 4 3 15 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=139750000000P
+ PS=980000U PD=1080000U
* device instance $13 r0 *1 3.25,0.56 nfet_01v8
M$13 9 5 10 15 nfet_01v8 L=150000U W=650000U AS=139750000000P AD=87750000000P
+ PS=1080000U PD=920000U
* device instance $14 r0 *1 3.67,0.56 nfet_01v8
M$14 1 8 9 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a32o_2

* cell sky130_fd_sc_hd__a221oi_2
* pin VGND
* pin C1
* pin Y
* pin B2
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a221oi_2 1 2 3 4 6 7 9 10 11 14
* net 1 VGND
* net 2 C1
* net 3 Y
* net 4 B2
* net 6 B1
* net 7 A2
* net 9 A1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.84,1.985 pfet_01v8_hvt
M$1 12 4 13 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=310000000000P PS=3790000U PD=2620000U
* device instance $2 r0 *1 2.26,1.985 pfet_01v8_hvt
M$2 13 6 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $5 r0 *1 3.6,1.985 pfet_01v8_hvt
M$5 10 7 13 11 pfet_01v8_hvt L=150000U W=2000000U AS=310000000000P
+ AD=420000000000P PS=2620000U PD=3840000U
* device instance $6 r0 *1 4.02,1.985 pfet_01v8_hvt
M$6 13 9 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $9 r0 *1 0.48,1.985 pfet_01v8_hvt
M$9 3 2 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=395000000000P PS=3810000U PD=3790000U
* device instance $11 r0 *1 0.48,0.56 nfet_01v8
M$11 3 2 1 14 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=344500000000P
+ PS=2760000U PD=2360000U
* device instance $13 r0 *1 1.84,0.56 nfet_01v8
M$13 5 4 1 14 nfet_01v8 L=150000U W=1300000U AS=344500000000P AD=201500000000P
+ PS=2360000U PD=1920000U
* device instance $14 r0 *1 2.26,0.56 nfet_01v8
M$14 3 6 5 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $17 r0 *1 3.6,0.56 nfet_01v8
M$17 8 7 1 14 nfet_01v8 L=150000U W=1300000U AS=201500000000P AD=256750000000P
+ PS=1920000U PD=2740000U
* device instance $18 r0 *1 4.02,0.56 nfet_01v8
M$18 3 9 8 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
.ENDS sky130_fd_sc_hd__a221oi_2

* cell sky130_fd_sc_hd__or2_2
* pin VPB
* pin A
* pin B
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__or2_2 1 2 4 5 6 7 8
* net 1 VPB
* net 2 A
* net 4 B
* net 5 X
* net 6 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.53,1.695 pfet_01v8_hvt
M$1 9 4 3 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 0.89,1.695 pfet_01v8_hvt
M$2 6 2 9 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=155750000000P
+ PS=630000U PD=1355000U
* device instance $3 r0 *1 1.395,1.985 pfet_01v8_hvt
M$3 5 3 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=290750000000P
+ AD=395000000000P PS=2625000U PD=3790000U
* device instance $5 r0 *1 0.47,0.445 nfet_01v8
M$5 3 4 7 8 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $6 r0 *1 0.89,0.445 nfet_01v8
M$6 7 2 3 8 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=106750000000P
+ PS=690000U PD=1005000U
* device instance $7 r0 *1 1.395,0.56 nfet_01v8
M$7 5 3 7 8 nfet_01v8 L=150000U W=1300000U AS=194500000000P AD=256750000000P
+ PS=1925000U PD=2740000U
.ENDS sky130_fd_sc_hd__or2_2

* cell sky130_fd_sc_hd__nand3_4
* pin VGND
* pin C
* pin B
* pin A
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand3_4 1 2 5 6 7 8 9 10
* net 1 VGND
* net 2 C
* net 5 B
* net 6 A
* net 7 VPWR
* net 8 Y
* net 9 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 2 7 9 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 8 5 7 9 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $9 r0 *1 4.35,1.985 pfet_01v8_hvt
M$9 8 6 7 9 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=675000000000P PS=6330000U PD=6350000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 1 2 3 10 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $17 r0 *1 2.15,0.56 nfet_01v8
M$17 4 5 3 10 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $21 r0 *1 4.35,0.56 nfet_01v8
M$21 8 6 4 10 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=438750000000P
+ PS=4580000U PD=4600000U
.ENDS sky130_fd_sc_hd__nand3_4

* cell sky130_fd_sc_hd__o32a_4
* pin VGND
* pin A1
* pin A2
* pin A3
* pin B1
* pin B2
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o32a_4 1 3 4 5 7 8 9 11 14 15
* net 1 VGND
* net 3 A1
* net 4 A2
* net 5 A3
* net 7 B1
* net 8 B2
* net 9 X
* net 11 VPWR
* net 14 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 11 3 10 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 12 4 10 14 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 4.03,1.985 pfet_01v8_hvt
M$5 11 7 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $7 r0 *1 4.87,1.985 pfet_01v8_hvt
M$7 6 8 13 14 pfet_01v8_hvt L=150000U W=2000000U AS=285000000000P
+ AD=410000000000P PS=2570000U PD=3820000U
* device instance $9 r0 *1 6.26,1.985 pfet_01v8_hvt
M$9 9 6 11 14 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=665000000000P PS=6330000U PD=6330000U
* device instance $13 r0 *1 2.67,1.985 pfet_01v8_hvt
M$13 6 5 12 14 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $15 r0 *1 6.26,0.56 nfet_01v8
M$15 9 6 1 15 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
* device instance $19 r0 *1 0.47,0.56 nfet_01v8
M$19 1 3 2 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $21 r0 *1 1.31,0.56 nfet_01v8
M$21 1 4 2 15 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=182000000000P
+ PS=1840000U PD=1860000U
* device instance $23 r0 *1 2.17,0.56 nfet_01v8
M$23 1 5 2 15 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=256750000000P
+ PS=1860000U PD=2740000U
* device instance $25 r0 *1 4.03,0.56 nfet_01v8
M$25 2 7 6 15 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $27 r0 *1 4.87,0.56 nfet_01v8
M$27 2 8 6 15 nfet_01v8 L=150000U W=1300000U AS=185250000000P AD=266500000000P
+ PS=1870000U PD=2770000U
.ENDS sky130_fd_sc_hd__o32a_4

* cell sky130_fd_sc_hd__o311a_1
* pin VGND
* pin X
* pin A1
* pin A2
* pin A3
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311a_1 1 2 5 6 7 8 9 11 12 15
* net 1 VGND
* net 2 X
* net 5 A1
* net 6 A2
* net 7 A3
* net 8 B1
* net 9 C1
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.48,1.985 pfet_01v8_hvt
M$1 11 4 2 12 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=312500000000P PS=2520000U PD=1625000U
* device instance $2 r0 *1 1.255,1.985 pfet_01v8_hvt
M$2 14 5 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=312500000000P
+ AD=180000000000P PS=1625000U PD=1360000U
* device instance $3 r0 *1 1.765,1.985 pfet_01v8_hvt
M$3 13 6 14 12 pfet_01v8_hvt L=150000U W=1000000U AS=180000000000P
+ AD=210000000000P PS=1360000U PD=1420000U
* device instance $4 r0 *1 2.335,1.985 pfet_01v8_hvt
M$4 4 7 13 12 pfet_01v8_hvt L=150000U W=1000000U AS=210000000000P
+ AD=137500000000P PS=1420000U PD=1275000U
* device instance $5 r0 *1 2.76,1.985 pfet_01v8_hvt
M$5 11 8 4 12 pfet_01v8_hvt L=150000U W=1000000U AS=137500000000P
+ AD=150000000000P PS=1275000U PD=1300000U
* device instance $6 r0 *1 3.21,1.985 pfet_01v8_hvt
M$6 4 9 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=150000000000P
+ AD=260000000000P PS=1300000U PD=2520000U
* device instance $7 r0 *1 0.48,0.56 nfet_01v8
M$7 1 4 2 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=203125000000P
+ PS=1820000U PD=1275000U
* device instance $8 r0 *1 1.255,0.56 nfet_01v8
M$8 3 5 1 15 nfet_01v8 L=150000U W=650000U AS=203125000000P AD=117000000000P
+ PS=1275000U PD=1010000U
* device instance $9 r0 *1 1.765,0.56 nfet_01v8
M$9 1 6 3 15 nfet_01v8 L=150000U W=650000U AS=117000000000P AD=136500000000P
+ PS=1010000U PD=1070000U
* device instance $10 r0 *1 2.335,0.56 nfet_01v8
M$10 3 7 1 15 nfet_01v8 L=150000U W=650000U AS=136500000000P AD=118625000000P
+ PS=1070000U PD=1015000U
* device instance $11 r0 *1 2.85,0.56 nfet_01v8
M$11 10 8 3 15 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=68250000000P
+ PS=1015000U PD=860000U
* device instance $12 r0 *1 3.21,0.56 nfet_01v8
M$12 4 9 10 15 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=169000000000P
+ PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o311a_1

* cell sky130_fd_sc_hd__o21a_1
* pin VPB
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o21a_1 1 2 3 4 5 7 8 10
* net 1 VPB
* net 2 B1
* net 3 A2
* net 4 A1
* net 5 VPWR
* net 7 X
* net 8 VGND
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 5 9 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=327500000000P PS=2560000U PD=1655000U
* device instance $2 r0 *1 1.295,1.985 pfet_01v8_hvt
M$2 9 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=327500000000P
+ AD=195000000000P PS=1655000U PD=1390000U
* device instance $3 r0 *1 1.835,1.985 pfet_01v8_hvt
M$3 11 3 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=152500000000P PS=1390000U PD=1305000U
* device instance $4 r0 *1 2.29,1.985 pfet_01v8_hvt
M$4 5 4 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=260000000000P PS=1305000U PD=2520000U
* device instance $5 r0 *1 1.41,0.56 nfet_01v8
M$5 6 2 9 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=100750000000P
+ PS=1820000U PD=960000U
* device instance $6 r0 *1 1.87,0.56 nfet_01v8
M$6 8 3 6 10 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=87750000000P
+ PS=960000U PD=920000U
* device instance $7 r0 *1 2.29,0.56 nfet_01v8
M$7 6 4 8 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $8 r0 *1 0.47,0.56 nfet_01v8
M$8 8 9 7 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__o21a_1

* cell sky130_fd_sc_hd__nor2_4
* pin VGND
* pin B
* pin Y
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor2_4 1 2 3 4 6 7 8
* net 1 VGND
* net 2 B
* net 3 Y
* net 4 A
* net 6 VPWR
* net 7 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 6 4 5 7 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $5 r0 *1 2.17,1.985 pfet_01v8_hvt
M$5 3 2 5 7 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=675000000000P PS=5080000U PD=6350000U
* device instance $9 r0 *1 0.49,0.56 nfet_01v8
M$9 3 4 1 8 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $13 r0 *1 2.17,0.56 nfet_01v8
M$13 3 2 1 8 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nor2_4

* cell sky130_fd_sc_hd__o2111ai_1
* pin VPB
* pin D1
* pin C1
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o2111ai_1 1 2 3 4 5 6 8 9 10 11
* net 1 VPB
* net 2 D1
* net 3 C1
* net 4 B1
* net 5 A2
* net 6 A1
* net 8 VPWR
* net 9 Y
* net 10 VGND
* device instance $1 r0 *1 0.67,1.985 pfet_01v8_hvt
M$1 9 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 1.1,1.985 pfet_01v8_hvt
M$2 8 3 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=195000000000P PS=1280000U PD=1390000U
* device instance $3 r0 *1 1.64,1.985 pfet_01v8_hvt
M$3 9 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=202500000000P PS=1390000U PD=1405000U
* device instance $4 r0 *1 2.195,1.985 pfet_01v8_hvt
M$4 12 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=202500000000P
+ AD=195000000000P PS=1405000U PD=1390000U
* device instance $5 r0 *1 2.735,1.985 pfet_01v8_hvt
M$5 8 6 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=265000000000P PS=1390000U PD=2530000U
* device instance $6 r0 *1 0.74,0.56 nfet_01v8
M$6 14 2 9 11 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=68250000000P
+ PS=1830000U PD=860000U
* device instance $7 r0 *1 1.1,0.56 nfet_01v8
M$7 13 3 14 11 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=126750000000P
+ PS=860000U PD=1040000U
* device instance $8 r0 *1 1.64,0.56 nfet_01v8
M$8 7 4 13 11 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=131625000000P
+ PS=1040000U PD=1055000U
* device instance $9 r0 *1 2.195,0.56 nfet_01v8
M$9 10 5 7 11 nfet_01v8 L=150000U W=650000U AS=131625000000P AD=126750000000P
+ PS=1055000U PD=1040000U
* device instance $10 r0 *1 2.735,0.56 nfet_01v8
M$10 7 6 10 11 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=172250000000P
+ PS=1040000U PD=1830000U
.ENDS sky130_fd_sc_hd__o2111ai_1

* cell sky130_fd_sc_hd__o211a_2
* pin VPB
* pin C1
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__o211a_2 1 2 3 4 5 7 9 10 11
* net 1 VPB
* net 2 C1
* net 3 B1
* net 4 A2
* net 5 A1
* net 7 VPWR
* net 9 VGND
* net 10 X
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 7 2 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 0.905,1.985 pfet_01v8_hvt
M$2 6 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=367500000000P PS=1280000U PD=1735000U
* device instance $3 r0 *1 1.79,1.985 pfet_01v8_hvt
M$3 12 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=367500000000P
+ AD=105000000000P PS=1735000U PD=1210000U
* device instance $4 r0 *1 2.15,1.985 pfet_01v8_hvt
M$4 7 5 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=195000000000P PS=1210000U PD=1390000U
* device instance $5 r0 *1 2.69,1.985 pfet_01v8_hvt
M$5 10 6 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=335000000000P
+ AD=405000000000P PS=2670000U PD=3810000U
* device instance $7 r0 *1 1.77,0.56 nfet_01v8
M$7 8 4 9 11 nfet_01v8 L=150000U W=650000U AS=165350000000P AD=91000000000P
+ PS=1820000U PD=930000U
* device instance $8 r0 *1 2.2,0.56 nfet_01v8
M$8 9 5 8 11 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=104000000000P
+ PS=930000U PD=970000U
* device instance $9 r0 *1 2.67,0.56 nfet_01v8
M$9 10 6 9 11 nfet_01v8 L=150000U W=1300000U AS=195000000000P AD=321750000000P
+ PS=1900000U PD=2940000U
* device instance $11 r0 *1 0.475,0.56 nfet_01v8
M$11 13 2 6 11 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=68250000000P
+ PS=1830000U PD=860000U
* device instance $12 r0 *1 0.835,0.56 nfet_01v8
M$12 8 3 13 11 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=165350000000P
+ PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o211a_2

* cell sky130_fd_sc_hd__a2bb2oi_1
* pin VGND
* pin Y
* pin B2
* pin A1_N
* pin A2_N
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a2bb2oi_1 1 3 4 5 6 7 10 11 13
* net 1 VGND
* net 3 Y
* net 4 B2
* net 5 A1_N
* net 6 A2_N
* net 7 B1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.91,1.985 pfet_01v8_hvt
M$1 9 2 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=340000000000P
+ AD=135000000000P PS=2680000U PD=1270000U
* device instance $2 r0 *1 2.33,1.985 pfet_01v8_hvt
M$2 10 4 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 2.75,1.985 pfet_01v8_hvt
M$3 9 7 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $4 r0 *1 0.47,1.985 pfet_01v8_hvt
M$4 12 5 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=105000000000P PS=2520000U PD=1210000U
* device instance $5 r0 *1 0.83,1.985 pfet_01v8_hvt
M$5 2 6 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 2 5 1 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 0.89,0.56 nfet_01v8
M$7 1 6 2 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=282750000000P
+ PS=920000U PD=1520000U
* device instance $8 r0 *1 1.91,0.56 nfet_01v8
M$8 3 2 1 13 nfet_01v8 L=150000U W=650000U AS=282750000000P AD=87750000000P
+ PS=1520000U PD=920000U
* device instance $9 r0 *1 2.33,0.56 nfet_01v8
M$9 8 4 3 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $10 r0 *1 2.75,0.56 nfet_01v8
M$10 1 7 8 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a2bb2oi_1

* cell sky130_fd_sc_hd__a31oi_2
* pin VGND
* pin Y
* pin A3
* pin A2
* pin A1
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a31oi_2 1 4 5 6 7 8 10 11 12
* net 1 VGND
* net 4 Y
* net 5 A3
* net 6 A2
* net 7 A1
* net 8 B1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 5 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 10 6 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 10 7 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=545000000000P
+ AD=590000000000P PS=3090000U PD=3180000U
* device instance $7 r0 *1 3.63,1.985 pfet_01v8_hvt
M$7 4 8 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=355000000000P
+ AD=435000000000P PS=2710000U PD=3870000U
* device instance $9 r0 *1 2.67,0.56 nfet_01v8
M$9 3 7 4 12 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=214500000000P
+ PS=2770000U PD=1960000U
* device instance $11 r0 *1 3.63,0.56 nfet_01v8
M$11 1 8 4 12 nfet_01v8 L=150000U W=1300000U AS=230750000000P AD=282750000000P
+ PS=2010000U PD=2820000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 1 5 2 12 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $15 r0 *1 1.31,0.56 nfet_01v8
M$15 3 6 2 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__a31oi_2

* cell sky130_fd_sc_hd__a21o_2
* pin VPB
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__a21o_2 1 3 4 5 7 8 9 10
* net 1 VPB
* net 3 B1
* net 4 A1
* net 5 A2
* net 7 VPWR
* net 8 VGND
* net 9 X
* device instance $1 r0 *1 1.855,1.985 pfet_01v8_hvt
M$1 6 3 2 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 2.285,1.985 pfet_01v8_hvt
M$2 7 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=157500000000P PS=1280000U PD=1315000U
* device instance $3 r0 *1 2.75,1.985 pfet_01v8_hvt
M$3 6 5 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=157500000000P
+ AD=260000000000P PS=1315000U PD=2520000U
* device instance $4 r0 *1 0.475,1.985 pfet_01v8_hvt
M$4 9 2 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=405000000000P PS=3810000U PD=3810000U
* device instance $6 r0 *1 0.645,0.56 nfet_01v8
M$6 9 2 8 10 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=201500000000P
+ PS=2760000U PD=1920000U
* device instance $8 r0 *1 1.565,0.56 nfet_01v8
M$8 2 3 8 10 nfet_01v8 L=150000U W=650000U AS=110500000000P AD=162500000000P
+ PS=990000U PD=1150000U
* device instance $9 r0 *1 2.215,0.56 nfet_01v8
M$9 11 4 2 10 nfet_01v8 L=150000U W=650000U AS=162500000000P AD=123500000000P
+ PS=1150000U PD=1030000U
* device instance $10 r0 *1 2.745,0.56 nfet_01v8
M$10 8 5 11 10 nfet_01v8 L=150000U W=650000U AS=123500000000P AD=172250000000P
+ PS=1030000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21o_2

* cell sky130_fd_sc_hd__a211o_1
* pin VPB
* pin B1
* pin C1
* pin A1
* pin A2
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a211o_1 1 2 3 4 5 7 8 9 11
* net 1 VPB
* net 2 B1
* net 3 C1
* net 4 A1
* net 5 A2
* net 7 VPWR
* net 8 X
* net 9 VGND
* device instance $1 r0 *1 1.425,1.985 pfet_01v8_hvt
M$1 7 5 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 1.855,1.985 pfet_01v8_hvt
M$2 10 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $3 r0 *1 2.285,1.985 pfet_01v8_hvt
M$3 12 2 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=155000000000P PS=1280000U PD=1310000U
* device instance $4 r0 *1 2.745,1.985 pfet_01v8_hvt
M$4 6 3 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=155000000000P
+ AD=265000000000P PS=1310000U PD=2530000U
* device instance $5 r0 *1 0.475,1.985 pfet_01v8_hvt
M$5 7 6 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=265000000000P PS=2530000U PD=2530000U
* device instance $6 r0 *1 0.475,0.56 nfet_01v8
M$6 9 6 8 11 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=260000000000P
+ PS=1830000U PD=1450000U
* device instance $7 r0 *1 1.425,0.56 nfet_01v8
M$7 13 5 9 11 nfet_01v8 L=150000U W=650000U AS=260000000000P AD=91000000000P
+ PS=1450000U PD=930000U
* device instance $8 r0 *1 1.855,0.56 nfet_01v8
M$8 6 4 13 11 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=91000000000P
+ PS=930000U PD=930000U
* device instance $9 r0 *1 2.285,0.56 nfet_01v8
M$9 9 2 6 11 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=100750000000P
+ PS=930000U PD=960000U
* device instance $10 r0 *1 2.745,0.56 nfet_01v8
M$10 6 3 9 11 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=172250000000P
+ PS=960000U PD=1830000U
.ENDS sky130_fd_sc_hd__a211o_1

* cell sky130_fd_sc_hd__o221a_1
* pin VGND
* pin X
* pin C1
* pin B1
* pin B2
* pin A2
* pin A1
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o221a_1 1 5 6 7 8 9 10 11 12 15
* net 1 VGND
* net 5 X
* net 6 C1
* net 7 B1
* net 8 B2
* net 9 A2
* net 10 A1
* net 11 VPB
* net 12 VPWR
* device instance $1 r0 *1 0.67,1.985 pfet_01v8_hvt
M$1 12 6 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=340000000000P
+ AD=165000000000P PS=2680000U PD=1330000U
* device instance $2 r0 *1 1.15,1.985 pfet_01v8_hvt
M$2 13 7 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=105000000000P PS=1330000U PD=1210000U
* device instance $3 r0 *1 1.51,1.985 pfet_01v8_hvt
M$3 2 8 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=412500000000P PS=1210000U PD=1825000U
* device instance $4 r0 *1 2.485,1.985 pfet_01v8_hvt
M$4 14 9 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=412500000000P
+ AD=105000000000P PS=1825000U PD=1210000U
* device instance $5 r0 *1 2.845,1.985 pfet_01v8_hvt
M$5 12 10 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=165000000000P PS=1210000U PD=1330000U
* device instance $6 r0 *1 3.325,1.985 pfet_01v8_hvt
M$6 5 2 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=280000000000P PS=1330000U PD=2560000U
* device instance $7 r0 *1 2.485,0.56 nfet_01v8
M$7 4 9 1 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 2.905,0.56 nfet_01v8
M$8 1 10 4 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $9 r0 *1 3.325,0.56 nfet_01v8
M$9 5 2 1 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=182000000000P
+ PS=920000U PD=1860000U
* device instance $10 r0 *1 0.67,0.56 nfet_01v8
M$10 3 6 2 15 nfet_01v8 L=150000U W=650000U AS=201500000000P AD=99125000000P
+ PS=1920000U PD=955000U
* device instance $11 r0 *1 1.125,0.56 nfet_01v8
M$11 4 7 3 15 nfet_01v8 L=150000U W=650000U AS=99125000000P AD=87750000000P
+ PS=955000U PD=920000U
* device instance $12 r0 *1 1.545,0.56 nfet_01v8
M$12 3 8 4 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221a_1

* cell sky130_fd_sc_hd__a21oi_4
* pin VGND
* pin Y
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a21oi_4 1 2 4 5 6 7 8 10
* net 1 VGND
* net 2 Y
* net 4 B1
* net 5 A2
* net 6 A1
* net 7 VPWR
* net 8 VPB
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 2 4 9 8 pfet_01v8_hvt L=150000U W=4000000U AS=680000000000P
+ AD=575000000000P PS=6360000U PD=5150000U
* device instance $5 r0 *1 2.225,1.985 pfet_01v8_hvt
M$5 7 5 9 8 pfet_01v8_hvt L=150000U W=4000000U AS=575000000000P
+ AD=690000000000P PS=5150000U PD=6380000U
* device instance $6 r0 *1 2.665,1.985 pfet_01v8_hvt
M$6 9 6 7 8 pfet_01v8_hvt L=150000U W=4000000U AS=565000000000P
+ AD=560000000000P PS=5130000U PD=5120000U
* device instance $13 r0 *1 0.475,0.56 nfet_01v8
M$13 2 4 1 10 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=377000000000P
+ PS=4620000U PD=3760000U
* device instance $17 r0 *1 2.235,0.56 nfet_01v8
M$17 3 5 1 10 nfet_01v8 L=150000U W=2600000U AS=377000000000P AD=445250000000P
+ PS=3760000U PD=4620000U
* device instance $18 r0 *1 2.665,0.56 nfet_01v8
M$18 2 6 3 10 nfet_01v8 L=150000U W=2600000U AS=364000000000P AD=364000000000P
+ PS=3720000U PD=3720000U
.ENDS sky130_fd_sc_hd__a21oi_4

* cell sky130_fd_sc_hd__a2111oi_0
* pin VGND
* pin D1
* pin Y
* pin A1
* pin C1
* pin B1
* pin A2
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a2111oi_0 1 2 3 4 6 7 8 9 10 14
* net 1 VGND
* net 2 D1
* net 3 Y
* net 4 A1
* net 6 C1
* net 7 B1
* net 8 A2
* net 9 VPB
* net 10 VPWR
* device instance $1 r0 *1 0.77,2.165 pfet_01v8_hvt
M$1 12 2 3 9 pfet_01v8_hvt L=150000U W=640000U AS=188800000000P AD=67200000000P
+ PS=1870000U PD=850000U
* device instance $2 r0 *1 1.13,2.165 pfet_01v8_hvt
M$2 13 6 12 9 pfet_01v8_hvt L=150000U W=640000U AS=67200000000P AD=67200000000P
+ PS=850000U PD=850000U
* device instance $3 r0 *1 1.49,2.165 pfet_01v8_hvt
M$3 11 7 13 9 pfet_01v8_hvt L=150000U W=640000U AS=67200000000P AD=89600000000P
+ PS=850000U PD=920000U
* device instance $4 r0 *1 1.92,2.165 pfet_01v8_hvt
M$4 10 4 11 9 pfet_01v8_hvt L=150000U W=640000U AS=89600000000P
+ AD=121600000000P PS=920000U PD=1020000U
* device instance $5 r0 *1 2.45,2.165 pfet_01v8_hvt
M$5 11 8 10 9 pfet_01v8_hvt L=150000U W=640000U AS=121600000000P
+ AD=195200000000P PS=1020000U PD=1890000U
* device instance $6 r0 *1 0.7,0.445 nfet_01v8
M$6 3 2 1 14 nfet_01v8 L=150000U W=420000U AS=126000000000P AD=58800000000P
+ PS=1440000U PD=700000U
* device instance $7 r0 *1 1.13,0.445 nfet_01v8
M$7 1 6 3 14 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=73500000000P
+ PS=700000U PD=770000U
* device instance $8 r0 *1 1.63,0.445 nfet_01v8
M$8 3 7 1 14 nfet_01v8 L=150000U W=420000U AS=73500000000P AD=58800000000P
+ PS=770000U PD=700000U
* device instance $9 r0 *1 2.06,0.445 nfet_01v8
M$9 5 4 3 14 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=44100000000P
+ PS=700000U PD=630000U
* device instance $10 r0 *1 2.42,0.445 nfet_01v8
M$10 1 8 5 14 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=119700000000P
+ PS=630000U PD=1410000U
.ENDS sky130_fd_sc_hd__a2111oi_0

* cell sky130_fd_sc_hd__o221ai_2
* pin VGND
* pin C1
* pin Y
* pin B1
* pin B2
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o221ai_2 1 3 4 6 7 8 9 10 13 14
* net 1 VGND
* net 3 C1
* net 4 Y
* net 6 B1
* net 7 B2
* net 8 A1
* net 9 A2
* net 10 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 4 3 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=530000000000P PS=3790000U PD=3060000U
* device instance $3 r0 *1 1.835,1.985 pfet_01v8_hvt
M$3 11 6 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=530000000000P
+ AD=310000000000P PS=3060000U PD=2620000U
* device instance $4 r0 *1 2.255,1.985 pfet_01v8_hvt
M$4 4 7 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $7 r0 *1 3.595,1.985 pfet_01v8_hvt
M$7 12 8 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=310000000000P
+ AD=420000000000P PS=2620000U PD=3840000U
* device instance $8 r0 *1 4.015,1.985 pfet_01v8_hvt
M$8 4 9 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $11 r0 *1 1.835,0.56 nfet_01v8
M$11 2 6 5 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=201500000000P
+ PS=2740000U PD=1920000U
* device instance $12 r0 *1 2.255,0.56 nfet_01v8
M$12 5 7 2 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $15 r0 *1 3.595,0.56 nfet_01v8
M$15 1 8 5 14 nfet_01v8 L=150000U W=1300000U AS=201500000000P AD=256750000000P
+ PS=1920000U PD=2740000U
* device instance $16 r0 *1 4.015,0.56 nfet_01v8
M$16 5 9 1 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $19 r0 *1 0.475,0.56 nfet_01v8
M$19 4 3 2 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
.ENDS sky130_fd_sc_hd__o221ai_2

* cell sky130_fd_sc_hd__o211a_4
* pin VGND
* pin X
* pin B1
* pin C1
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o211a_4 1 2 5 6 7 8 11 12 15
* net 1 VGND
* net 2 X
* net 5 B1
* net 6 C1
* net 7 A1
* net 8 A2
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.86,1.985 pfet_01v8_hvt
M$1 2 3 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=560000000000P PS=6370000U PD=5120000U
* device instance $5 r0 *1 2.58,1.985 pfet_01v8_hvt
M$5 3 5 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=335000000000P
+ AD=412500000000P PS=2670000U PD=2825000U
* device instance $6 r0 *1 3.235,1.985 pfet_01v8_hvt
M$6 11 6 3 12 pfet_01v8_hvt L=150000U W=2000000U AS=392500000000P
+ AD=335000000000P PS=2785000U PD=2670000U
* device instance $9 r0 *1 4.675,1.985 pfet_01v8_hvt
M$9 13 7 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=160000000000P
+ AD=140000000000P PS=1320000U PD=1280000U
* device instance $10 r0 *1 5.105,1.985 pfet_01v8_hvt
M$10 3 8 13 12 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $11 r0 *1 5.535,1.985 pfet_01v8_hvt
M$11 14 8 3 12 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $12 r0 *1 5.965,1.985 pfet_01v8_hvt
M$12 11 7 14 12 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=265000000000P PS=1280000U PD=2530000U
* device instance $13 r0 *1 2.71,0.56 nfet_01v8
M$13 9 5 4 15 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=68250000000P
+ PS=1830000U PD=860000U
* device instance $14 r0 *1 3.07,0.56 nfet_01v8
M$14 3 6 9 15 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=144625000000P
+ PS=860000U PD=1095000U
* device instance $15 r0 *1 3.665,0.56 nfet_01v8
M$15 10 6 3 15 nfet_01v8 L=150000U W=650000U AS=144625000000P AD=91000000000P
+ PS=1095000U PD=930000U
* device instance $16 r0 *1 4.095,0.56 nfet_01v8
M$16 4 5 10 15 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=104000000000P
+ PS=930000U PD=970000U
* device instance $17 r0 *1 4.565,0.56 nfet_01v8
M$17 1 7 4 15 nfet_01v8 L=150000U W=1300000U AS=195000000000P AD=299000000000P
+ PS=1900000U PD=2870000U
* device instance $18 r0 *1 5.105,0.56 nfet_01v8
M$18 4 8 1 15 nfet_01v8 L=150000U W=1300000U AS=217750000000P AD=182000000000P
+ PS=1970000U PD=1860000U
* device instance $21 r0 *1 0.47,0.56 nfet_01v8
M$21 2 3 1 15 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=455000000000P
+ PS=4580000U PD=4650000U
.ENDS sky130_fd_sc_hd__o211a_4

* cell sky130_fd_sc_hd__o21ba_2
* pin VPB
* pin B1_N
* pin A1
* pin A2
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__o21ba_2 1 2 3 5 7 8 9 11
* net 1 VPB
* net 2 B1_N
* net 3 A1
* net 5 A2
* net 7 VPWR
* net 8 VGND
* net 9 X
* device instance $1 r0 *1 0.47,1.695 pfet_01v8_hvt
M$1 7 2 4 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=145750000000P
+ PS=1360000U PD=1335000U
* device instance $2 r0 *1 0.955,1.985 pfet_01v8_hvt
M$2 9 6 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=280750000000P
+ AD=530000000000P PS=2605000U PD=3060000U
* device instance $4 r0 *1 2.315,1.985 pfet_01v8_hvt
M$4 6 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=395000000000P
+ AD=165000000000P PS=1790000U PD=1330000U
* device instance $5 r0 *1 2.795,1.985 pfet_01v8_hvt
M$5 12 5 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=105000000000P PS=1330000U PD=1210000U
* device instance $6 r0 *1 3.155,1.985 pfet_01v8_hvt
M$6 7 3 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=280000000000P PS=1210000U PD=2560000U
* device instance $7 r0 *1 2.315,0.56 nfet_01v8
M$7 10 4 6 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=105625000000P
+ PS=1820000U PD=975000U
* device instance $8 r0 *1 2.79,0.56 nfet_01v8
M$8 8 5 10 11 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=87750000000P
+ PS=975000U PD=920000U
* device instance $9 r0 *1 3.21,0.56 nfet_01v8
M$9 10 3 8 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $10 r0 *1 0.47,0.675 nfet_01v8
M$10 4 2 8 11 nfet_01v8 L=150000U W=420000U AS=97000000000P AD=109200000000P
+ PS=975000U PD=1360000U
* device instance $11 r0 *1 0.945,0.56 nfet_01v8
M$11 9 6 8 11 nfet_01v8 L=150000U W=1300000U AS=184750000000P AD=256750000000P
+ PS=1895000U PD=2740000U
.ENDS sky130_fd_sc_hd__o21ba_2

* cell sky130_fd_sc_hd__inv_2
* pin VPB
* pin A
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__inv_2 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 VGND
* net 4 VPWR
* net 5 Y
* device instance $1 r0 *1 0.48,1.985 pfet_01v8_hvt
M$1 5 2 4 1 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $3 r0 *1 0.48,0.56 nfet_01v8
M$3 5 2 3 6 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
.ENDS sky130_fd_sc_hd__inv_2

* cell sky130_fd_sc_hd__o221a_2
* pin VGND
* pin C1
* pin B1
* pin B2
* pin A2
* pin A1
* pin X
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o221a_2 1 2 5 7 8 9 10 11 12 15
* net 1 VGND
* net 2 C1
* net 5 B1
* net 7 B2
* net 8 A2
* net 9 A1
* net 10 X
* net 11 VPB
* net 12 VPWR
* device instance $1 r0 *1 0.63,1.985 pfet_01v8_hvt
M$1 12 2 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=325000000000P
+ AD=165000000000P PS=2650000U PD=1330000U
* device instance $2 r0 *1 1.11,1.985 pfet_01v8_hvt
M$2 13 5 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=112500000000P PS=1330000U PD=1225000U
* device instance $3 r0 *1 1.485,1.985 pfet_01v8_hvt
M$3 3 7 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=112500000000P
+ AD=387500000000P PS=1225000U PD=1775000U
* device instance $4 r0 *1 2.41,1.985 pfet_01v8_hvt
M$4 14 8 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=387500000000P
+ AD=105000000000P PS=1775000U PD=1210000U
* device instance $5 r0 *1 2.77,1.985 pfet_01v8_hvt
M$5 12 9 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=165000000000P PS=1210000U PD=1330000U
* device instance $6 r0 *1 3.25,1.985 pfet_01v8_hvt
M$6 10 3 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=300000000000P
+ AD=395000000000P PS=2600000U PD=3790000U
* device instance $8 r0 *1 2.41,0.56 nfet_01v8
M$8 6 8 1 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $9 r0 *1 2.83,0.56 nfet_01v8
M$9 1 9 6 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $10 r0 *1 3.25,0.56 nfet_01v8
M$10 10 3 1 15 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $12 r0 *1 0.63,0.56 nfet_01v8
M$12 4 2 3 15 nfet_01v8 L=150000U W=650000U AS=237250000000P AD=87750000000P
+ PS=2030000U PD=920000U
* device instance $13 r0 *1 1.05,0.56 nfet_01v8
M$13 6 5 4 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $14 r0 *1 1.47,0.56 nfet_01v8
M$14 4 7 6 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221a_2

* cell sky130_fd_sc_hd__o21bai_4
* pin VGND
* pin B1_N
* pin Y
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o21bai_4 1 2 5 6 7 8 10 11
* net 1 VGND
* net 2 B1_N
* net 5 Y
* net 6 A2
* net 7 A1
* net 8 VPWR
* net 10 VPB
* device instance $1 r0 *1 3.14,1.985 pfet_01v8_hvt
M$1 5 6 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 4.82,1.985 pfet_01v8_hvt
M$5 8 7 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=685000000000P PS=5080000U PD=6370000U
* device instance $9 r0 *1 0.52,1.985 pfet_01v8_hvt
M$9 8 2 3 10 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=135000000000P PS=2560000U PD=1270000U
* device instance $10 r0 *1 0.94,1.985 pfet_01v8_hvt
M$10 5 3 8 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $14 r0 *1 0.52,0.56 nfet_01v8
M$14 3 2 1 11 nfet_01v8 L=150000U W=650000U AS=182000000000P AD=169000000000P
+ PS=1860000U PD=1820000U
* device instance $15 r0 *1 1.46,0.56 nfet_01v8
M$15 5 3 4 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $19 r0 *1 3.14,0.56 nfet_01v8
M$19 1 6 4 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $23 r0 *1 4.82,0.56 nfet_01v8
M$23 1 7 4 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__o21bai_4

* cell sky130_fd_sc_hd__and4_1
* pin VPB
* pin D
* pin C
* pin B
* pin A
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__and4_1 1 3 4 5 6 7 8 9 10
* net 1 VPB
* net 3 D
* net 4 C
* net 5 B
* net 6 A
* net 7 VGND
* net 8 VPWR
* net 9 X
* device instance $1 r0 *1 0.47,2.275 pfet_01v8_hvt
M$1 2 6 8 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=73500000000P
+ PS=1360000U PD=770000U
* device instance $2 r0 *1 0.97,2.275 pfet_01v8_hvt
M$2 8 5 2 1 pfet_01v8_hvt L=150000U W=420000U AS=73500000000P AD=77700000000P
+ PS=770000U PD=790000U
* device instance $3 r0 *1 1.49,2.275 pfet_01v8_hvt
M$3 2 4 8 1 pfet_01v8_hvt L=150000U W=420000U AS=77700000000P AD=58800000000P
+ PS=790000U PD=700000U
* device instance $4 r0 *1 1.92,2.275 pfet_01v8_hvt
M$4 2 3 8 1 pfet_01v8_hvt L=150000U W=420000U AS=312450000000P AD=58800000000P
+ PS=1680000U PD=700000U
* device instance $5 r0 *1 2.75,1.985 pfet_01v8_hvt
M$5 9 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=312450000000P
+ AD=260000000000P PS=1680000U PD=2520000U
* device instance $6 r0 *1 0.47,0.445 nfet_01v8
M$6 13 6 2 10 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=60900000000P
+ PS=1360000U PD=710000U
* device instance $7 r0 *1 0.91,0.445 nfet_01v8
M$7 11 5 13 10 nfet_01v8 L=150000U W=420000U AS=60900000000P AD=79800000000P
+ PS=710000U PD=800000U
* device instance $8 r0 *1 1.44,0.445 nfet_01v8
M$8 12 4 11 10 nfet_01v8 L=150000U W=420000U AS=79800000000P AD=69300000000P
+ PS=800000U PD=750000U
* device instance $9 r0 *1 1.92,0.445 nfet_01v8
M$9 7 3 12 10 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=196275000000P
+ PS=750000U PD=1330000U
* device instance $10 r0 *1 2.75,0.56 nfet_01v8
M$10 9 2 7 10 nfet_01v8 L=150000U W=650000U AS=196275000000P AD=169000000000P
+ PS=1330000U PD=1820000U
.ENDS sky130_fd_sc_hd__and4_1

* cell sky130_fd_sc_hd__nor3b_2
* pin VGND
* pin Y
* pin A
* pin B
* pin C_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor3b_2 1 2 3 4 6 9 10 11
* net 1 VGND
* net 2 Y
* net 3 A
* net 4 B
* net 6 C_N
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 9 3 7 10 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 1.33,1.985 pfet_01v8_hvt
M$3 8 4 7 10 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $5 r0 *1 2.73,1.985 pfet_01v8_hvt
M$5 2 5 8 10 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=415000000000P PS=3830000U PD=3830000U
* device instance $7 r0 *1 4.13,1.695 pfet_01v8_hvt
M$7 9 6 5 10 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=109200000000P PS=1360000U PD=1360000U
* device instance $8 r0 *1 4.13,0.675 nfet_01v8
M$8 1 6 5 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $9 r0 *1 2.73,0.56 nfet_01v8
M$9 2 5 1 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=269750000000P
+ PS=2740000U PD=2780000U
* device instance $11 r0 *1 0.49,0.56 nfet_01v8
M$11 2 3 1 11 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $13 r0 *1 1.33,0.56 nfet_01v8
M$13 2 4 1 11 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nor3b_2

* cell sky130_fd_sc_hd__nand3_2
* pin VGND
* pin Y
* pin A
* pin B
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand3_2 1 3 5 6 7 8 9 10
* net 1 VGND
* net 3 Y
* net 5 A
* net 6 B
* net 7 C
* net 8 VPWR
* net 9 VPB
* device instance $1 r0 *1 2.67,1.985 pfet_01v8_hvt
M$1 3 7 8 9 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=445000000000P PS=3790000U PD=3890000U
* device instance $3 r0 *1 0.47,1.985 pfet_01v8_hvt
M$3 3 5 8 9 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $5 r0 *1 1.31,1.985 pfet_01v8_hvt
M$5 3 6 8 9 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $7 r0 *1 2.67,0.56 nfet_01v8
M$7 4 7 1 10 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=289250000000P
+ PS=2740000U PD=2840000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 3 5 2 10 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $11 r0 *1 1.31,0.56 nfet_01v8
M$11 4 6 2 10 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nand3_2

* cell sky130_fd_sc_hd__and2_1
* pin VPB
* pin A
* pin B
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__and2_1 1 2 3 4 5 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 4 X
* net 5 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.65,2.065 pfet_01v8_hvt
M$1 6 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=117600000000P AD=56700000000P
+ PS=1400000U PD=690000U
* device instance $2 r0 *1 1.07,2.065 pfet_01v8_hvt
M$2 6 3 5 1 pfet_01v8_hvt L=150000U W=420000U AS=166550000000P AD=56700000000P
+ PS=1390000U PD=690000U
* device instance $3 r0 *1 1.61,1.985 pfet_01v8_hvt
M$3 4 6 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=166550000000P
+ AD=475000000000P PS=1390000U PD=2950000U
* device instance $4 r0 *1 0.65,0.585 nfet_01v8
M$4 9 2 6 8 nfet_01v8 L=150000U W=420000U AS=117600000000P AD=56700000000P
+ PS=1400000U PD=690000U
* device instance $5 r0 *1 1.07,0.585 nfet_01v8
M$5 9 3 7 8 nfet_01v8 L=150000U W=420000U AS=111800000000P AD=56700000000P
+ PS=1040000U PD=690000U
* device instance $6 r0 *1 1.61,0.56 nfet_01v8
M$6 4 6 7 8 nfet_01v8 L=150000U W=650000U AS=111800000000P AD=182000000000P
+ PS=1040000U PD=1860000U
.ENDS sky130_fd_sc_hd__and2_1

* cell sky130_fd_sc_hd__a21boi_2
* pin VGND
* pin B1_N
* pin Y
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a21boi_2 1 2 4 5 6 9 10 12
* net 1 VGND
* net 2 B1_N
* net 4 Y
* net 5 A2
* net 6 A1
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 1.42,1.985 pfet_01v8_hvt
M$1 4 3 11 10 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 2.26,1.985 pfet_01v8_hvt
M$3 9 5 11 10 pfet_01v8_hvt L=150000U W=2000000U AS=275000000000P
+ AD=420000000000P PS=2550000U PD=3840000U
* device instance $4 r0 *1 2.68,1.985 pfet_01v8_hvt
M$4 11 6 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=275000000000P
+ AD=280000000000P PS=2550000U PD=2560000U
* device instance $7 r0 *1 0.475,2.1 pfet_01v8_hvt
M$7 3 2 9 10 pfet_01v8_hvt L=150000U W=420000U AS=111300000000P
+ AD=111300000000P PS=1370000U PD=1370000U
* device instance $8 r0 *1 0.68,0.445 nfet_01v8
M$8 1 2 3 12 nfet_01v8 L=150000U W=420000U AS=126000000000P AD=183125000000P
+ PS=1440000U PD=1240000U
* device instance $9 r0 *1 1.42,0.56 nfet_01v8
M$9 4 3 1 12 nfet_01v8 L=150000U W=1300000U AS=270875000000P AD=195000000000P
+ PS=2160000U PD=1900000U
* device instance $11 r0 *1 2.32,0.56 nfet_01v8
M$11 8 5 1 12 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=68250000000P
+ PS=980000U PD=860000U
* device instance $12 r0 *1 2.68,0.56 nfet_01v8
M$12 4 6 8 12 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=91000000000P
+ PS=860000U PD=930000U
* device instance $13 r0 *1 3.11,0.56 nfet_01v8
M$13 7 6 4 12 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=91000000000P
+ PS=930000U PD=930000U
* device instance $14 r0 *1 3.54,0.56 nfet_01v8
M$14 1 5 7 12 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=185250000000P
+ PS=930000U PD=1870000U
.ENDS sky130_fd_sc_hd__a21boi_2

* cell sky130_fd_sc_hd__o211a_1
* pin VGND
* pin X
* pin A1
* pin A2
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o211a_1 1 2 5 6 7 8 10 11 13
* net 1 VGND
* net 2 X
* net 5 A1
* net 6 A2
* net 7 B1
* net 8 C1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.41,1.985 pfet_01v8_hvt
M$1 12 5 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=162500000000P PS=2520000U PD=1325000U
* device instance $2 r0 *1 1.885,1.985 pfet_01v8_hvt
M$2 4 6 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=162500000000P
+ AD=220000000000P PS=1325000U PD=1440000U
* device instance $3 r0 *1 2.475,1.985 pfet_01v8_hvt
M$3 10 7 4 11 pfet_01v8_hvt L=150000U W=1000000U AS=220000000000P
+ AD=175000000000P PS=1440000U PD=1350000U
* device instance $4 r0 *1 2.975,1.985 pfet_01v8_hvt
M$4 4 8 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=175000000000P
+ AD=300000000000P PS=1350000U PD=2600000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 10 4 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $6 r0 *1 1.41,0.56 nfet_01v8
M$6 1 5 3 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=105625000000P
+ PS=1820000U PD=975000U
* device instance $7 r0 *1 1.885,0.56 nfet_01v8
M$7 3 6 1 13 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=143000000000P
+ PS=975000U PD=1090000U
* device instance $8 r0 *1 2.475,0.56 nfet_01v8
M$8 9 7 3 13 nfet_01v8 L=150000U W=650000U AS=143000000000P AD=113750000000P
+ PS=1090000U PD=1000000U
* device instance $9 r0 *1 2.975,0.56 nfet_01v8
M$9 4 8 9 13 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=195000000000P
+ PS=1000000U PD=1900000U
* device instance $10 r0 *1 0.47,0.56 nfet_01v8
M$10 1 4 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__o211a_1

* cell sky130_fd_sc_hd__o21ai_2
* pin VPB
* pin A1
* pin A2
* pin B1
* pin VGND
* pin Y
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o21ai_2 1 2 3 4 7 8 9 10
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 B1
* net 7 VGND
* net 8 Y
* net 9 VPWR
* device instance $1 r0 *1 0.485,1.985 pfet_01v8_hvt
M$1 6 2 9 1 pfet_01v8_hvt L=150000U W=2000000U AS=440000000000P
+ AD=300000000000P PS=3880000U PD=2600000U
* device instance $2 r0 *1 0.915,1.985 pfet_01v8_hvt
M$2 8 3 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=315000000000P PS=2560000U PD=2630000U
* device instance $5 r0 *1 2.315,1.985 pfet_01v8_hvt
M$5 8 4 9 1 pfet_01v8_hvt L=150000U W=2000000U AS=300000000000P
+ AD=405000000000P PS=2600000U PD=3810000U
* device instance $7 r0 *1 0.485,0.56 nfet_01v8
M$7 7 2 5 10 nfet_01v8 L=150000U W=1300000U AS=299000000000P AD=182000000000P
+ PS=2870000U PD=1860000U
* device instance $8 r0 *1 0.915,0.56 nfet_01v8
M$8 5 3 7 10 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=217750000000P
+ PS=1860000U PD=1970000U
* device instance $11 r0 *1 2.315,0.56 nfet_01v8
M$11 8 4 5 10 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=263250000000P
+ PS=1860000U PD=2760000U
.ENDS sky130_fd_sc_hd__o21ai_2

* cell sky130_fd_sc_hd__or2_0
* pin VPB
* pin B
* pin A
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__or2_0 1 2 3 4 6 7 8
* net 1 VPB
* net 2 B
* net 3 A
* net 4 X
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.675,1.985 pfet_01v8_hvt
M$1 9 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 1.035,1.985 pfet_01v8_hvt
M$2 7 3 9 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=98950000000P
+ PS=630000U PD=975000U
* device instance $3 r0 *1 1.52,2.095 pfet_01v8_hvt
M$3 4 5 7 1 pfet_01v8_hvt L=150000U W=640000U AS=98950000000P AD=217600000000P
+ PS=975000U PD=1960000U
* device instance $4 r0 *1 0.615,0.675 nfet_01v8
M$4 5 2 6 8 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $5 r0 *1 1.035,0.675 nfet_01v8
M$5 6 3 5 8 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=70350000000P
+ PS=690000U PD=755000U
* device instance $6 r0 *1 1.52,0.675 nfet_01v8
M$6 4 5 6 8 nfet_01v8 L=150000U W=420000U AS=70350000000P AD=109200000000P
+ PS=755000U PD=1360000U
.ENDS sky130_fd_sc_hd__or2_0

* cell sky130_fd_sc_hd__o2bb2ai_1
* pin VPB
* pin A1_N
* pin A2_N
* pin B2
* pin B1
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o2bb2ai_1 1 2 3 4 5 6 8 10 11
* net 1 VPB
* net 2 A1_N
* net 3 A2_N
* net 4 B2
* net 5 B1
* net 6 VPWR
* net 8 Y
* net 10 VGND
* device instance $1 r0 *1 0.485,1.985 pfet_01v8_hvt
M$1 7 2 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=275000000000P
+ AD=135000000000P PS=2550000U PD=1270000U
* device instance $2 r0 *1 0.905,1.985 pfet_01v8_hvt
M$2 6 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=420000000000P PS=1270000U PD=1840000U
* device instance $3 r0 *1 1.895,1.985 pfet_01v8_hvt
M$3 8 7 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=420000000000P
+ AD=135000000000P PS=1840000U PD=1270000U
* device instance $4 r0 *1 2.315,1.985 pfet_01v8_hvt
M$4 12 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $5 r0 *1 2.735,1.985 pfet_01v8_hvt
M$5 6 5 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=275000000000P PS=1270000U PD=2550000U
* device instance $6 r0 *1 1.895,0.56 nfet_01v8
M$6 9 7 8 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 2.315,0.56 nfet_01v8
M$7 10 4 9 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $8 r0 *1 2.735,0.56 nfet_01v8
M$8 9 5 10 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $9 r0 *1 0.485,0.56 nfet_01v8
M$9 13 2 10 11 nfet_01v8 L=150000U W=650000U AS=178750000000P AD=68250000000P
+ PS=1850000U PD=860000U
* device instance $10 r0 *1 0.845,0.56 nfet_01v8
M$10 7 3 13 11 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=240500000000P
+ PS=860000U PD=2040000U
.ENDS sky130_fd_sc_hd__o2bb2ai_1

* cell sky130_fd_sc_hd__a22oi_2
* pin VGND
* pin B2
* pin B1
* pin Y
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a22oi_2 1 3 4 5 7 8 10 11 12
* net 1 VGND
* net 3 B2
* net 4 B1
* net 5 Y
* net 7 A1
* net 8 A2
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.67,1.985 pfet_01v8_hvt
M$1 10 7 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 3.51,1.985 pfet_01v8_hvt
M$3 10 8 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 9 3 5 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $7 r0 *1 1.31,1.985 pfet_01v8_hvt
M$7 9 4 5 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $9 r0 *1 2.67,0.56 nfet_01v8
M$9 5 7 6 12 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $11 r0 *1 3.51,0.56 nfet_01v8
M$11 1 8 6 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 1 3 2 12 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $15 r0 *1 1.31,0.56 nfet_01v8
M$15 5 4 2 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__a22oi_2

* cell sky130_fd_sc_hd__clkinvlp_4
* pin VPB
* pin A
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__clkinvlp_4 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 VPWR
* net 4 VGND
* net 5 Y
* device instance $1 r0 *1 0.525,1.985 pfet_01v8_hvt
M$1 5 2 3 1 pfet_01v8_hvt L=250000U W=4000000U AS=685000000000P
+ AD=685000000000P PS=6370000U PD=6370000U
* device instance $5 r0 *1 0.475,0.51 nfet_01v8
M$5 8 2 4 6 nfet_01v8 L=150000U W=550000U AS=145750000000P AD=57750000000P
+ PS=1630000U PD=760000U
* device instance $6 r0 *1 0.835,0.51 nfet_01v8
M$6 5 2 8 6 nfet_01v8 L=150000U W=550000U AS=57750000000P AD=77000000000P
+ PS=760000U PD=830000U
* device instance $7 r0 *1 1.265,0.51 nfet_01v8
M$7 7 2 5 6 nfet_01v8 L=150000U W=550000U AS=77000000000P AD=57750000000P
+ PS=830000U PD=760000U
* device instance $8 r0 *1 1.625,0.51 nfet_01v8
M$8 4 2 7 6 nfet_01v8 L=150000U W=550000U AS=57750000000P AD=145750000000P
+ PS=760000U PD=1630000U
.ENDS sky130_fd_sc_hd__clkinvlp_4

* cell sky130_fd_sc_hd__a2bb2oi_2
* pin VGND
* pin Y
* pin B1
* pin B2
* pin A1_N
* pin A2_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a2bb2oi_2 1 3 5 6 7 8 10 11 13
* net 1 VGND
* net 3 Y
* net 5 B1
* net 6 B2
* net 7 A1_N
* net 8 A2_N
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 3.645,1.985 pfet_01v8_hvt
M$1 10 7 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 4.485,1.985 pfet_01v8_hvt
M$3 4 8 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $5 r0 *1 0.605,1.985 pfet_01v8_hvt
M$5 10 5 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $6 r0 *1 1.025,1.985 pfet_01v8_hvt
M$6 12 6 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $9 r0 *1 2.285,1.985 pfet_01v8_hvt
M$9 3 4 12 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $11 r0 *1 0.605,0.56 nfet_01v8
M$11 2 5 1 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $12 r0 *1 1.025,0.56 nfet_01v8
M$12 3 6 2 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $15 r0 *1 2.285,0.56 nfet_01v8
M$15 3 4 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=344500000000P
+ PS=1840000U PD=2360000U
* device instance $17 r0 *1 3.645,0.56 nfet_01v8
M$17 4 7 1 13 nfet_01v8 L=150000U W=1300000U AS=344500000000P AD=175500000000P
+ PS=2360000U PD=1840000U
* device instance $19 r0 *1 4.485,0.56 nfet_01v8
M$19 4 8 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
.ENDS sky130_fd_sc_hd__a2bb2oi_2

* cell sky130_fd_sc_hd__and4_2
* pin VGND
* pin B
* pin C
* pin X
* pin A
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__and4_2 1 3 4 5 6 7 11 12 13
* net 1 VGND
* net 3 B
* net 4 C
* net 5 X
* net 6 A
* net 7 D
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.47,2.275 pfet_01v8_hvt
M$1 2 6 11 12 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=74550000000P PS=1360000U PD=775000U
* device instance $2 r0 *1 0.975,2.275 pfet_01v8_hvt
M$2 11 3 2 12 pfet_01v8_hvt L=150000U W=420000U AS=74550000000P AD=77700000000P
+ PS=775000U PD=790000U
* device instance $3 r0 *1 1.495,2.275 pfet_01v8_hvt
M$3 2 4 11 12 pfet_01v8_hvt L=150000U W=420000U AS=77700000000P AD=58800000000P
+ PS=790000U PD=700000U
* device instance $4 r0 *1 1.925,2.275 pfet_01v8_hvt
M$4 2 7 11 12 pfet_01v8_hvt L=150000U W=420000U AS=279950000000P
+ AD=58800000000P PS=1615000U PD=700000U
* device instance $5 r0 *1 2.69,1.985 pfet_01v8_hvt
M$5 5 2 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=444950000000P
+ AD=465000000000P PS=2945000U PD=3930000U
* device instance $7 r0 *1 0.47,0.445 nfet_01v8
M$7 8 6 2 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=61950000000P
+ PS=1360000U PD=715000U
* device instance $8 r0 *1 0.915,0.445 nfet_01v8
M$8 9 3 8 13 nfet_01v8 L=150000U W=420000U AS=61950000000P AD=79800000000P
+ PS=715000U PD=800000U
* device instance $9 r0 *1 1.445,0.445 nfet_01v8
M$9 10 4 9 13 nfet_01v8 L=150000U W=420000U AS=79800000000P AD=69300000000P
+ PS=800000U PD=750000U
* device instance $10 r0 *1 1.925,0.445 nfet_01v8
M$10 1 7 10 13 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=175150000000P
+ PS=750000U PD=1265000U
* device instance $11 r0 *1 2.69,0.56 nfet_01v8
M$11 5 2 1 13 nfet_01v8 L=150000U W=1300000U AS=282400000000P AD=302250000000P
+ PS=2245000U PD=2880000U
.ENDS sky130_fd_sc_hd__and4_2

* cell sky130_fd_sc_hd__o32ai_4
* pin VGND
* pin B1
* pin A2
* pin A1
* pin Y
* pin A3
* pin B2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o32ai_4 1 2 3 4 6 7 8 12 13 14
* net 1 VGND
* net 2 B1
* net 3 A2
* net 4 A1
* net 6 Y
* net 7 A3
* net 8 B2
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 8.245,1.985 pfet_01v8_hvt
M$1 11 4 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=712500000000P
+ AD=712500000000P PS=6425000U PD=6425000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 6 8 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=547500000000P PS=6330000U PD=5095000U
* device instance $9 r0 *1 2.165,1.985 pfet_01v8_hvt
M$9 12 2 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=547500000000P
+ AD=665000000000P PS=5095000U PD=6330000U
* device instance $13 r0 *1 4.365,1.985 pfet_01v8_hvt
M$13 6 7 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $17 r0 *1 6.045,1.985 pfet_01v8_hvt
M$17 11 3 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 0.47,0.56 nfet_01v8
M$21 6 8 5 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=355875000000P
+ PS=4580000U PD=3695000U
* device instance $25 r0 *1 2.165,0.56 nfet_01v8
M$25 6 2 5 14 nfet_01v8 L=150000U W=2600000U AS=355875000000P AD=351000000000P
+ PS=3695000U PD=3680000U
* device instance $29 r0 *1 3.845,0.56 nfet_01v8
M$29 1 7 5 14 nfet_01v8 L=150000U W=2600000U AS=403000000000P AD=520000000000P
+ PS=3840000U PD=4200000U
* device instance $33 r0 *1 6.045,0.56 nfet_01v8
M$33 1 3 5 14 nfet_01v8 L=150000U W=2600000U AS=468000000000P AD=520000000000P
+ PS=4040000U PD=4200000U
* device instance $37 r0 *1 8.245,0.56 nfet_01v8
M$37 1 4 5 14 nfet_01v8 L=150000U W=2600000U AS=550875000000P AD=463125000000P
+ PS=4295000U PD=4675000U
.ENDS sky130_fd_sc_hd__o32ai_4

* cell sky130_fd_sc_hd__o31ai_1
* pin VPB
* pin A1
* pin A2
* pin A3
* pin B1
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__o31ai_1 1 2 3 4 5 6 7 9 10
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 A3
* net 5 B1
* net 6 VPWR
* net 7 VGND
* net 9 Y
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 12 2 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 11 3 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 9 4 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=392500000000P PS=1270000U PD=1785000U
* device instance $4 r0 *1 2.245,1.985 pfet_01v8_hvt
M$4 6 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=392500000000P
+ AD=300000000000P PS=1785000U PD=2600000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 8 2 7 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $6 r0 *1 0.89,0.56 nfet_01v8
M$6 7 3 8 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $7 r0 *1 1.31,0.56 nfet_01v8
M$7 8 4 7 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=198250000000P
+ PS=920000U PD=1260000U
* device instance $8 r0 *1 2.07,0.56 nfet_01v8
M$8 9 5 8 10 nfet_01v8 L=150000U W=650000U AS=198250000000P AD=221000000000P
+ PS=1260000U PD=1980000U
.ENDS sky130_fd_sc_hd__o31ai_1

* cell sky130_fd_sc_hd__a221o_1
* pin VGND
* pin B1
* pin A1
* pin X
* pin C1
* pin B2
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a221o_1 1 3 4 5 8 9 10 13 14 15
* net 1 VGND
* net 3 B1
* net 4 A1
* net 5 X
* net 8 C1
* net 9 B2
* net 10 A2
* net 13 VPWR
* net 14 VPB
* device instance $1 r0 *1 2.25,1.985 pfet_01v8_hvt
M$1 12 4 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=165000000000P PS=2520000U PD=1330000U
* device instance $2 r0 *1 2.73,1.985 pfet_01v8_hvt
M$2 13 10 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=157500000000P PS=1330000U PD=1315000U
* device instance $3 r0 *1 3.195,1.985 pfet_01v8_hvt
M$3 5 2 13 14 pfet_01v8_hvt L=150000U W=1000000U AS=157500000000P
+ AD=260000000000P PS=1315000U PD=2520000U
* device instance $4 r0 *1 0.47,1.985 pfet_01v8_hvt
M$4 11 8 2 14 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $5 r0 *1 0.89,1.985 pfet_01v8_hvt
M$5 12 9 11 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $6 r0 *1 1.31,1.985 pfet_01v8_hvt
M$6 11 3 12 14 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $7 r0 *1 2.25,0.56 nfet_01v8
M$7 7 4 2 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $8 r0 *1 2.73,0.56 nfet_01v8
M$8 1 10 7 15 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=102375000000P
+ PS=980000U PD=965000U
* device instance $9 r0 *1 3.195,0.56 nfet_01v8
M$9 5 2 1 15 nfet_01v8 L=150000U W=650000U AS=102375000000P AD=169000000000P
+ PS=965000U PD=1820000U
* device instance $10 r0 *1 0.47,0.56 nfet_01v8
M$10 1 8 2 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $11 r0 *1 0.95,0.56 nfet_01v8
M$11 6 9 1 15 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=68250000000P
+ PS=980000U PD=860000U
* device instance $12 r0 *1 1.31,0.56 nfet_01v8
M$12 2 3 6 15 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=169000000000P
+ PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__a221o_1

* cell sky130_fd_sc_hd__o22ai_4
* pin VGND
* pin B1
* pin B2
* pin A1
* pin A2
* pin Y
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o22ai_4 1 2 3 5 6 7 9 10 12
* net 1 VGND
* net 2 B1
* net 3 B2
* net 5 A1
* net 6 A2
* net 7 Y
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.5,1.985 pfet_01v8_hvt
M$1 8 5 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=695000000000P
+ AD=565000000000P PS=6390000U PD=5130000U
* device instance $4 r0 *1 1.76,1.985 pfet_01v8_hvt
M$4 7 6 8 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $9 r0 *1 3.91,1.985 pfet_01v8_hvt
M$9 11 2 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=565000000000P
+ AD=665000000000P PS=5130000U PD=6330000U
* device instance $12 r0 *1 5.17,1.985 pfet_01v8_hvt
M$12 7 3 11 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $17 r0 *1 0.5,0.56 nfet_01v8
M$17 1 5 4 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=367250000000P
+ PS=4580000U PD=3730000U
* device instance $20 r0 *1 1.76,0.56 nfet_01v8
M$20 4 6 1 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $25 r0 *1 3.91,0.56 nfet_01v8
M$25 7 2 4 12 nfet_01v8 L=150000U W=2600000U AS=367250000000P AD=432250000000P
+ PS=3730000U PD=4580000U
* device instance $28 r0 *1 5.17,0.56 nfet_01v8
M$28 4 3 7 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
.ENDS sky130_fd_sc_hd__o22ai_4

* cell sky130_fd_sc_hd__nor4_4
* pin VGND
* pin C
* pin Y
* pin A
* pin B
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor4_4 1 2 3 4 6 7 8 11 12
* net 1 VGND
* net 2 C
* net 3 Y
* net 4 A
* net 6 B
* net 7 D
* net 8 VPWR
* net 11 VPB
* device instance $1 r0 *1 4.37,1.985 pfet_01v8_hvt
M$1 9 2 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 6.05,1.985 pfet_01v8_hvt
M$5 3 7 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $9 r0 *1 0.49,1.985 pfet_01v8_hvt
M$9 8 4 5 11 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $13 r0 *1 2.17,1.985 pfet_01v8_hvt
M$13 9 6 5 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $17 r0 *1 0.49,0.56 nfet_01v8
M$17 3 4 1 12 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $21 r0 *1 2.17,0.56 nfet_01v8
M$21 3 6 1 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=520000000000P
+ PS=3680000U PD=4200000U
* device instance $25 r0 *1 4.37,0.56 nfet_01v8
M$25 3 2 1 12 nfet_01v8 L=150000U W=2600000U AS=520000000000P AD=351000000000P
+ PS=4200000U PD=3680000U
* device instance $29 r0 *1 6.05,0.56 nfet_01v8
M$29 3 7 1 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nor4_4

* cell sky130_fd_sc_hd__nor2b_2
* pin VPB
* pin B_N
* pin A
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__nor2b_2 1 2 4 5 7 8 9
* net 1 VPB
* net 2 B_N
* net 4 A
* net 5 VGND
* net 7 VPWR
* net 8 Y
* device instance $1 r0 *1 2.69,2.275 pfet_01v8_hvt
M$1 7 2 3 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $2 r0 *1 0.49,1.985 pfet_01v8_hvt
M$2 7 4 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $4 r0 *1 1.33,1.985 pfet_01v8_hvt
M$4 8 3 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $6 r0 *1 2.69,0.675 nfet_01v8
M$6 5 2 3 9 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $7 r0 *1 0.49,0.56 nfet_01v8
M$7 8 4 5 9 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=175500000000P
+ PS=2770000U PD=1840000U
* device instance $9 r0 *1 1.33,0.56 nfet_01v8
M$9 8 3 5 9 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nor2b_2

* cell sky130_fd_sc_hd__nor4_2
* pin VGND
* pin Y
* pin A
* pin B
* pin C
* pin D
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor4_2 1 2 3 4 5 6 8 11 12
* net 1 VGND
* net 2 Y
* net 3 A
* net 4 B
* net 5 C
* net 6 D
* net 8 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.73,1.985 pfet_01v8_hvt
M$1 9 5 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 3.57,1.985 pfet_01v8_hvt
M$3 2 6 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 0.49,1.985 pfet_01v8_hvt
M$5 8 3 7 11 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $7 r0 *1 1.33,1.985 pfet_01v8_hvt
M$7 9 4 7 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $9 r0 *1 2.73,0.56 nfet_01v8
M$9 2 5 1 12 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $11 r0 *1 3.57,0.56 nfet_01v8
M$11 2 6 1 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $13 r0 *1 0.49,0.56 nfet_01v8
M$13 2 3 1 12 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $15 r0 *1 1.33,0.56 nfet_01v8
M$15 2 4 1 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
.ENDS sky130_fd_sc_hd__nor4_2

* cell sky130_fd_sc_hd__or3_1
* pin VPB
* pin A
* pin B
* pin C
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__or3_1 1 2 3 4 5 6 7 9
* net 1 VPB
* net 2 A
* net 3 B
* net 4 C
* net 5 X
* net 6 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.48,1.695 pfet_01v8_hvt
M$1 11 4 8 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 0.84,1.695 pfet_01v8_hvt
M$2 10 3 11 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $3 r0 *1 1.32,1.695 pfet_01v8_hvt
M$3 6 2 10 1 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P AD=148250000000P
+ PS=750000U PD=1340000U
* device instance $4 r0 *1 1.81,1.985 pfet_01v8_hvt
M$4 5 8 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=148250000000P
+ AD=280000000000P PS=1340000U PD=2560000U
* device instance $5 r0 *1 0.48,0.475 nfet_01v8
M$5 7 4 8 9 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $6 r0 *1 0.9,0.475 nfet_01v8
M$6 8 3 7 9 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $7 r0 *1 1.32,0.475 nfet_01v8
M$7 8 2 7 9 nfet_01v8 L=150000U W=420000U AS=101875000000P AD=56700000000P
+ PS=990000U PD=690000U
* device instance $8 r0 *1 1.81,0.56 nfet_01v8
M$8 5 8 7 9 nfet_01v8 L=150000U W=650000U AS=101875000000P AD=182000000000P
+ PS=990000U PD=1860000U
.ENDS sky130_fd_sc_hd__or3_1

* cell sky130_fd_sc_hd__nand3_1
* pin VPB
* pin A
* pin B
* pin C
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__nand3_1 1 2 3 4 5 6 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 4 C
* net 5 Y
* net 6 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 5 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 6 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $3 r0 *1 1.37,1.985 pfet_01v8_hvt
M$3 5 2 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=260000000000P PS=1330000U PD=2520000U
* device instance $4 r0 *1 0.47,0.56 nfet_01v8
M$4 10 4 7 8 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $5 r0 *1 0.89,0.56 nfet_01v8
M$5 9 3 10 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $6 r0 *1 1.37,0.56 nfet_01v8
M$6 5 2 9 8 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=169000000000P
+ PS=980000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand3_1

* cell sky130_fd_sc_hd__nor4_1
* pin VPB
* pin D
* pin B
* pin A
* pin C
* pin VGND
* pin Y
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor4_1 1 2 3 4 5 6 7 8 9
* net 1 VPB
* net 2 D
* net 3 B
* net 4 A
* net 5 C
* net 6 VGND
* net 7 Y
* net 8 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 11 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=130000000000P PS=2520000U PD=1260000U
* device instance $2 r0 *1 0.88,1.985 pfet_01v8_hvt
M$2 10 5 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=130000000000P
+ AD=190000000000P PS=1260000U PD=1380000U
* device instance $3 r0 *1 1.41,1.985 pfet_01v8_hvt
M$3 12 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=190000000000P
+ AD=135000000000P PS=1380000U PD=1270000U
* device instance $4 r0 *1 1.83,1.985 pfet_01v8_hvt
M$4 8 4 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 7 2 6 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=118625000000P
+ PS=1820000U PD=1015000U
* device instance $6 r0 *1 0.985,0.56 nfet_01v8
M$6 6 5 7 9 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=89375000000P
+ PS=1015000U PD=925000U
* device instance $7 r0 *1 1.41,0.56 nfet_01v8
M$7 7 3 6 9 nfet_01v8 L=150000U W=650000U AS=89375000000P AD=87750000000P
+ PS=925000U PD=920000U
* device instance $8 r0 *1 1.83,0.56 nfet_01v8
M$8 6 4 7 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor4_1

* cell sky130_fd_sc_hd__ha_1
* pin VGND
* pin SUM
* pin COUT
* pin A
* pin B
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__ha_1 1 2 5 8 9 10 11 13
* net 1 VGND
* net 2 SUM
* net 5 COUT
* net 8 A
* net 9 B
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 3 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=236050000000P PS=2520000U PD=1765000U
* device instance $2 r0 *1 1.385,2.275 pfet_01v8_hvt
M$2 3 7 10 11 pfet_01v8_hvt L=150000U W=420000U AS=236050000000P
+ AD=56700000000P PS=1765000U PD=690000U
* device instance $3 r0 *1 1.805,2.275 pfet_01v8_hvt
M$3 12 9 3 11 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P AD=84000000000P
+ PS=690000U PD=820000U
* device instance $4 r0 *1 2.355,2.275 pfet_01v8_hvt
M$4 10 8 12 11 pfet_01v8_hvt L=150000U W=420000U AS=84000000000P
+ AD=149100000000P PS=820000U PD=1130000U
* device instance $5 r0 *1 3.215,2.275 pfet_01v8_hvt
M$5 7 9 10 11 pfet_01v8_hvt L=150000U W=420000U AS=149100000000P
+ AD=60900000000P PS=1130000U PD=710000U
* device instance $6 r0 *1 3.655,2.275 pfet_01v8_hvt
M$6 7 8 10 11 pfet_01v8_hvt L=150000U W=420000U AS=140750000000P
+ AD=60900000000P PS=1325000U PD=710000U
* device instance $7 r0 *1 4.13,1.985 pfet_01v8_hvt
M$7 5 7 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=140750000000P
+ AD=260000000000P PS=1325000U PD=2520000U
* device instance $8 r0 *1 3.295,0.445 nfet_01v8
M$8 6 9 7 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $9 r0 *1 3.655,0.445 nfet_01v8
M$9 1 8 6 13 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=97000000000P
+ PS=630000U PD=975000U
* device instance $10 r0 *1 4.13,0.56 nfet_01v8
M$10 5 7 1 13 nfet_01v8 L=150000U W=650000U AS=97000000000P AD=169000000000P
+ PS=975000U PD=1820000U
* device instance $11 r0 *1 1.41,0.445 nfet_01v8
M$11 4 7 3 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $12 r0 *1 1.83,0.445 nfet_01v8
M$12 1 9 4 13 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $13 r0 *1 2.25,0.445 nfet_01v8
M$13 4 8 1 13 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $14 r0 *1 0.47,0.56 nfet_01v8
M$14 1 3 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__ha_1

* cell sky130_fd_sc_hd__fa_1
* pin VGND
* pin COUT
* pin SUM
* pin A
* pin CIN
* pin B
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__fa_1 1 2 7 11 12 13 16 17 21
* net 1 VGND
* net 2 COUT
* net 7 SUM
* net 11 A
* net 12 CIN
* net 13 B
* net 16 VPWR
* net 17 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 16 3 2 17 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=147850000000P PS=2520000U PD=1345000U
* device instance $2 r0 *1 0.965,2.275 pfet_01v8_hvt
M$2 18 11 16 17 pfet_01v8_hvt L=150000U W=420000U AS=147850000000P
+ AD=63000000000P PS=1345000U PD=720000U
* device instance $3 r0 *1 1.415,2.275 pfet_01v8_hvt
M$3 3 13 18 17 pfet_01v8_hvt L=150000U W=420000U AS=63000000000P
+ AD=56700000000P PS=720000U PD=690000U
* device instance $4 r0 *1 1.835,2.275 pfet_01v8_hvt
M$4 14 12 3 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
* device instance $5 r0 *1 2.255,2.275 pfet_01v8_hvt
M$5 16 11 14 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
* device instance $6 r0 *1 2.675,2.275 pfet_01v8_hvt
M$6 14 13 16 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=109200000000P PS=690000U PD=1360000U
* device instance $7 r0 *1 3.615,2.275 pfet_01v8_hvt
M$7 15 13 16 17 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
* device instance $8 r0 *1 4.035,2.275 pfet_01v8_hvt
M$8 16 12 15 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
* device instance $9 r0 *1 4.455,2.275 pfet_01v8_hvt
M$9 15 11 16 17 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P
+ AD=61950000000P PS=690000U PD=715000U
* device instance $10 r0 *1 4.9,2.275 pfet_01v8_hvt
M$10 6 3 15 17 pfet_01v8_hvt L=150000U W=420000U AS=61950000000P
+ AD=69300000000P PS=715000U PD=750000U
* device instance $11 r0 *1 5.38,2.275 pfet_01v8_hvt
M$11 19 12 6 17 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P
+ AD=44100000000P PS=750000U PD=630000U
* device instance $12 r0 *1 5.74,2.275 pfet_01v8_hvt
M$12 20 13 19 17 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P
+ AD=69300000000P PS=630000U PD=750000U
* device instance $13 r0 *1 6.22,2.275 pfet_01v8_hvt
M$13 20 11 16 17 pfet_01v8_hvt L=150000U W=420000U AS=147850000000P
+ AD=69300000000P PS=1345000U PD=750000U
* device instance $14 r0 *1 6.715,1.985 pfet_01v8_hvt
M$14 7 6 16 17 pfet_01v8_hvt L=150000U W=1000000U AS=147850000000P
+ AD=260000000000P PS=1345000U PD=2520000U
* device instance $15 r0 *1 0.965,0.445 nfet_01v8
M$15 8 11 1 21 nfet_01v8 L=150000U W=420000U AS=102350000000P AD=63000000000P
+ PS=995000U PD=720000U
* device instance $16 r0 *1 1.415,0.445 nfet_01v8
M$16 3 13 8 21 nfet_01v8 L=150000U W=420000U AS=63000000000P AD=56700000000P
+ PS=720000U PD=690000U
* device instance $17 r0 *1 1.835,0.445 nfet_01v8
M$17 4 12 3 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $18 r0 *1 2.255,0.445 nfet_01v8
M$18 1 11 4 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $19 r0 *1 2.675,0.445 nfet_01v8
M$19 4 13 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=109200000000P
+ PS=690000U PD=1360000U
* device instance $20 r0 *1 0.47,0.56 nfet_01v8
M$20 1 3 2 21 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=102350000000P
+ PS=1820000U PD=995000U
* device instance $21 r0 *1 3.615,0.445 nfet_01v8
M$21 5 13 1 21 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $22 r0 *1 4.035,0.445 nfet_01v8
M$22 1 12 5 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=56700000000P
+ PS=690000U PD=690000U
* device instance $23 r0 *1 4.455,0.445 nfet_01v8
M$23 5 11 1 21 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=61950000000P
+ PS=690000U PD=715000U
* device instance $24 r0 *1 4.9,0.445 nfet_01v8
M$24 6 3 5 21 nfet_01v8 L=150000U W=420000U AS=61950000000P AD=69300000000P
+ PS=715000U PD=750000U
* device instance $25 r0 *1 5.38,0.445 nfet_01v8
M$25 10 12 6 21 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=44100000000P
+ PS=750000U PD=630000U
* device instance $26 r0 *1 5.74,0.445 nfet_01v8
M$26 9 13 10 21 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=69300000000P
+ PS=630000U PD=750000U
* device instance $27 r0 *1 6.22,0.445 nfet_01v8
M$27 1 11 9 21 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=102350000000P
+ PS=750000U PD=995000U
* device instance $28 r0 *1 6.715,0.56 nfet_01v8
M$28 7 6 1 21 nfet_01v8 L=150000U W=650000U AS=102350000000P AD=169000000000P
+ PS=995000U PD=1820000U
.ENDS sky130_fd_sc_hd__fa_1

* cell sky130_fd_sc_hd__a311o_1
* pin VPB
* pin C1
* pin B1
* pin A1
* pin A2
* pin A3
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a311o_1 1 2 3 4 5 6 7 8 10 12
* net 1 VPB
* net 2 C1
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 A3
* net 7 X
* net 8 VGND
* net 10 VPWR
* device instance $1 r0 *1 0.495,1.985 pfet_01v8_hvt
M$1 10 11 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=285000000000P
+ AD=142500000000P PS=2570000U PD=1285000U
* device instance $2 r0 *1 0.93,1.985 pfet_01v8_hvt
M$2 9 6 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=142500000000P
+ AD=165000000000P PS=1285000U PD=1330000U
* device instance $3 r0 *1 1.41,1.985 pfet_01v8_hvt
M$3 10 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=305000000000P PS=1330000U PD=1610000U
* device instance $4 r0 *1 2.17,1.985 pfet_01v8_hvt
M$4 9 4 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=305000000000P
+ AD=162500000000P PS=1610000U PD=1325000U
* device instance $5 r0 *1 2.645,1.985 pfet_01v8_hvt
M$5 13 3 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=162500000000P
+ AD=207500000000P PS=1325000U PD=1415000U
* device instance $6 r0 *1 3.21,1.985 pfet_01v8_hvt
M$6 11 2 13 1 pfet_01v8_hvt L=150000U W=1000000U AS=207500000000P
+ AD=260000000000P PS=1415000U PD=2520000U
* device instance $7 r0 *1 0.47,0.56 nfet_01v8
M$7 8 11 7 12 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=112125000000P
+ PS=1820000U PD=995000U
* device instance $8 r0 *1 0.965,0.56 nfet_01v8
M$8 15 6 8 12 nfet_01v8 L=150000U W=650000U AS=112125000000P AD=125125000000P
+ PS=995000U PD=1035000U
* device instance $9 r0 *1 1.5,0.56 nfet_01v8
M$9 14 5 15 12 nfet_01v8 L=150000U W=650000U AS=125125000000P AD=169000000000P
+ PS=1035000U PD=1170000U
* device instance $10 r0 *1 2.17,0.56 nfet_01v8
M$10 11 4 14 12 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=105625000000P
+ PS=1170000U PD=975000U
* device instance $11 r0 *1 2.645,0.56 nfet_01v8
M$11 8 3 11 12 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=134875000000P
+ PS=975000U PD=1065000U
* device instance $12 r0 *1 3.21,0.56 nfet_01v8
M$12 11 2 8 12 nfet_01v8 L=150000U W=650000U AS=134875000000P AD=169000000000P
+ PS=1065000U PD=1820000U
.ENDS sky130_fd_sc_hd__a311o_1

* cell sky130_fd_sc_hd__a22oi_4
* pin VGND
* pin B1
* pin A1
* pin B2
* pin Y
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a22oi_4 1 2 3 5 6 8 10 11 12
* net 1 VGND
* net 2 B1
* net 3 A1
* net 5 B2
* net 6 Y
* net 8 A2
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 6 5 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 6 2 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=800000000000P PS=5080000U PD=5600000U
* device instance $9 r0 *1 4.35,1.985 pfet_01v8_hvt
M$9 10 3 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=800000000000P
+ AD=540000000000P PS=5600000U PD=5080000U
* device instance $13 r0 *1 6.03,1.985 pfet_01v8_hvt
M$13 10 8 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=705000000000P PS=5080000U PD=6410000U
* device instance $17 r0 *1 4.35,0.56 nfet_01v8
M$17 6 3 7 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $21 r0 *1 6.03,0.56 nfet_01v8
M$21 1 8 7 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $25 r0 *1 0.47,0.56 nfet_01v8
M$25 1 5 4 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $29 r0 *1 2.15,0.56 nfet_01v8
M$29 6 2 4 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__a22oi_4

* cell sky130_fd_sc_hd__a21boi_4
* pin VGND
* pin Y
* pin B1_N
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a21boi_4 1 3 5 6 7 8 9 11
* net 1 VGND
* net 3 Y
* net 5 B1_N
* net 6 A2
* net 7 A1
* net 8 VPWR
* net 9 VPB
* device instance $1 r0 *1 1.455,1.985 pfet_01v8_hvt
M$1 3 2 10 9 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=575000000000P PS=6370000U PD=5150000U
* device instance $5 r0 *1 3.205,1.985 pfet_01v8_hvt
M$5 8 6 10 9 pfet_01v8_hvt L=150000U W=4000000U AS=575000000000P
+ AD=690000000000P PS=5150000U PD=6380000U
* device instance $6 r0 *1 3.645,1.985 pfet_01v8_hvt
M$6 10 7 8 9 pfet_01v8_hvt L=150000U W=4000000U AS=565000000000P
+ AD=560000000000P PS=5130000U PD=5120000U
* device instance $13 r0 *1 0.505,1.985 pfet_01v8_hvt
M$13 8 5 2 9 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=265000000000P PS=2530000U PD=2530000U
* device instance $14 r0 *1 0.625,0.56 nfet_01v8
M$14 1 5 2 11 nfet_01v8 L=150000U W=650000U AS=269750000000P AD=123500000000P
+ PS=2130000U PD=1030000U
* device instance $15 r0 *1 1.155,0.56 nfet_01v8
M$15 3 2 1 11 nfet_01v8 L=150000U W=2600000U AS=396500000000P AD=474500000000P
+ PS=3820000U PD=4060000U
* device instance $19 r0 *1 3.215,0.56 nfet_01v8
M$19 4 6 1 11 nfet_01v8 L=150000U W=2600000U AS=474500000000P AD=445250000000P
+ PS=4060000U PD=4620000U
* device instance $20 r0 *1 3.645,0.56 nfet_01v8
M$20 3 7 4 11 nfet_01v8 L=150000U W=2600000U AS=364000000000P AD=364000000000P
+ PS=3720000U PD=3720000U
.ENDS sky130_fd_sc_hd__a21boi_4

* cell sky130_fd_sc_hd__a41oi_4
* pin VGND
* pin B1
* pin A1
* pin A2
* pin Y
* pin A3
* pin A4
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a41oi_4 1 2 3 4 5 9 10 12 13 14
* net 1 VGND
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 Y
* net 9 A3
* net 10 A4
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 5 2 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=695000000000P PS=6330000U PD=5390000U
* device instance $5 r0 *1 2.46,1.985 pfet_01v8_hvt
M$5 12 3 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=865000000000P
+ AD=757500000000P PS=5730000U PD=5515000U
* device instance $9 r0 *1 4.575,1.985 pfet_01v8_hvt
M$9 12 4 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=790000000000P
+ AD=752500000000P PS=5580000U PD=5505000U
* device instance $13 r0 *1 6.68,1.985 pfet_01v8_hvt
M$13 12 9 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=550000000000P
+ AD=540000000000P PS=5100000U PD=5080000U
* device instance $17 r0 *1 8.36,1.985 pfet_01v8_hvt
M$17 12 10 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=695000000000P PS=5080000U PD=6390000U
* device instance $21 r0 *1 6.68,0.56 nfet_01v8
M$21 7 9 8 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $25 r0 *1 8.36,0.56 nfet_01v8
M$25 1 10 8 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=451750000000P
+ PS=3680000U PD=4640000U
* device instance $29 r0 *1 2.8,0.56 nfet_01v8
M$29 5 3 6 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $33 r0 *1 4.48,0.56 nfet_01v8
M$33 7 4 6 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $37 r0 *1 0.47,0.56 nfet_01v8
M$37 5 2 1 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=432250000000P
+ PS=4580000U PD=4580000U
.ENDS sky130_fd_sc_hd__a41oi_4

* cell sky130_fd_sc_hd__nand2b_4
* pin VGND
* pin B
* pin Y
* pin A_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand2b_4 1 2 5 6 7 8 9
* net 1 VGND
* net 2 B
* net 5 Y
* net 6 A_N
* net 7 VPWR
* net 8 VPB
* device instance $1 r0 *1 1.41,1.985 pfet_01v8_hvt
M$1 5 3 7 8 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=547500000000P PS=6330000U PD=5095000U
* device instance $5 r0 *1 3.105,1.985 pfet_01v8_hvt
M$5 5 2 7 8 pfet_01v8_hvt L=150000U W=4000000U AS=547500000000P
+ AD=795000000000P PS=5095000U PD=6590000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 7 6 3 8 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $10 r0 *1 1.41,0.56 nfet_01v8
M$10 5 3 4 9 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=355875000000P
+ PS=4580000U PD=3695000U
* device instance $14 r0 *1 3.105,0.56 nfet_01v8
M$14 1 2 4 9 nfet_01v8 L=150000U W=2600000U AS=355875000000P AD=516750000000P
+ PS=3695000U PD=4840000U
* device instance $18 r0 *1 0.47,0.56 nfet_01v8
M$18 1 6 3 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2b_4

* cell sky130_fd_sc_hd__o41ai_1
* pin VGND
* pin Y
* pin B1
* pin A4
* pin A3
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o41ai_1 1 2 4 5 6 7 8 9 10 14
* net 1 VGND
* net 2 Y
* net 4 B1
* net 5 A4
* net 6 A3
* net 7 A2
* net 8 A1
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 2 4 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 11 5 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=312500000000P PS=1270000U PD=1625000U
* device instance $3 r0 *1 1.665,1.985 pfet_01v8_hvt
M$3 13 6 11 10 pfet_01v8_hvt L=150000U W=1000000U AS=312500000000P
+ AD=135000000000P PS=1625000U PD=1270000U
* device instance $4 r0 *1 2.085,1.985 pfet_01v8_hvt
M$4 12 7 13 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=175000000000P PS=1270000U PD=1350000U
* device instance $5 r0 *1 2.585,1.985 pfet_01v8_hvt
M$5 9 8 12 10 pfet_01v8_hvt L=150000U W=1000000U AS=175000000000P
+ AD=280000000000P PS=1350000U PD=2560000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 3 4 2 14 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=203125000000P
+ PS=1820000U PD=1275000U
* device instance $7 r0 *1 1.245,0.56 nfet_01v8
M$7 1 5 3 14 nfet_01v8 L=150000U W=650000U AS=203125000000P AD=87750000000P
+ PS=1275000U PD=920000U
* device instance $8 r0 *1 1.665,0.56 nfet_01v8
M$8 3 6 1 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $9 r0 *1 2.085,0.56 nfet_01v8
M$9 1 7 3 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=113750000000P
+ PS=920000U PD=1000000U
* device instance $10 r0 *1 2.585,0.56 nfet_01v8
M$10 3 8 1 14 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=182000000000P
+ PS=1000000U PD=1860000U
.ENDS sky130_fd_sc_hd__o41ai_1

* cell sky130_fd_sc_hd__o32a_1
* pin VGND
* pin X
* pin A1
* pin A2
* pin A3
* pin B2
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o32a_1 1 2 5 6 7 8 9 10 11 15
* net 1 VGND
* net 2 X
* net 5 A1
* net 6 A2
* net 7 A3
* net 8 B2
* net 9 B1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.64,1.985 pfet_01v8_hvt
M$1 10 4 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=335000000000P
+ AD=135000000000P PS=2670000U PD=1270000U
* device instance $2 r0 *1 1.06,1.985 pfet_01v8_hvt
M$2 13 5 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $3 r0 *1 1.54,1.985 pfet_01v8_hvt
M$3 12 6 13 11 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=195000000000P PS=1330000U PD=1390000U
* device instance $4 r0 *1 2.08,1.985 pfet_01v8_hvt
M$4 4 7 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=195000000000P PS=1390000U PD=1390000U
* device instance $5 r0 *1 2.62,1.985 pfet_01v8_hvt
M$5 14 8 4 11 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=205000000000P PS=1390000U PD=1410000U
* device instance $6 r0 *1 3.18,1.985 pfet_01v8_hvt
M$6 10 9 14 11 pfet_01v8_hvt L=150000U W=1000000U AS=205000000000P
+ AD=290000000000P PS=1410000U PD=2580000U
* device instance $7 r0 *1 0.64,0.56 nfet_01v8
M$7 1 4 2 15 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 1.06,0.56 nfet_01v8
M$8 3 5 1 15 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $9 r0 *1 1.54,0.56 nfet_01v8
M$9 1 6 3 15 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=126750000000P
+ PS=980000U PD=1040000U
* device instance $10 r0 *1 2.08,0.56 nfet_01v8
M$10 3 7 1 15 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=126750000000P
+ PS=1040000U PD=1040000U
* device instance $11 r0 *1 2.62,0.56 nfet_01v8
M$11 4 8 3 15 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=133250000000P
+ PS=1040000U PD=1060000U
* device instance $12 r0 *1 3.18,0.56 nfet_01v8
M$12 3 9 4 15 nfet_01v8 L=150000U W=650000U AS=133250000000P AD=188500000000P
+ PS=1060000U PD=1880000U
.ENDS sky130_fd_sc_hd__o32a_1

* cell sky130_fd_sc_hd__mux2i_1
* pin VGND
* pin Y
* pin A0
* pin A1
* pin S
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2i_1 1 3 6 7 8 10 11 13
* net 1 VGND
* net 3 Y
* net 6 A0
* net 7 A1
* net 8 S
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 3.21,1.985 pfet_01v8_hvt
M$1 10 8 5 11 pfet_01v8_hvt L=150000U W=1000000U AS=290000000000P
+ AD=260000000000P PS=2580000U PD=2520000U
* device instance $2 r0 *1 0.49,1.985 pfet_01v8_hvt
M$2 3 6 9 11 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=152500000000P PS=2560000U PD=1305000U
* device instance $3 r0 *1 0.945,1.985 pfet_01v8_hvt
M$3 12 7 3 11 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=197500000000P PS=1305000U PD=1395000U
* device instance $4 r0 *1 1.49,1.985 pfet_01v8_hvt
M$4 10 5 12 11 pfet_01v8_hvt L=150000U W=1000000U AS=197500000000P
+ AD=300000000000P PS=1395000U PD=1600000U
* device instance $5 r0 *1 2.24,1.985 pfet_01v8_hvt
M$5 9 8 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=300000000000P
+ AD=260000000000P PS=1600000U PD=2520000U
* device instance $6 r0 *1 3.21,0.56 nfet_01v8
M$6 1 8 5 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
* device instance $7 r0 *1 1.85,0.56 nfet_01v8
M$7 1 5 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $8 r0 *1 2.27,0.56 nfet_01v8
M$8 4 8 1 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 3 6 2 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $10 r0 *1 0.89,0.56 nfet_01v8
M$10 4 7 3 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=182000000000P
+ PS=920000U PD=1860000U
.ENDS sky130_fd_sc_hd__mux2i_1

* cell sky130_fd_sc_hd__o22ai_1
* pin VPB
* pin B1
* pin B2
* pin A2
* pin A1
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o22ai_1 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 B1
* net 3 B2
* net 4 A2
* net 5 A1
* net 7 Y
* net 8 VGND
* net 9 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 12 2 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=112500000000P PS=2520000U PD=1225000U
* device instance $2 r0 *1 0.845,1.985 pfet_01v8_hvt
M$2 7 3 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=112500000000P
+ AD=232500000000P PS=1225000U PD=1465000U
* device instance $3 r0 *1 1.46,1.985 pfet_01v8_hvt
M$3 11 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=232500000000P
+ AD=105000000000P PS=1465000U PD=1210000U
* device instance $4 r0 *1 1.82,1.985 pfet_01v8_hvt
M$4 9 5 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=270000000000P PS=1210000U PD=2540000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 7 2 6 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=92625000000P
+ PS=1820000U PD=935000U
* device instance $6 r0 *1 0.905,0.56 nfet_01v8
M$6 6 3 7 10 nfet_01v8 L=150000U W=650000U AS=92625000000P AD=115375000000P
+ PS=935000U PD=1005000U
* device instance $7 r0 *1 1.41,0.56 nfet_01v8
M$7 8 4 6 10 nfet_01v8 L=150000U W=650000U AS=115375000000P AD=87750000000P
+ PS=1005000U PD=920000U
* device instance $8 r0 *1 1.83,0.56 nfet_01v8
M$8 6 5 8 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22ai_1

* cell sky130_fd_sc_hd__o22a_1
* pin VPB
* pin B1
* pin B2
* pin A2
* pin A1
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__o22a_1 1 2 3 4 5 6 7 10 11
* net 1 VPB
* net 2 B1
* net 3 B2
* net 4 A2
* net 5 A1
* net 6 X
* net 7 VGND
* net 10 VPWR
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 10 8 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=280000000000P
+ AD=372500000000P PS=2560000U PD=1745000U
* device instance $2 r0 *1 1.385,1.985 pfet_01v8_hvt
M$2 13 2 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=372500000000P
+ AD=117500000000P PS=1745000U PD=1235000U
* device instance $3 r0 *1 1.77,1.985 pfet_01v8_hvt
M$3 8 3 13 1 pfet_01v8_hvt L=150000U W=1000000U AS=117500000000P
+ AD=235000000000P PS=1235000U PD=1470000U
* device instance $4 r0 *1 2.39,1.985 pfet_01v8_hvt
M$4 12 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=235000000000P
+ AD=105000000000P PS=1470000U PD=1210000U
* device instance $5 r0 *1 2.75,1.985 pfet_01v8_hvt
M$5 10 5 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $6 r0 *1 1.41,0.56 nfet_01v8
M$6 8 2 9 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 1.83,0.56 nfet_01v8
M$7 9 3 8 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=113750000000P
+ PS=920000U PD=1000000U
* device instance $8 r0 *1 2.33,0.56 nfet_01v8
M$8 7 4 9 11 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=87750000000P
+ PS=1000000U PD=920000U
* device instance $9 r0 *1 2.75,0.56 nfet_01v8
M$9 9 5 7 11 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
* device instance $10 r0 *1 0.47,0.56 nfet_01v8
M$10 7 8 6 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22a_1

* cell sky130_fd_sc_hd__a22o_1
* pin VPB
* pin B2
* pin B1
* pin A1
* pin A2
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a22o_1 1 2 3 4 5 6 9 10 11
* net 1 VPB
* net 2 B2
* net 3 B1
* net 4 A1
* net 5 A2
* net 6 VGND
* net 9 X
* net 10 VPWR
* device instance $1 r0 *1 1.82,1.985 pfet_01v8_hvt
M$1 7 4 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=252900000000P
+ AD=160000000000P PS=2520000U PD=1320000U
* device instance $2 r0 *1 2.29,1.985 pfet_01v8_hvt
M$2 10 5 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=160000000000P
+ AD=155000000000P PS=1320000U PD=1310000U
* device instance $3 r0 *1 2.75,1.985 pfet_01v8_hvt
M$3 9 8 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=155000000000P
+ AD=260000000000P PS=1310000U PD=2520000U
* device instance $4 r0 *1 0.47,1.985 pfet_01v8_hvt
M$4 7 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $5 r0 *1 0.89,1.985 pfet_01v8_hvt
M$5 8 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=252850000000P PS=1270000U PD=2520000U
* device instance $6 r0 *1 1.79,0.56 nfet_01v8
M$6 12 4 8 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=113750000000P
+ PS=1820000U PD=1000000U
* device instance $7 r0 *1 2.29,0.56 nfet_01v8
M$7 6 5 12 11 nfet_01v8 L=150000U W=650000U AS=113750000000P AD=100750000000P
+ PS=1000000U PD=960000U
* device instance $8 r0 *1 2.75,0.56 nfet_01v8
M$8 9 8 6 11 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=169000000000P
+ PS=960000U PD=1820000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 13 2 6 11 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=74750000000P
+ PS=1820000U PD=880000U
* device instance $10 r0 *1 0.85,0.56 nfet_01v8
M$10 8 3 13 11 nfet_01v8 L=150000U W=650000U AS=74750000000P AD=169000000000P
+ PS=880000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22o_1

* cell sky130_fd_sc_hd__nor3_2
* pin VGND
* pin A
* pin Y
* pin B
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor3_2 1 2 3 4 5 7 9 10
* net 1 VGND
* net 2 A
* net 3 Y
* net 4 B
* net 5 C
* net 7 VPWR
* net 9 VPB
* device instance $1 r0 *1 2.71,1.985 pfet_01v8_hvt
M$1 3 5 8 9 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=395000000000P PS=3790000U PD=3790000U
* device instance $3 r0 *1 0.49,1.985 pfet_01v8_hvt
M$3 7 2 6 9 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $5 r0 *1 1.33,1.985 pfet_01v8_hvt
M$5 8 4 6 9 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $7 r0 *1 2.71,0.56 nfet_01v8
M$7 3 5 1 10 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
* device instance $9 r0 *1 0.49,0.56 nfet_01v8
M$9 3 2 1 10 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=175500000000P
+ PS=2770000U PD=1840000U
* device instance $11 r0 *1 1.33,0.56 nfet_01v8
M$11 3 4 1 10 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nor3_2

* cell sky130_fd_sc_hd__mux2i_4
* pin VGND
* pin A0
* pin Y
* pin A1
* pin S
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2i_4 1 2 3 7 8 10 11 13
* net 1 VGND
* net 2 A0
* net 3 Y
* net 7 A1
* net 8 S
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 4.35,1.985 pfet_01v8_hvt
M$1 9 8 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 6.03,1.985 pfet_01v8_hvt
M$5 12 6 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=567500000000P
+ AD=590000000000P PS=5135000U PD=5180000U
* device instance $9 r0 *1 7.81,1.985 pfet_01v8_hvt
M$9 6 8 10 11 pfet_01v8_hvt L=150000U W=1000000U AS=157500000000P
+ AD=260000000000P PS=1315000U PD=2520000U
* device instance $10 r0 *1 0.47,1.985 pfet_01v8_hvt
M$10 9 2 3 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $14 r0 *1 2.15,1.985 pfet_01v8_hvt
M$14 12 7 3 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $18 r0 *1 4.35,0.56 nfet_01v8
M$18 5 8 1 13 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $22 r0 *1 6.03,0.56 nfet_01v8
M$22 4 6 1 13 nfet_01v8 L=150000U W=2600000U AS=368875000000P AD=383500000000P
+ PS=3735000U PD=3780000U
* device instance $26 r0 *1 7.81,0.56 nfet_01v8
M$26 6 8 1 13 nfet_01v8 L=150000U W=650000U AS=102375000000P AD=169000000000P
+ PS=965000U PD=1820000U
* device instance $27 r0 *1 0.47,0.56 nfet_01v8
M$27 4 2 3 13 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $31 r0 *1 2.15,0.56 nfet_01v8
M$31 5 7 3 13 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__mux2i_4

* cell sky130_fd_sc_hd__o211ai_4
* pin VGND
* pin A1
* pin A2
* pin C1
* pin B1
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o211ai_4 1 2 3 4 6 10 11 12 14
* net 1 VGND
* net 2 A1
* net 3 A2
* net 4 C1
* net 6 B1
* net 10 VPWR
* net 11 Y
* net 12 VPB
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 13 2 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=580000000000P PS=6370000U PD=5160000U
* device instance $4 r0 *1 1.765,1.985 pfet_01v8_hvt
M$4 11 3 13 12 pfet_01v8_hvt L=150000U W=4000000U AS=560000000000P
+ AD=560000000000P PS=5120000U PD=5120000U
* device instance $9 r0 *1 3.955,1.985 pfet_01v8_hvt
M$9 11 6 10 12 pfet_01v8_hvt L=150000U W=4000000U AS=575000000000P AD=1.09e+12P
+ PS=5150000U PD=7180000U
* device instance $12 r0 *1 5.235,1.985 pfet_01v8_hvt
M$12 10 4 11 12 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $17 r0 *1 0.475,0.56 nfet_01v8
M$17 1 2 5 14 nfet_01v8 L=150000U W=2600000U AS=448500000000P AD=373750000000P
+ PS=4630000U PD=3750000U
* device instance $20 r0 *1 1.765,0.56 nfet_01v8
M$20 5 3 1 14 nfet_01v8 L=150000U W=2600000U AS=364000000000P AD=367250000000P
+ PS=3720000U PD=3730000U
* device instance $25 r0 *1 3.955,0.56 nfet_01v8
M$25 7 6 5 14 nfet_01v8 L=150000U W=1300000U AS=191750000000P AD=182000000000P
+ PS=1890000U PD=1860000U
* device instance $27 r0 *1 4.815,0.56 nfet_01v8
M$27 9 6 5 14 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=87750000000P
+ PS=930000U PD=920000U
* device instance $28 r0 *1 5.235,0.56 nfet_01v8
M$28 11 4 9 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $29 r0 *1 5.655,0.56 nfet_01v8
M$29 7 4 11 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $31 r0 *1 6.495,0.56 nfet_01v8
M$31 8 4 11 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=104000000000P
+ PS=920000U PD=970000U
* device instance $32 r0 *1 6.965,0.56 nfet_01v8
M$32 5 6 8 14 nfet_01v8 L=150000U W=650000U AS=104000000000P AD=256750000000P
+ PS=970000U PD=2090000U
.ENDS sky130_fd_sc_hd__o211ai_4

* cell sky130_fd_sc_hd__a221oi_1
* pin VGND
* pin Y
* pin B1
* pin A1
* pin C1
* pin B2
* pin A2
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a221oi_1 1 2 3 4 5 6 7 10 11 14
* net 1 VGND
* net 2 Y
* net 3 B1
* net 4 A1
* net 5 C1
* net 6 B2
* net 7 A2
* net 10 VPB
* net 11 VPWR
* device instance $1 r0 *1 2.25,1.985 pfet_01v8_hvt
M$1 13 4 11 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=152500000000P PS=2520000U PD=1305000U
* device instance $2 r0 *1 2.705,1.985 pfet_01v8_hvt
M$2 11 7 13 10 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=305000000000P PS=1305000U PD=2610000U
* device instance $3 r0 *1 0.47,1.985 pfet_01v8_hvt
M$3 12 5 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $4 r0 *1 0.89,1.985 pfet_01v8_hvt
M$4 13 6 12 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $5 r0 *1 1.31,1.985 pfet_01v8_hvt
M$5 12 3 13 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $6 r0 *1 2.25,0.56 nfet_01v8
M$6 9 4 2 14 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=99125000000P
+ PS=1820000U PD=955000U
* device instance $7 r0 *1 2.705,0.56 nfet_01v8
M$7 1 7 9 14 nfet_01v8 L=150000U W=650000U AS=99125000000P AD=198250000000P
+ PS=955000U PD=1910000U
* device instance $8 r0 *1 0.47,0.56 nfet_01v8
M$8 1 5 2 14 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=105625000000P
+ PS=1820000U PD=975000U
* device instance $9 r0 *1 0.945,0.56 nfet_01v8
M$9 8 6 1 14 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=69875000000P
+ PS=975000U PD=865000U
* device instance $10 r0 *1 1.31,0.56 nfet_01v8
M$10 2 3 8 14 nfet_01v8 L=150000U W=650000U AS=69875000000P AD=169000000000P
+ PS=865000U PD=1820000U
.ENDS sky130_fd_sc_hd__a221oi_1

* cell sky130_fd_sc_hd__and3_2
* pin VPB
* pin A
* pin B
* pin C
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__and3_2 1 2 3 4 6 7 8 9
* net 1 VPB
* net 2 A
* net 3 B
* net 4 C
* net 6 VGND
* net 7 VPWR
* net 8 X
* device instance $1 r0 *1 1.375,1.695 pfet_01v8_hvt
M$1 7 4 5 1 pfet_01v8_hvt L=150000U W=420000U AS=74375000000P AD=150750000000P
+ PS=815000U PD=1345000U
* device instance $2 r0 *1 0.48,1.765 pfet_01v8_hvt
M$2 7 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $3 r0 *1 0.9,1.765 pfet_01v8_hvt
M$3 7 3 5 1 pfet_01v8_hvt L=150000U W=420000U AS=74375000000P AD=56700000000P
+ PS=815000U PD=690000U
* device instance $4 r0 *1 1.87,1.985 pfet_01v8_hvt
M$4 8 5 7 1 pfet_01v8_hvt L=150000U W=2000000U AS=285750000000P
+ AD=395000000000P PS=2615000U PD=3790000U
* device instance $6 r0 *1 0.485,0.475 nfet_01v8
M$6 11 2 5 9 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $7 r0 *1 0.845,0.475 nfet_01v8
M$7 10 3 11 9 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=53550000000P
+ PS=630000U PD=675000U
* device instance $8 r0 *1 1.25,0.475 nfet_01v8
M$8 10 4 6 9 nfet_01v8 L=150000U W=420000U AS=130400000000P AD=53550000000P
+ PS=1105000U PD=675000U
* device instance $9 r0 *1 1.855,0.56 nfet_01v8
M$9 8 5 6 9 nfet_01v8 L=150000U W=1300000U AS=218150000000P AD=266500000000P
+ PS=2025000U PD=2770000U
.ENDS sky130_fd_sc_hd__and3_2

* cell sky130_fd_sc_hd__o2111a_1
* pin VGND
* pin X
* pin C1
* pin B1
* pin D1
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o2111a_1 1 2 4 5 7 8 9 12 13 14
* net 1 VGND
* net 2 X
* net 4 C1
* net 5 B1
* net 7 D1
* net 8 A2
* net 9 A1
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 12 3 2 13 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=382500000000P PS=2520000U PD=1765000U
* device instance $2 r0 *1 1.385,1.985 pfet_01v8_hvt
M$2 3 7 12 13 pfet_01v8_hvt L=150000U W=1000000U AS=382500000000P
+ AD=217500000000P PS=1765000U PD=1435000U
* device instance $3 r0 *1 1.97,1.985 pfet_01v8_hvt
M$3 12 4 3 13 pfet_01v8_hvt L=150000U W=1000000U AS=217500000000P
+ AD=305000000000P PS=1435000U PD=1610000U
* device instance $4 r0 *1 2.73,1.985 pfet_01v8_hvt
M$4 3 5 12 13 pfet_01v8_hvt L=150000U W=1000000U AS=305000000000P
+ AD=212500000000P PS=1610000U PD=1425000U
* device instance $5 r0 *1 3.305,1.985 pfet_01v8_hvt
M$5 15 8 3 13 pfet_01v8_hvt L=150000U W=1000000U AS=212500000000P
+ AD=105000000000P PS=1425000U PD=1210000U
* device instance $6 r0 *1 3.665,1.985 pfet_01v8_hvt
M$6 12 9 15 13 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=265000000000P PS=1210000U PD=2530000U
* device instance $7 r0 *1 1.455,0.56 nfet_01v8
M$7 11 7 3 14 nfet_01v8 L=150000U W=650000U AS=198250000000P AD=118625000000P
+ PS=1910000U PD=1015000U
* device instance $8 r0 *1 1.97,0.56 nfet_01v8
M$8 10 4 11 14 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=118625000000P
+ PS=1015000U PD=1015000U
* device instance $9 r0 *1 2.485,0.56 nfet_01v8
M$9 6 5 10 14 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=198250000000P
+ PS=1015000U PD=1260000U
* device instance $10 r0 *1 3.245,0.56 nfet_01v8
M$10 1 8 6 14 nfet_01v8 L=150000U W=650000U AS=198250000000P AD=87750000000P
+ PS=1260000U PD=920000U
* device instance $11 r0 *1 3.665,0.56 nfet_01v8
M$11 6 9 1 14 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=172250000000P
+ PS=920000U PD=1830000U
* device instance $12 r0 *1 0.47,0.56 nfet_01v8
M$12 1 3 2 14 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__o2111a_1

* cell sky130_fd_sc_hd__o211ai_2
* pin VGND
* pin Y
* pin A1
* pin C1
* pin B1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o211ai_2 1 3 5 6 7 8 9 11 12
* net 1 VGND
* net 3 Y
* net 5 A1
* net 6 C1
* net 7 B1
* net 8 A2
* net 9 VPWR
* net 11 VPB
* device instance $1 r0 *1 2.775,1.985 pfet_01v8_hvt
M$1 3 8 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=280000000000P PS=3810000U PD=2560000U
* device instance $3 r0 *1 3.635,1.985 pfet_01v8_hvt
M$3 9 5 10 11 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=405000000000P PS=2560000U PD=3810000U
* device instance $5 r0 *1 0.495,1.985 pfet_01v8_hvt
M$5 3 6 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=280000000000P PS=3810000U PD=2560000U
* device instance $7 r0 *1 1.355,1.985 pfet_01v8_hvt
M$7 3 7 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=405000000000P PS=2560000U PD=3810000U
* device instance $9 r0 *1 2.775,0.56 nfet_01v8
M$9 4 8 1 12 nfet_01v8 L=150000U W=1300000U AS=276250000000P AD=182000000000P
+ PS=2800000U PD=1860000U
* device instance $11 r0 *1 3.635,0.56 nfet_01v8
M$11 4 5 1 12 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=276250000000P
+ PS=1860000U PD=2800000U
* device instance $13 r0 *1 0.495,0.56 nfet_01v8
M$13 3 6 2 12 nfet_01v8 L=150000U W=1300000U AS=276250000000P AD=182000000000P
+ PS=2800000U PD=1860000U
* device instance $15 r0 *1 1.355,0.56 nfet_01v8
M$15 4 7 2 12 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=276250000000P
+ PS=1860000U PD=2800000U
.ENDS sky130_fd_sc_hd__o211ai_2

* cell sky130_fd_sc_hd__xnor2_2
* pin VGND
* pin Y
* pin B
* pin A
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__xnor2_2 1 5 6 7 8 9 11
* net 1 VGND
* net 5 Y
* net 6 B
* net 7 A
* net 8 VPB
* net 9 VPWR
* device instance $1 r0 *1 4.96,1.985 pfet_01v8_hvt
M$1 5 3 9 8 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=415000000000P PS=3790000U PD=3830000U
* device instance $3 r0 *1 2.725,1.985 pfet_01v8_hvt
M$3 9 7 10 8 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $5 r0 *1 3.565,1.985 pfet_01v8_hvt
M$5 5 6 10 8 pfet_01v8_hvt L=150000U W=2000000U AS=287500000000P
+ AD=412500000000P PS=2575000U PD=3825000U
* device instance $7 r0 *1 0.485,1.985 pfet_01v8_hvt
M$7 9 6 3 8 pfet_01v8_hvt L=150000U W=2000000U AS=410000000000P
+ AD=270000000000P PS=3820000U PD=2540000U
* device instance $9 r0 *1 1.325,1.985 pfet_01v8_hvt
M$9 9 7 3 8 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $11 r0 *1 4.96,0.56 nfet_01v8
M$11 4 3 5 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
* device instance $13 r0 *1 2.725,0.56 nfet_01v8
M$13 4 7 1 11 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $15 r0 *1 3.565,0.56 nfet_01v8
M$15 4 6 1 11 nfet_01v8 L=150000U W=1300000U AS=186875000000P AD=268125000000P
+ PS=1875000U PD=2775000U
* device instance $17 r0 *1 0.485,0.56 nfet_01v8
M$17 3 6 2 11 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=175500000000P
+ PS=2770000U PD=1840000U
* device instance $19 r0 *1 1.325,0.56 nfet_01v8
M$19 1 7 2 11 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
.ENDS sky130_fd_sc_hd__xnor2_2

* cell sky130_fd_sc_hd__o311ai_4
* pin VGND
* pin A1
* pin A2
* pin A3
* pin B1
* pin C1
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311ai_4 1 2 4 5 7 8 10 12 13 14
* net 1 VGND
* net 2 A1
* net 4 A2
* net 5 A3
* net 7 B1
* net 8 C1
* net 10 VPWR
* net 12 Y
* net 13 VPB
* device instance $1 r0 *1 4.43,1.985 pfet_01v8_hvt
M$1 11 5 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=550000000000P PS=6330000U PD=5100000U
* device instance $5 r0 *1 6.13,1.985 pfet_01v8_hvt
M$5 10 7 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=550000000000P
+ AD=540000000000P PS=5100000U PD=5080000U
* device instance $9 r0 *1 7.81,1.985 pfet_01v8_hvt
M$9 10 8 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $13 r0 *1 0.55,1.985 pfet_01v8_hvt
M$13 10 2 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $17 r0 *1 2.23,1.985 pfet_01v8_hvt
M$17 11 4 9 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 6.17,0.56 nfet_01v8
M$21 3 7 6 14 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $25 r0 *1 7.85,0.56 nfet_01v8
M$25 12 8 6 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=445250000000P
+ PS=3680000U PD=4620000U
* device instance $29 r0 *1 0.55,0.56 nfet_01v8
M$29 3 2 1 14 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $33 r0 *1 2.23,0.56 nfet_01v8
M$33 3 4 1 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=357500000000P
+ PS=3680000U PD=3700000U
* device instance $37 r0 *1 3.93,0.56 nfet_01v8
M$37 3 5 1 14 nfet_01v8 L=150000U W=2600000U AS=357500000000P AD=445250000000P
+ PS=3700000U PD=4620000U
.ENDS sky130_fd_sc_hd__o311ai_4

* cell sky130_fd_sc_hd__and2_2
* pin VPB
* pin A
* pin B
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__and2_2 1 2 3 5 6 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 5 VPWR
* net 6 X
* net 7 VGND
* device instance $1 r0 *1 0.66,2.065 pfet_01v8_hvt
M$1 4 2 5 1 pfet_01v8_hvt L=150000U W=420000U AS=117600000000P AD=56700000000P
+ PS=1400000U PD=690000U
* device instance $2 r0 *1 1.08,2.065 pfet_01v8_hvt
M$2 4 3 5 1 pfet_01v8_hvt L=150000U W=420000U AS=166550000000P AD=56700000000P
+ PS=1390000U PD=690000U
* device instance $3 r0 *1 1.62,1.985 pfet_01v8_hvt
M$3 6 4 5 1 pfet_01v8_hvt L=150000U W=2000000U AS=361550000000P
+ AD=575000000000P PS=2780000U PD=4150000U
* device instance $5 r0 *1 0.66,0.585 nfet_01v8
M$5 9 2 4 8 nfet_01v8 L=150000U W=420000U AS=117600000000P AD=56700000000P
+ PS=1400000U PD=690000U
* device instance $6 r0 *1 1.08,0.585 nfet_01v8
M$6 9 3 7 8 nfet_01v8 L=150000U W=420000U AS=111800000000P AD=56700000000P
+ PS=1040000U PD=690000U
* device instance $7 r0 *1 1.62,0.56 nfet_01v8
M$7 6 4 7 8 nfet_01v8 L=150000U W=1300000U AS=238550000000P AD=373750000000P
+ PS=2080000U PD=3100000U
.ENDS sky130_fd_sc_hd__and2_2

* cell sky130_fd_sc_hd__o311ai_2
* pin VGND
* pin Y
* pin A1
* pin A2
* pin A3
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o311ai_2 1 4 5 6 7 8 9 11 13 14
* net 1 VGND
* net 4 Y
* net 5 A1
* net 6 A2
* net 7 A3
* net 8 B1
* net 9 C1
* net 11 VPWR
* net 13 VPB
* device instance $1 r0 *1 2.79,1.985 pfet_01v8_hvt
M$1 12 7 4 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 3.63,1.985 pfet_01v8_hvt
M$3 11 8 4 13 pfet_01v8_hvt L=150000U W=2000000U AS=440000000000P
+ AD=510000000000P PS=2880000U PD=3020000U
* device instance $5 r0 *1 4.95,1.985 pfet_01v8_hvt
M$5 11 9 4 13 pfet_01v8_hvt L=150000U W=2000000U AS=340000000000P
+ AD=395000000000P PS=2680000U PD=3790000U
* device instance $7 r0 *1 0.59,1.985 pfet_01v8_hvt
M$7 11 5 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $9 r0 *1 1.43,1.985 pfet_01v8_hvt
M$9 12 6 10 13 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $11 r0 *1 4.97,0.56 nfet_01v8
M$11 3 9 4 14 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=256750000000P
+ PS=2780000U PD=2740000U
* device instance $13 r0 *1 0.61,0.56 nfet_01v8
M$13 1 5 2 14 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $15 r0 *1 1.45,0.56 nfet_01v8
M$15 1 6 2 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $17 r0 *1 2.29,0.56 nfet_01v8
M$17 1 7 2 14 nfet_01v8 L=150000U W=1300000U AS=318500000000P AD=318500000000P
+ PS=2280000U PD=2280000U
* device instance $19 r0 *1 3.57,0.56 nfet_01v8
M$19 3 8 2 14 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
.ENDS sky130_fd_sc_hd__o311ai_2

* cell sky130_fd_sc_hd__a311oi_4
* pin VGND
* pin A3
* pin C1
* pin A2
* pin A1
* pin Y
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a311oi_4 1 2 3 5 7 8 9 10 13 14
* net 1 VGND
* net 2 A3
* net 3 C1
* net 5 A2
* net 7 A1
* net 8 Y
* net 9 B1
* net 10 VPWR
* net 13 VPB
* device instance $1 r0 *1 6.03,1.985 pfet_01v8_hvt
M$1 11 9 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=650000000000P PS=6330000U PD=5300000U
* device instance $5 r0 *1 7.93,1.985 pfet_01v8_hvt
M$5 8 3 12 13 pfet_01v8_hvt L=150000U W=4000000U AS=650000000000P
+ AD=665000000000P PS=5300000U PD=6330000U
* device instance $9 r0 *1 0.47,1.985 pfet_01v8_hvt
M$9 11 2 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $13 r0 *1 2.15,1.985 pfet_01v8_hvt
M$13 11 5 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $17 r0 *1 3.83,1.985 pfet_01v8_hvt
M$17 11 7 10 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 4.35,0.56 nfet_01v8
M$21 6 7 8 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $25 r0 *1 6.03,0.56 nfet_01v8
M$25 1 9 8 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=422500000000P
+ PS=3680000U PD=3900000U
* device instance $29 r0 *1 7.93,0.56 nfet_01v8
M$29 1 3 8 14 nfet_01v8 L=150000U W=2600000U AS=422500000000P AD=432250000000P
+ PS=3900000U PD=4580000U
* device instance $33 r0 *1 0.47,0.56 nfet_01v8
M$33 1 2 4 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $37 r0 *1 2.15,0.56 nfet_01v8
M$37 6 5 4 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__a311oi_4

* cell sky130_fd_sc_hd__o2111ai_2
* pin VGND
* pin D1
* pin Y
* pin C1
* pin B1
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o2111ai_2 1 2 4 5 7 9 10 11 13 14
* net 1 VGND
* net 2 D1
* net 4 Y
* net 5 C1
* net 7 B1
* net 9 A2
* net 10 A1
* net 11 VPWR
* net 13 VPB
* device instance $1 r0 *1 3.69,1.985 pfet_01v8_hvt
M$1 4 9 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=435000000000P
+ AD=280000000000P PS=3870000U PD=2560000U
* device instance $3 r0 *1 4.55,1.985 pfet_01v8_hvt
M$3 11 10 12 13 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=470000000000P PS=2560000U PD=3940000U
* device instance $5 r0 *1 0.555,1.985 pfet_01v8_hvt
M$5 4 2 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=280000000000P PS=3810000U PD=2560000U
* device instance $7 r0 *1 1.415,1.985 pfet_01v8_hvt
M$7 4 5 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=280000000000P PS=2560000U PD=2560000U
* device instance $9 r0 *1 2.275,1.985 pfet_01v8_hvt
M$9 4 7 11 13 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=405000000000P PS=2560000U PD=3810000U
* device instance $11 r0 *1 2.83,0.56 nfet_01v8
M$11 6 7 8 14 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=182000000000P
+ PS=2770000U PD=1860000U
* device instance $13 r0 *1 3.69,0.56 nfet_01v8
M$13 1 9 8 14 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=182000000000P
+ PS=1860000U PD=1860000U
* device instance $15 r0 *1 4.55,0.56 nfet_01v8
M$15 1 10 8 14 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=305500000000P
+ PS=1860000U PD=2890000U
* device instance $17 r0 *1 0.555,0.56 nfet_01v8
M$17 4 2 3 14 nfet_01v8 L=150000U W=1300000U AS=315250000000P AD=182000000000P
+ PS=2920000U PD=1860000U
* device instance $19 r0 *1 1.415,0.56 nfet_01v8
M$19 6 5 3 14 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=282750000000P
+ PS=1860000U PD=2820000U
.ENDS sky130_fd_sc_hd__o2111ai_2

* cell sky130_fd_sc_hd__buf_6
* pin VGND
* pin A
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__buf_6 1 2 4 5 6 7
* net 1 VGND
* net 2 A
* net 4 X
* net 5 VPWR
* net 6 VPB
* device instance $1 r0 *1 0.73,1.985 pfet_01v8_hvt
M$1 3 2 5 6 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.57,1.985 pfet_01v8_hvt
M$3 4 3 5 6 pfet_01v8_hvt L=150000U W=6000000U AS=810000000000P
+ AD=935000000000P PS=7620000U PD=8870000U
* device instance $9 r0 *1 0.73,0.56 nfet_01v8
M$9 3 2 1 7 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $11 r0 *1 1.57,0.56 nfet_01v8
M$11 4 3 1 7 nfet_01v8 L=150000U W=3900000U AS=526500000000P AD=607750000000P
+ PS=5520000U PD=6420000U
.ENDS sky130_fd_sc_hd__buf_6

* cell sky130_fd_sc_hd__nor4b_2
* pin VGND
* pin Y
* pin A
* pin B
* pin C
* pin D_N
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor4b_2 1 2 4 5 6 7 11 12 13
* net 1 VGND
* net 2 Y
* net 4 A
* net 5 B
* net 6 C
* net 7 D_N
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 2.705,1.985 pfet_01v8_hvt
M$1 9 6 10 12 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 3.545,1.985 pfet_01v8_hvt
M$3 2 3 10 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 11 4 8 12 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $7 r0 *1 1.31,1.985 pfet_01v8_hvt
M$7 9 5 8 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $9 r0 *1 4.905,2.275 pfet_01v8_hvt
M$9 11 7 3 12 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=109200000000P PS=1360000U PD=1360000U
* device instance $10 r0 *1 4.905,0.675 nfet_01v8
M$10 1 7 3 13 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
* device instance $11 r0 *1 2.705,0.56 nfet_01v8
M$11 2 6 1 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $13 r0 *1 3.545,0.56 nfet_01v8
M$13 2 3 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
* device instance $15 r0 *1 0.47,0.56 nfet_01v8
M$15 2 4 1 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $17 r0 *1 1.31,0.56 nfet_01v8
M$17 2 5 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nor4b_2

* cell sky130_fd_sc_hd__o211ai_1
* pin VPB
* pin A1
* pin A2
* pin B1
* pin C1
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o211ai_1 1 2 3 4 5 7 8 9 10
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 B1
* net 5 C1
* net 7 Y
* net 8 VPWR
* net 9 VGND
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 11 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=105000000000P PS=2530000U PD=1210000U
* device instance $2 r0 *1 0.835,1.985 pfet_01v8_hvt
M$2 7 3 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=195000000000P PS=1210000U PD=1390000U
* device instance $3 r0 *1 1.375,1.985 pfet_01v8_hvt
M$3 8 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=195000000000P PS=1390000U PD=1390000U
* device instance $4 r0 *1 1.915,1.985 pfet_01v8_hvt
M$4 7 5 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=635000000000P PS=1390000U PD=3270000U
* device instance $5 r0 *1 0.475,0.56 nfet_01v8
M$5 9 2 6 10 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=126750000000P
+ PS=1830000U PD=1040000U
* device instance $6 r0 *1 1.015,0.56 nfet_01v8
M$6 6 3 9 10 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=126750000000P
+ PS=1040000U PD=1040000U
* device instance $7 r0 *1 1.555,0.56 nfet_01v8
M$7 12 4 6 10 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=68250000000P
+ PS=1040000U PD=860000U
* device instance $8 r0 *1 1.915,0.56 nfet_01v8
M$8 7 5 12 10 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=393250000000P
+ PS=860000U PD=2510000U
.ENDS sky130_fd_sc_hd__o211ai_1

* cell sky130_fd_sc_hd__nor3_4
* pin VGND
* pin A
* pin Y
* pin B
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nor3_4 1 2 3 4 5 7 9 10
* net 1 VGND
* net 2 A
* net 3 Y
* net 4 B
* net 5 C
* net 7 VPWR
* net 9 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 7 2 6 9 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $5 r0 *1 2.17,1.985 pfet_01v8_hvt
M$5 8 4 6 9 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $8 r0 *1 3.43,1.985 pfet_01v8_hvt
M$8 3 5 8 9 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $13 r0 *1 0.49,0.56 nfet_01v8
M$13 3 2 1 10 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $17 r0 *1 2.17,0.56 nfet_01v8
M$17 3 4 1 10 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $20 r0 *1 3.43,0.56 nfet_01v8
M$20 1 5 3 10 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
.ENDS sky130_fd_sc_hd__nor3_4

* cell sky130_fd_sc_hd__a211oi_2
* pin VGND
* pin Y
* pin C1
* pin B1
* pin A1
* pin A2
* pin VPB
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a211oi_2 1 2 4 5 6 7 10 11 12
* net 1 VGND
* net 2 Y
* net 4 C1
* net 5 B1
* net 6 A1
* net 7 A2
* net 10 VPB
* net 11 VPWR
* device instance $1 r0 *1 2.765,1.985 pfet_01v8_hvt
M$1 9 6 11 10 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=280000000000P PS=3810000U PD=2560000U
* device instance $3 r0 *1 3.625,1.985 pfet_01v8_hvt
M$3 9 7 11 10 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=405000000000P PS=2560000U PD=3810000U
* device instance $5 r0 *1 0.525,1.985 pfet_01v8_hvt
M$5 2 4 8 10 pfet_01v8_hvt L=150000U W=2000000U AS=405000000000P
+ AD=280000000000P PS=3810000U PD=2560000U
* device instance $7 r0 *1 1.385,1.985 pfet_01v8_hvt
M$7 9 5 8 10 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=405000000000P PS=2560000U PD=3810000U
* device instance $9 r0 *1 2.765,0.56 nfet_01v8
M$9 2 6 3 12 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=182000000000P
+ PS=2760000U PD=1860000U
* device instance $11 r0 *1 3.625,0.56 nfet_01v8
M$11 1 7 3 12 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=263250000000P
+ PS=1860000U PD=2760000U
* device instance $13 r0 *1 0.525,0.56 nfet_01v8
M$13 2 4 1 12 nfet_01v8 L=150000U W=1300000U AS=263250000000P AD=182000000000P
+ PS=2760000U PD=1860000U
* device instance $15 r0 *1 1.385,0.56 nfet_01v8
M$15 2 5 1 12 nfet_01v8 L=150000U W=1300000U AS=182000000000P AD=263250000000P
+ PS=1860000U PD=2760000U
.ENDS sky130_fd_sc_hd__a211oi_2

* cell sky130_fd_sc_hd__a211oi_1
* pin VPB
* pin A2
* pin A1
* pin C1
* pin B1
* pin VGND
* pin Y
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__a211oi_1 1 2 3 4 5 6 7 9 10
* net 1 VPB
* net 2 A2
* net 3 A1
* net 4 C1
* net 5 B1
* net 6 VGND
* net 7 Y
* net 9 VPWR
* device instance $1 r0 *1 0.62,1.985 pfet_01v8_hvt
M$1 9 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 1.05,1.985 pfet_01v8_hvt
M$2 8 3 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=140000000000P PS=1280000U PD=1280000U
* device instance $3 r0 *1 1.48,1.985 pfet_01v8_hvt
M$3 11 5 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=155000000000P PS=1280000U PD=1310000U
* device instance $4 r0 *1 1.94,1.985 pfet_01v8_hvt
M$4 7 4 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=155000000000P
+ AD=265000000000P PS=1310000U PD=2530000U
* device instance $5 r0 *1 0.62,0.56 nfet_01v8
M$5 12 2 6 10 nfet_01v8 L=150000U W=650000U AS=266500000000P AD=91000000000P
+ PS=2120000U PD=930000U
* device instance $6 r0 *1 1.05,0.56 nfet_01v8
M$6 7 3 12 10 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=91000000000P
+ PS=930000U PD=930000U
* device instance $7 r0 *1 1.48,0.56 nfet_01v8
M$7 6 5 7 10 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=100750000000P
+ PS=930000U PD=960000U
* device instance $8 r0 *1 1.94,0.56 nfet_01v8
M$8 7 4 6 10 nfet_01v8 L=150000U W=650000U AS=100750000000P AD=172250000000P
+ PS=960000U PD=1830000U
.ENDS sky130_fd_sc_hd__a211oi_1

* cell sky130_fd_sc_hd__a32oi_4
* pin VGND
* pin B2
* pin B1
* pin A2
* pin Y
* pin A1
* pin A3
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a32oi_4 1 2 3 4 6 7 10 12 13 14
* net 1 VGND
* net 2 B2
* net 3 B1
* net 4 A2
* net 6 Y
* net 7 A1
* net 10 A3
* net 12 VPWR
* net 13 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 6 2 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 6 3 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=550000000000P PS=5080000U PD=5100000U
* device instance $9 r0 *1 3.85,1.985 pfet_01v8_hvt
M$9 12 7 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=752500000000P
+ AD=860000000000P PS=5505000U PD=5720000U
* device instance $13 r0 *1 6.17,1.985 pfet_01v8_hvt
M$13 12 4 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=657500000000P
+ AD=800000000000P PS=5315000U PD=5600000U
* device instance $17 r0 *1 8.37,1.985 pfet_01v8_hvt
M$17 12 10 11 13 pfet_01v8_hvt L=150000U W=4000000U AS=800000000000P
+ AD=665000000000P PS=5600000U PD=6330000U
* device instance $21 r0 *1 8.37,0.56 nfet_01v8
M$21 9 10 1 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=445250000000P
+ PS=4580000U PD=4620000U
* device instance $25 r0 *1 4.35,0.56 nfet_01v8
M$25 6 7 8 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=396500000000P
+ PS=4580000U PD=3820000U
* device instance $29 r0 *1 6.17,0.56 nfet_01v8
M$29 9 4 8 14 nfet_01v8 L=150000U W=2600000U AS=396500000000P AD=432250000000P
+ PS=3820000U PD=4580000U
* device instance $33 r0 *1 0.47,0.56 nfet_01v8
M$33 1 2 5 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $37 r0 *1 2.15,0.56 nfet_01v8
M$37 6 3 5 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__a32oi_4

* cell sky130_fd_sc_hd__o21ai_4
* pin VGND
* pin A2
* pin B1
* pin A1
* pin Y
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o21ai_4 1 2 3 5 6 7 8 10
* net 1 VGND
* net 2 A2
* net 3 B1
* net 5 A1
* net 6 Y
* net 7 VPWR
* net 8 VPB
* device instance $1 r0 *1 0.5,1.985 pfet_01v8_hvt
M$1 9 5 7 8 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=580000000000P PS=6370000U PD=5160000U
* device instance $4 r0 *1 1.79,1.985 pfet_01v8_hvt
M$4 6 2 9 8 pfet_01v8_hvt L=150000U W=4000000U AS=560000000000P
+ AD=560000000000P PS=5120000U PD=5120000U
* device instance $9 r0 *1 3.98,1.985 pfet_01v8_hvt
M$9 6 3 7 8 pfet_01v8_hvt L=150000U W=4000000U AS=580000000000P
+ AD=685000000000P PS=5160000U PD=6370000U
* device instance $13 r0 *1 0.5,0.56 nfet_01v8
M$13 1 5 4 10 nfet_01v8 L=150000U W=2600000U AS=458250000000P AD=364000000000P
+ PS=4660000U PD=3720000U
* device instance $16 r0 *1 1.79,0.56 nfet_01v8
M$16 4 2 1 10 nfet_01v8 L=150000U W=2600000U AS=364000000000P AD=377000000000P
+ PS=3720000U PD=3760000U
* device instance $21 r0 *1 3.98,0.56 nfet_01v8
M$21 6 3 4 10 nfet_01v8 L=150000U W=2600000U AS=364000000000P AD=458250000000P
+ PS=3720000U PD=4660000U
.ENDS sky130_fd_sc_hd__o21ai_4

* cell sky130_fd_sc_hd__a211oi_4
* pin VGND
* pin A2
* pin A1
* pin Y
* pin B1
* pin C1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a211oi_4 1 2 4 5 6 7 8 9 14
* net 1 VGND
* net 2 A2
* net 4 A1
* net 5 Y
* net 6 B1
* net 7 C1
* net 8 VPWR
* net 9 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 2 10 9 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $4 r0 *1 1.73,1.985 pfet_01v8_hvt
M$4 10 4 8 9 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $9 r0 *1 3.83,1.985 pfet_01v8_hvt
M$9 11 6 10 9 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $11 r0 *1 4.67,1.985 pfet_01v8_hvt
M$11 13 6 10 9 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=150000000000P PS=1270000U PD=1300000U
* device instance $12 r0 *1 5.12,1.985 pfet_01v8_hvt
M$12 5 7 13 9 pfet_01v8_hvt L=150000U W=1000000U AS=150000000000P
+ AD=140000000000P PS=1300000U PD=1280000U
* device instance $13 r0 *1 5.55,1.985 pfet_01v8_hvt
M$13 11 7 5 9 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=290000000000P PS=2560000U PD=2580000U
* device instance $15 r0 *1 6.43,1.985 pfet_01v8_hvt
M$15 12 7 5 9 pfet_01v8_hvt L=150000U W=1000000U AS=150000000000P
+ AD=155000000000P PS=1300000U PD=1310000U
* device instance $16 r0 *1 6.89,1.985 pfet_01v8_hvt
M$16 10 6 12 9 pfet_01v8_hvt L=150000U W=1000000U AS=155000000000P
+ AD=260000000000P PS=1310000U PD=2520000U
* device instance $17 r0 *1 0.47,0.56 nfet_01v8
M$17 3 2 1 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $20 r0 *1 1.73,0.56 nfet_01v8
M$20 5 4 3 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $25 r0 *1 3.83,0.56 nfet_01v8
M$25 5 6 1 14 nfet_01v8 L=150000U W=2600000U AS=378625000000P AD=477750000000P
+ PS=3765000U PD=4720000U
* device instance $28 r0 *1 5.17,0.56 nfet_01v8
M$28 1 7 5 14 nfet_01v8 L=150000U W=2600000U AS=352625000000P AD=354250000000P
+ PS=3685000U PD=3690000U
.ENDS sky130_fd_sc_hd__a211oi_4

* cell sky130_fd_sc_hd__nand4_4
* pin VGND
* pin D
* pin A
* pin C
* pin B
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand4_4 1 2 3 5 7 9 10 11 12
* net 1 VGND
* net 2 D
* net 3 A
* net 5 C
* net 7 B
* net 9 VPWR
* net 10 Y
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 2 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 10 5 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=800000000000P PS=5080000U PD=5600000U
* device instance $9 r0 *1 4.35,1.985 pfet_01v8_hvt
M$9 10 7 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=800000000000P
+ AD=570000000000P PS=5600000U PD=5140000U
* device instance $13 r0 *1 6.09,1.985 pfet_01v8_hvt
M$13 10 3 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=570000000000P
+ AD=665000000000P PS=5140000U PD=6330000U
* device instance $17 r0 *1 4.35,0.56 nfet_01v8
M$17 6 7 8 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=370500000000P
+ PS=4580000U PD=3740000U
* device instance $21 r0 *1 6.09,0.56 nfet_01v8
M$21 10 3 8 12 nfet_01v8 L=150000U W=2600000U AS=370500000000P AD=432250000000P
+ PS=3740000U PD=4580000U
* device instance $25 r0 *1 0.47,0.56 nfet_01v8
M$25 1 2 4 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $29 r0 *1 2.15,0.56 nfet_01v8
M$29 6 5 4 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nand4_4

* cell sky130_fd_sc_hd__nor2_2
* pin VGND
* pin 
* pin Y
* pin VPB
* pin A
* pin B
* pin VPWR
.SUBCKT sky130_fd_sc_hd__nor2_2 1 2 3 4 5 6 8
* net 1 VGND
* net 3 Y
* net 4 VPB
* net 5 A
* net 6 B
* net 8 VPWR
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 8 5 7 4 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=270000000000P PS=3830000U PD=2540000U
* device instance $3 r0 *1 1.33,1.985 pfet_01v8_hvt
M$3 3 6 7 4 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 0.49,0.56 nfet_01v8
M$5 3 5 1 2 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $7 r0 *1 1.33,0.56 nfet_01v8
M$7 3 6 1 2 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nor2_2

* cell sky130_fd_sc_hd__nand2_4
* pin VGND
* pin B
* pin Y
* pin A
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand2_4 1 3 4 5 6 7 8
* net 1 VGND
* net 3 B
* net 4 Y
* net 5 A
* net 6 VPWR
* net 7 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 4 3 6 7 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 4 5 6 7 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $9 r0 *1 0.47,0.56 nfet_01v8
M$9 1 3 2 8 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $13 r0 *1 2.15,0.56 nfet_01v8
M$13 4 5 2 8 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__nand2_4

* cell sky130_fd_sc_hd__xnor2_4
* pin VGND
* pin B
* pin A
* pin Y
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__xnor2_4 1 2 3 7 8 10 11
* net 1 VGND
* net 2 B
* net 3 A
* net 7 Y
* net 8 VPWR
* net 10 VPB
* device instance $1 r0 *1 8.335,1.985 pfet_01v8_hvt
M$1 8 5 7 10 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=685000000000P PS=6370000U PD=6370000U
* device instance $5 r0 *1 0.545,1.985 pfet_01v8_hvt
M$5 8 2 5 10 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $9 r0 *1 2.225,1.985 pfet_01v8_hvt
M$9 8 3 5 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $13 r0 *1 4.435,1.985 pfet_01v8_hvt
M$13 8 3 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $17 r0 *1 6.115,1.985 pfet_01v8_hvt
M$17 7 2 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 8.335,0.56 nfet_01v8
M$21 7 5 6 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=445250000000P
+ PS=4580000U PD=4620000U
* device instance $25 r0 *1 4.435,0.56 nfet_01v8
M$25 6 3 1 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $29 r0 *1 6.115,0.56 nfet_01v8
M$29 6 2 1 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $33 r0 *1 0.545,0.56 nfet_01v8
M$33 5 2 4 11 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=351000000000P
+ PS=4620000U PD=3680000U
* device instance $37 r0 *1 2.225,0.56 nfet_01v8
M$37 1 3 4 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__xnor2_4

* cell sky130_fd_sc_hd__nand2_2
* pin VGND
* pin 
* pin B
* pin Y
* pin A
* pin VPB
* pin VPWR
.SUBCKT sky130_fd_sc_hd__nand2_2 1 2 4 5 6 7 8
* net 1 VGND
* net 4 B
* net 5 Y
* net 6 A
* net 7 VPB
* net 8 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 5 4 8 7 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 5 6 8 7 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 1 4 3 2 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $7 r0 *1 1.31,0.56 nfet_01v8
M$7 5 6 3 2 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__nand2_2

* cell sky130_fd_sc_hd__xor2_4
* pin VGND
* pin A
* pin B
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__xor2_4 1 2 3 6 8 10 11
* net 1 VGND
* net 2 A
* net 3 B
* net 6 X
* net 8 VPWR
* net 10 VPB
* device instance $1 r0 *1 8.255,1.985 pfet_01v8_hvt
M$1 9 4 6 10 pfet_01v8_hvt L=150000U W=4000000U AS=677450000000P
+ AD=685000000000P PS=6370000U PD=6370000U
* device instance $5 r0 *1 4.365,1.985 pfet_01v8_hvt
M$5 8 3 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $9 r0 *1 6.045,1.985 pfet_01v8_hvt
M$9 8 2 9 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=661800000000P PS=5080000U PD=6330000U
* device instance $13 r0 *1 0.485,1.985 pfet_01v8_hvt
M$13 8 2 7 10 pfet_01v8_hvt L=150000U W=4000000U AS=680000000000P
+ AD=540000000000P PS=6360000U PD=5080000U
* device instance $17 r0 *1 2.165,1.985 pfet_01v8_hvt
M$17 4 3 7 10 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $21 r0 *1 8.255,0.56 nfet_01v8
M$21 6 4 1 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=445250000000P
+ PS=4580000U PD=4620000U
* device instance $25 r0 *1 4.365,0.56 nfet_01v8
M$25 6 3 5 11 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $29 r0 *1 6.045,0.56 nfet_01v8
M$29 1 2 5 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
* device instance $33 r0 *1 0.485,0.56 nfet_01v8
M$33 4 2 1 11 nfet_01v8 L=150000U W=2600000U AS=442000000000P AD=351000000000P
+ PS=4610000U PD=3680000U
* device instance $37 r0 *1 2.165,0.56 nfet_01v8
M$37 4 3 1 11 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__xor2_4

* cell sky130_fd_sc_hd__buf_4
* pin VPB
* pin A
* pin VPWR
* pin VGND
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__buf_4 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 VPWR
* net 5 VGND
* net 6 X
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 4 3 2 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 6 2 4 1 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $6 r0 *1 0.47,0.56 nfet_01v8
M$6 5 3 2 7 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 0.89,0.56 nfet_01v8
M$7 6 2 5 7 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__buf_4

* cell sky130_fd_sc_hd__and2_0
* pin VPB
* pin A
* pin B
* pin X
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__and2_0 1 2 3 5 6 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 5 X
* net 6 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.54,2.275 pfet_01v8_hvt
M$1 4 2 6 1 pfet_01v8_hvt L=150000U W=420000U AS=111300000000P AD=60900000000P
+ PS=1370000U PD=710000U
* device instance $2 r0 *1 0.98,2.275 pfet_01v8_hvt
M$2 4 3 6 1 pfet_01v8_hvt L=150000U W=420000U AS=184100000000P AD=60900000000P
+ PS=1260000U PD=710000U
* device instance $3 r0 *1 1.75,2.165 pfet_01v8_hvt
M$3 5 4 6 1 pfet_01v8_hvt L=150000U W=640000U AS=184100000000P AD=169600000000P
+ PS=1260000U PD=1810000U
* device instance $4 r0 *1 0.54,0.445 nfet_01v8
M$4 9 2 4 8 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=44100000000P
+ PS=1370000U PD=630000U
* device instance $5 r0 *1 0.9,0.445 nfet_01v8
M$5 7 3 9 8 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=96600000000P
+ PS=630000U PD=880000U
* device instance $6 r0 *1 1.51,0.445 nfet_01v8
M$6 5 4 7 8 nfet_01v8 L=150000U W=420000U AS=96600000000P AD=111300000000P
+ PS=880000U PD=1370000U
.ENDS sky130_fd_sc_hd__and2_0

* cell sky130_fd_sc_hd__nand4_2
* pin VGND
* pin D
* pin C
* pin B
* pin A
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__nand4_2 1 5 6 7 8 9 10 11 12
* net 1 VGND
* net 5 D
* net 6 C
* net 7 B
* net 8 A
* net 9 VPWR
* net 10 Y
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 5 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 10 6 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=350000000000P PS=2540000U PD=2700000U
* device instance $5 r0 *1 2.31,1.985 pfet_01v8_hvt
M$5 10 7 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=350000000000P
+ AD=470000000000P PS=2700000U PD=2940000U
* device instance $7 r0 *1 3.55,1.985 pfet_01v8_hvt
M$7 10 8 9 11 pfet_01v8_hvt L=150000U W=2000000U AS=470000000000P
+ AD=555000000000P PS=2940000U PD=4110000U
* device instance $9 r0 *1 2.71,0.56 nfet_01v8
M$9 3 7 4 12 nfet_01v8 L=150000U W=1300000U AS=269750000000P AD=175500000000P
+ PS=2780000U PD=1840000U
* device instance $11 r0 *1 3.55,0.56 nfet_01v8
M$11 10 8 4 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=321750000000P
+ PS=1840000U PD=2940000U
* device instance $13 r0 *1 0.47,0.56 nfet_01v8
M$13 1 5 2 12 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $15 r0 *1 1.31,0.56 nfet_01v8
M$15 3 6 2 12 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
.ENDS sky130_fd_sc_hd__nand4_2

* cell sky130_fd_sc_hd__and3_1
* pin VGND
* pin B
* pin X
* pin A
* pin C
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__and3_1 1 2 3 6 7 9 10 11
* net 1 VGND
* net 2 B
* net 3 X
* net 6 A
* net 7 C
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.47,1.71 pfet_01v8_hvt
M$1 9 6 8 10 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $2 r0 *1 0.89,1.71 pfet_01v8_hvt
M$2 8 2 9 10 pfet_01v8_hvt L=150000U W=420000U AS=56700000000P AD=66150000000P
+ PS=690000U PD=735000U
* device instance $3 r0 *1 1.355,1.71 pfet_01v8_hvt
M$3 8 7 9 10 pfet_01v8_hvt L=150000U W=420000U AS=142225000000P AD=66150000000P
+ PS=1335000U PD=735000U
* device instance $4 r0 *1 1.83,1.985 pfet_01v8_hvt
M$4 3 8 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=142225000000P
+ AD=260000000000P PS=1335000U PD=2520000U
* device instance $5 r0 *1 0.47,0.445 nfet_01v8
M$5 5 6 8 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $6 r0 *1 0.83,0.445 nfet_01v8
M$6 4 2 5 11 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=44100000000P
+ PS=630000U PD=630000U
* device instance $7 r0 *1 1.19,0.445 nfet_01v8
M$7 1 7 4 11 nfet_01v8 L=150000U W=420000U AS=44100000000P AD=131650000000P
+ PS=630000U PD=1140000U
* device instance $8 r0 *1 1.83,0.56 nfet_01v8
M$8 3 8 1 11 nfet_01v8 L=150000U W=650000U AS=131650000000P AD=169000000000P
+ PS=1140000U PD=1820000U
.ENDS sky130_fd_sc_hd__and3_1

* cell sky130_fd_sc_hd__o21ai_1
* pin VPB
* pin A1
* pin B1
* pin A2
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__o21ai_1 1 2 3 4 5 7 8 9
* net 1 VPB
* net 2 A1
* net 3 B1
* net 4 A2
* net 5 VPWR
* net 7 VGND
* net 8 Y
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=105000000000P PS=2520000U PD=1210000U
* device instance $2 r0 *1 0.83,1.985 pfet_01v8_hvt
M$2 8 4 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=174000000000P PS=1210000U PD=1390000U
* device instance $3 r0 *1 1.37,2.135 pfet_01v8_hvt
M$3 5 3 8 1 pfet_01v8_hvt L=150000U W=700000U AS=174000000000P AD=182000000000P
+ PS=1390000U PD=1920000U
* device instance $4 r0 *1 0.47,0.56 nfet_01v8
M$4 7 2 6 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=107250000000P
+ PS=1820000U PD=980000U
* device instance $5 r0 *1 0.95,0.56 nfet_01v8
M$5 6 4 7 9 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=87750000000P
+ PS=980000U PD=920000U
* device instance $6 r0 *1 1.37,0.56 nfet_01v8
M$6 8 3 6 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o21ai_1

* cell sky130_fd_sc_hd__or2_1
* pin VPB
* pin B
* pin A
* pin X
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__or2_1 1 2 3 4 5 7 8
* net 1 VPB
* net 2 B
* net 3 A
* net 4 X
* net 5 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.675,1.695 pfet_01v8_hvt
M$1 9 2 6 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=44100000000P
+ PS=1360000U PD=630000U
* device instance $2 r0 *1 1.035,1.695 pfet_01v8_hvt
M$2 7 3 9 1 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P AD=145750000000P
+ PS=630000U PD=1335000U
* device instance $3 r0 *1 1.52,1.985 pfet_01v8_hvt
M$3 4 6 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=145750000000P
+ AD=340000000000P PS=1335000U PD=2680000U
* device instance $4 r0 *1 0.615,0.445 nfet_01v8
M$4 6 2 5 8 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=56700000000P
+ PS=1360000U PD=690000U
* device instance $5 r0 *1 1.035,0.445 nfet_01v8
M$5 5 3 6 8 nfet_01v8 L=150000U W=420000U AS=56700000000P AD=100250000000P
+ PS=690000U PD=985000U
* device instance $6 r0 *1 1.52,0.56 nfet_01v8
M$6 4 6 5 8 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=169000000000P
+ PS=985000U PD=1820000U
.ENDS sky130_fd_sc_hd__or2_1

* cell sky130_fd_sc_hd__xor2_1
* pin VPB
* pin B
* pin A
* pin VPWR
* pin X
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__xor2_1 1 2 3 6 7 8 9
* net 1 VPB
* net 2 B
* net 3 A
* net 6 VPWR
* net 7 X
* net 8 VGND
* device instance $1 r0 *1 2.71,1.985 pfet_01v8_hvt
M$1 7 4 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=300000000000P PS=2520000U PD=2600000U
* device instance $2 r0 *1 0.51,1.985 pfet_01v8_hvt
M$2 10 2 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $3 r0 *1 0.93,1.985 pfet_01v8_hvt
M$3 6 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $4 r0 *1 1.35,1.985 pfet_01v8_hvt
M$4 5 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $5 r0 *1 1.77,1.985 pfet_01v8_hvt
M$5 6 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $6 r0 *1 0.51,0.56 nfet_01v8
M$6 4 2 8 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 0.93,0.56 nfet_01v8
M$7 8 3 4 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $8 r0 *1 1.35,0.56 nfet_01v8
M$8 11 3 8 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $9 r0 *1 1.77,0.56 nfet_01v8
M$9 7 2 11 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=250250000000P
+ PS=920000U PD=1420000U
* device instance $10 r0 *1 2.69,0.56 nfet_01v8
M$10 8 4 7 9 nfet_01v8 L=150000U W=650000U AS=250250000000P AD=208000000000P
+ PS=1420000U PD=1940000U
.ENDS sky130_fd_sc_hd__xor2_1

* cell sky130_fd_sc_hd__buf_2
* pin VPB
* pin A
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__buf_2 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 VGND
* net 5 X
* net 6 VPWR
* device instance $1 r0 *1 0.47,2.125 pfet_01v8_hvt
M$1 2 3 6 1 pfet_01v8_hvt L=150000U W=640000U AS=149000000000P AD=166400000000P
+ PS=1325000U PD=1800000U
* device instance $2 r0 *1 0.945,1.985 pfet_01v8_hvt
M$2 5 2 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=284000000000P
+ AD=400000000000P PS=2595000U PD=3800000U
* device instance $4 r0 *1 0.47,0.445 nfet_01v8
M$4 4 3 2 7 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=97000000000P
+ PS=1360000U PD=975000U
* device instance $5 r0 *1 0.945,0.56 nfet_01v8
M$5 5 2 4 7 nfet_01v8 L=150000U W=1300000U AS=184750000000P AD=260000000000P
+ PS=1895000U PD=2750000U
.ENDS sky130_fd_sc_hd__buf_2

* cell sky130_fd_sc_hd__inv_1
* pin VPB
* pin A
* pin VPWR
* pin VGND
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__inv_1 1 2 3 4 5 6
* net 1 VPB
* net 2 A
* net 3 VPWR
* net 4 VGND
* net 5 Y
* device instance $1 r0 *1 0.675,1.985 pfet_01v8_hvt
M$1 5 2 3 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $2 r0 *1 0.675,0.56 nfet_01v8
M$2 5 2 4 6 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=169000000000P
+ PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__inv_1

* cell sky130_fd_sc_hd__a31o_1
* pin VGND
* pin X
* pin A3
* pin A2
* pin A1
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a31o_1 1 2 6 7 8 9 11 12 13
* net 1 VGND
* net 2 X
* net 6 A3
* net 7 A2
* net 8 A1
* net 9 B1
* net 11 VPWR
* net 12 VPB
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 11 3 2 12 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=172500000000P PS=2530000U PD=1345000U
* device instance $2 r0 *1 0.97,1.985 pfet_01v8_hvt
M$2 10 6 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=172500000000P
+ AD=160000000000P PS=1345000U PD=1320000U
* device instance $3 r0 *1 1.44,1.985 pfet_01v8_hvt
M$3 11 7 10 12 pfet_01v8_hvt L=150000U W=1000000U AS=160000000000P
+ AD=165000000000P PS=1320000U PD=1330000U
* device instance $4 r0 *1 1.92,1.985 pfet_01v8_hvt
M$4 10 8 11 12 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=165000000000P PS=1330000U PD=1330000U
* device instance $5 r0 *1 2.4,1.985 pfet_01v8_hvt
M$5 3 9 10 12 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=320000000000P PS=1330000U PD=2640000U
* device instance $6 r0 *1 0.475,0.56 nfet_01v8
M$6 1 3 2 13 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=112125000000P
+ PS=1830000U PD=995000U
* device instance $7 r0 *1 0.97,0.56 nfet_01v8
M$7 4 6 1 13 nfet_01v8 L=150000U W=650000U AS=112125000000P AD=104000000000P
+ PS=995000U PD=970000U
* device instance $8 r0 *1 1.44,0.56 nfet_01v8
M$8 5 7 4 13 nfet_01v8 L=150000U W=650000U AS=104000000000P AD=107250000000P
+ PS=970000U PD=980000U
* device instance $9 r0 *1 1.92,0.56 nfet_01v8
M$9 3 8 5 13 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=107250000000P
+ PS=980000U PD=980000U
* device instance $10 r0 *1 2.4,0.56 nfet_01v8
M$10 1 9 3 13 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=208000000000P
+ PS=980000U PD=1940000U
.ENDS sky130_fd_sc_hd__a31o_1

* cell sky130_fd_sc_hd__a21oi_1
* pin VPB
* pin B1
* pin A1
* pin A2
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__a21oi_1 1 2 3 4 5 7 8 9
* net 1 VPB
* net 2 B1
* net 3 A1
* net 4 A2
* net 5 VGND
* net 7 VPWR
* net 8 Y
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 6 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=140000000000P PS=2530000U PD=1280000U
* device instance $2 r0 *1 0.92,1.985 pfet_01v8_hvt
M$2 7 3 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=147500000000P PS=1280000U PD=1295000U
* device instance $3 r0 *1 1.365,1.985 pfet_01v8_hvt
M$3 6 4 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=147500000000P
+ AD=265000000000P PS=1295000U PD=2530000U
* device instance $4 r0 *1 0.49,0.56 nfet_01v8
M$4 8 2 5 9 nfet_01v8 L=150000U W=650000U AS=172250000000P AD=91000000000P
+ PS=1830000U PD=930000U
* device instance $5 r0 *1 0.92,0.56 nfet_01v8
M$5 10 3 8 9 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=95875000000P
+ PS=930000U PD=945000U
* device instance $6 r0 *1 1.365,0.56 nfet_01v8
M$6 5 4 10 9 nfet_01v8 L=150000U W=650000U AS=95875000000P AD=172250000000P
+ PS=945000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21oi_1

* cell sky130_fd_sc_hd__o21ai_0
* pin VPB
* pin A1
* pin A2
* pin B1
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__o21ai_0 1 2 3 4 5 6 8 9
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 B1
* net 5 VPWR
* net 6 Y
* net 8 VGND
* device instance $1 r0 *1 0.525,2.165 pfet_01v8_hvt
M$1 10 2 5 1 pfet_01v8_hvt L=150000U W=640000U AS=169600000000P AD=76800000000P
+ PS=1810000U PD=880000U
* device instance $2 r0 *1 0.915,2.165 pfet_01v8_hvt
M$2 6 3 10 1 pfet_01v8_hvt L=150000U W=640000U AS=76800000000P AD=89600000000P
+ PS=880000U PD=920000U
* device instance $3 r0 *1 1.345,2.165 pfet_01v8_hvt
M$3 5 4 6 1 pfet_01v8_hvt L=150000U W=640000U AS=89600000000P AD=182400000000P
+ PS=920000U PD=1850000U
* device instance $4 r0 *1 0.5,0.445 nfet_01v8
M$4 8 2 7 9 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=58800000000P
+ PS=1370000U PD=700000U
* device instance $5 r0 *1 0.93,0.445 nfet_01v8
M$5 7 3 8 9 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=58800000000P
+ PS=700000U PD=700000U
* device instance $6 r0 *1 1.36,0.445 nfet_01v8
M$6 6 4 7 9 nfet_01v8 L=150000U W=420000U AS=58800000000P AD=111300000000P
+ PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__o21ai_0

* cell sky130_fd_sc_hd__nand4_1
* pin VPB
* pin C
* pin A
* pin B
* pin D
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__nand4_1 1 2 3 4 5 6 7 8 9
* net 1 VPB
* net 2 C
* net 3 A
* net 4 B
* net 5 D
* net 6 VPWR
* net 7 Y
* net 8 VGND
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 7 5 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 6 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 7 4 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $4 r0 *1 1.79,1.985 pfet_01v8_hvt
M$4 6 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=300000000000P PS=1330000U PD=2600000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 12 5 8 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $6 r0 *1 0.89,0.56 nfet_01v8
M$6 11 2 12 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $7 r0 *1 1.31,0.56 nfet_01v8
M$7 10 4 11 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $8 r0 *1 1.79,0.56 nfet_01v8
M$8 7 3 10 9 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=195000000000P
+ PS=980000U PD=1900000U
.ENDS sky130_fd_sc_hd__nand4_1

* cell sky130_fd_sc_hd__nor3_1
* pin VPB
* pin A
* pin B
* pin C
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor3_1 1 2 3 4 5 6 7 8
* net 1 VPB
* net 2 A
* net 3 B
* net 4 C
* net 5 Y
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 4 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 9 3 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=135000000000P PS=1270000U PD=1270000U
* device instance $3 r0 *1 1.31,1.985 pfet_01v8_hvt
M$3 7 2 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $4 r0 *1 0.47,0.56 nfet_01v8
M$4 6 4 5 8 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $5 r0 *1 0.89,0.56 nfet_01v8
M$5 5 3 6 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=87750000000P
+ PS=920000U PD=920000U
* device instance $6 r0 *1 1.31,0.56 nfet_01v8
M$6 6 2 5 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor3_1

* cell sky130_fd_sc_hd__clkbuf_4
* pin VPB
* pin A
* pin VGND
* pin X
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__clkbuf_4 1 3 4 5 6 7
* net 1 VPB
* net 3 A
* net 4 VGND
* net 5 X
* net 6 VPWR
* device instance $1 r0 *1 0.475,1.985 pfet_01v8_hvt
M$1 6 3 2 1 pfet_01v8_hvt L=150000U W=1000000U AS=265000000000P
+ AD=165000000000P PS=2530000U PD=1330000U
* device instance $2 r0 *1 0.955,1.985 pfet_01v8_hvt
M$2 5 2 6 1 pfet_01v8_hvt L=150000U W=4000000U AS=585000000000P
+ AD=720000000000P PS=5170000U PD=6440000U
* device instance $6 r0 *1 0.475,0.445 nfet_01v8
M$6 4 3 2 7 nfet_01v8 L=150000U W=420000U AS=111300000000P AD=70350000000P
+ PS=1370000U PD=755000U
* device instance $7 r0 *1 0.96,0.445 nfet_01v8
M$7 5 2 4 7 nfet_01v8 L=150000U W=1680000U AS=246750000000P AD=298200000000P
+ PS=2855000U PD=3520000U
.ENDS sky130_fd_sc_hd__clkbuf_4

* cell sky130_fd_sc_hd__buf_16
* pin VGND
* pin A
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__buf_16 1 2 4 5 6 7
* net 1 VGND
* net 2 A
* net 4 X
* net 5 VPWR
* net 6 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 3 2 5 6 pfet_01v8_hvt L=150000U W=6000000U AS=935000000000P
+ AD=810000000000P PS=8870000U PD=7620000U
* device instance $7 r0 *1 2.99,1.985 pfet_01v8_hvt
M$7 4 3 5 6 pfet_01v8_hvt L=150000U W=16000000U AS=2.16e+12P AD=2.285e+12P
+ PS=20320000U PD=21570000U
* device instance $23 r0 *1 0.47,0.56 nfet_01v8
M$23 3 2 1 7 nfet_01v8 L=150000U W=3900000U AS=607750000000P AD=526500000000P
+ PS=6420000U PD=5520000U
* device instance $29 r0 *1 2.99,0.56 nfet_01v8
M$29 4 3 1 7 nfet_01v8 L=150000U W=10400000U AS=1.404e+12P AD=1.48525e+12P
+ PS=14720000U PD=15620000U
.ENDS sky130_fd_sc_hd__buf_16

* cell sky130_fd_sc_hd__nor4b_1
* pin VPB
* pin C
* pin B
* pin A
* pin D_N
* pin VGND
* pin Y
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor4b_1 1 2 3 4 5 6 7 8 10
* net 1 VPB
* net 2 C
* net 3 B
* net 4 A
* net 5 D_N
* net 6 VGND
* net 7 Y
* net 8 VPWR
* device instance $1 r0 *1 2.535,1.89 pfet_01v8_hvt
M$1 9 5 8 1 pfet_01v8_hvt L=150000U W=420000U AS=145750000000P AD=109200000000P
+ PS=1335000U PD=1360000U
* device instance $2 r0 *1 0.73,1.985 pfet_01v8_hvt
M$2 13 9 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=520000000000P
+ AD=135000000000P PS=3040000U PD=1270000U
* device instance $3 r0 *1 1.15,1.985 pfet_01v8_hvt
M$3 12 2 13 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $4 r0 *1 1.63,1.985 pfet_01v8_hvt
M$4 11 3 12 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=135000000000P PS=1330000U PD=1270000U
* device instance $5 r0 *1 2.05,1.985 pfet_01v8_hvt
M$5 8 4 11 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=145750000000P PS=1270000U PD=1335000U
* device instance $6 r0 *1 0.73,0.56 nfet_01v8
M$6 7 9 6 10 nfet_01v8 L=150000U W=650000U AS=182000000000P AD=87750000000P
+ PS=1860000U PD=920000U
* device instance $7 r0 *1 1.15,0.56 nfet_01v8
M$7 6 2 7 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $8 r0 *1 1.63,0.56 nfet_01v8
M$8 7 3 6 10 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=87750000000P
+ PS=980000U PD=920000U
* device instance $9 r0 *1 2.05,0.56 nfet_01v8
M$9 6 4 7 10 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=100250000000P
+ PS=920000U PD=985000U
* device instance $10 r0 *1 2.535,0.675 nfet_01v8
M$10 9 5 6 10 nfet_01v8 L=150000U W=420000U AS=100250000000P AD=109200000000P
+ PS=985000U PD=1360000U
.ENDS sky130_fd_sc_hd__nor4b_1

* cell sky130_fd_sc_hd__o21bai_2
* pin VGND
* pin Y
* pin B1_N
* pin A2
* pin A1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o21bai_2 1 4 5 6 7 8 10 11
* net 1 VGND
* net 4 Y
* net 5 B1_N
* net 6 A2
* net 7 A1
* net 8 VPWR
* net 10 VPB
* device instance $1 r0 *1 2.32,1.985 pfet_01v8_hvt
M$1 4 6 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $3 r0 *1 3.16,1.985 pfet_01v8_hvt
M$3 8 7 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=415000000000P PS=2540000U PD=3830000U
* device instance $5 r0 *1 0.475,1.695 pfet_01v8_hvt
M$5 8 5 2 10 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P
+ AD=145750000000P PS=1360000U PD=1335000U
* device instance $6 r0 *1 0.96,1.985 pfet_01v8_hvt
M$6 4 2 8 10 pfet_01v8_hvt L=150000U W=2000000U AS=280750000000P
+ AD=395000000000P PS=2605000U PD=3790000U
* device instance $8 r0 *1 1.48,0.56 nfet_01v8
M$8 4 2 3 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $10 r0 *1 2.32,0.56 nfet_01v8
M$10 1 6 3 11 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $12 r0 *1 3.16,0.56 nfet_01v8
M$12 1 7 3 11 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=269750000000P
+ PS=1840000U PD=2780000U
* device instance $14 r0 *1 0.475,0.675 nfet_01v8
M$14 2 5 1 11 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=109200000000P
+ PS=1360000U PD=1360000U
.ENDS sky130_fd_sc_hd__o21bai_2

* cell sky130_fd_sc_hd__mux2i_2
* pin VGND
* pin S
* pin A0
* pin A1
* pin VPWR
* pin Y
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2i_2 1 2 6 7 8 11 12 13
* net 1 VGND
* net 2 S
* net 6 A0
* net 7 A1
* net 8 VPWR
* net 11 Y
* net 12 VPB
* device instance $1 r0 *1 3.09,1.985 pfet_01v8_hvt
M$1 9 6 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=290000000000P PS=3790000U PD=2580000U
* device instance $3 r0 *1 3.97,1.985 pfet_01v8_hvt
M$3 10 7 11 12 pfet_01v8_hvt L=150000U W=2000000U AS=292500000000P
+ AD=592500000000P PS=2585000U PD=4185000U
* device instance $5 r0 *1 0.47,1.985 pfet_01v8_hvt
M$5 8 2 3 12 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $6 r0 *1 0.89,1.985 pfet_01v8_hvt
M$6 9 2 8 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=270000000000P PS=2540000U PD=2540000U
* device instance $8 r0 *1 1.73,1.985 pfet_01v8_hvt
M$8 10 3 8 12 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $10 r0 *1 3.09,0.56 nfet_01v8
M$10 5 6 11 13 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=188500000000P
+ PS=2740000U PD=1880000U
* device instance $12 r0 *1 3.97,0.56 nfet_01v8
M$12 4 7 11 13 nfet_01v8 L=150000U W=1300000U AS=190125000000P AD=385125000000P
+ PS=1885000U PD=3135000U
* device instance $14 r0 *1 0.47,0.56 nfet_01v8
M$14 1 2 3 13 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $15 r0 *1 0.89,0.56 nfet_01v8
M$15 4 2 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=175500000000P
+ PS=1840000U PD=1840000U
* device instance $17 r0 *1 1.73,0.56 nfet_01v8
M$17 5 3 1 13 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__mux2i_2

* cell sky130_fd_sc_hd__mux2_1
* pin VGND
* pin X
* pin A1
* pin A0
* pin S
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__mux2_1 1 2 3 5 9 10 11 14
* net 1 VGND
* net 2 X
* net 3 A1
* net 5 A0
* net 9 S
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 1.015,2.08 pfet_01v8_hvt
M$1 12 9 10 11 pfet_01v8_hvt L=150000U W=420000U AS=158350000000P
+ AD=76650000000P PS=1395000U PD=785000U
* device instance $2 r0 *1 1.53,2.08 pfet_01v8_hvt
M$2 4 5 12 11 pfet_01v8_hvt L=150000U W=420000U AS=76650000000P
+ AD=193200000000P PS=785000U PD=1340000U
* device instance $3 r0 *1 2.6,2.08 pfet_01v8_hvt
M$3 13 3 4 11 pfet_01v8_hvt L=150000U W=420000U AS=193200000000P
+ AD=44100000000P PS=1340000U PD=630000U
* device instance $4 r0 *1 2.96,2.08 pfet_01v8_hvt
M$4 10 6 13 11 pfet_01v8_hvt L=150000U W=420000U AS=44100000000P
+ AD=69300000000P PS=630000U PD=750000U
* device instance $5 r0 *1 3.44,2.08 pfet_01v8_hvt
M$5 6 9 10 11 pfet_01v8_hvt L=150000U W=420000U AS=69300000000P
+ AD=117600000000P PS=750000U PD=1400000U
* device instance $6 r0 *1 0.47,1.985 pfet_01v8_hvt
M$6 10 4 2 11 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=158350000000P PS=2520000U PD=1395000U
* device instance $7 r0 *1 1.015,0.445 nfet_01v8
M$7 7 9 1 14 nfet_01v8 L=150000U W=420000U AS=112850000000P AD=69300000000P
+ PS=1045000U PD=750000U
* device instance $8 r0 *1 1.495,0.445 nfet_01v8
M$8 4 3 7 14 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=99750000000P
+ PS=750000U PD=895000U
* device instance $9 r0 *1 2.12,0.445 nfet_01v8
M$9 8 5 4 14 nfet_01v8 L=150000U W=420000U AS=99750000000P AD=69300000000P
+ PS=895000U PD=750000U
* device instance $10 r0 *1 2.6,0.445 nfet_01v8
M$10 1 6 8 14 nfet_01v8 L=150000U W=420000U AS=69300000000P AD=144900000000P
+ PS=750000U PD=1110000U
* device instance $11 r0 *1 3.44,0.445 nfet_01v8
M$11 6 9 1 14 nfet_01v8 L=150000U W=420000U AS=144900000000P AD=109200000000P
+ PS=1110000U PD=1360000U
* device instance $12 r0 *1 0.47,0.56 nfet_01v8
M$12 1 4 2 14 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=112850000000P
+ PS=1820000U PD=1045000U
.ENDS sky130_fd_sc_hd__mux2_1

* cell sky130_fd_sc_hd__a31oi_1
* pin VPB
* pin A3
* pin A2
* pin A1
* pin B1
* pin VGND
* pin VPWR
* pin Y
* pin 
.SUBCKT sky130_fd_sc_hd__a31oi_1 1 2 3 4 5 6 8 9 10
* net 1 VPB
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 B1
* net 6 VGND
* net 8 VPWR
* net 9 Y
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 7 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.89,1.985 pfet_01v8_hvt
M$2 8 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=152500000000P PS=1270000U PD=1305000U
* device instance $3 r0 *1 1.345,1.985 pfet_01v8_hvt
M$3 7 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=152500000000P
+ AD=162500000000P PS=1305000U PD=1325000U
* device instance $4 r0 *1 1.82,1.985 pfet_01v8_hvt
M$4 9 5 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=162500000000P
+ AD=270000000000P PS=1325000U PD=2540000U
* device instance $5 r0 *1 0.47,0.56 nfet_01v8
M$5 12 2 6 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=68250000000P
+ PS=1820000U PD=860000U
* device instance $6 r0 *1 0.83,0.56 nfet_01v8
M$6 11 3 12 10 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=118625000000P
+ PS=860000U PD=1015000U
* device instance $7 r0 *1 1.345,0.56 nfet_01v8
M$7 9 4 11 10 nfet_01v8 L=150000U W=650000U AS=118625000000P AD=105625000000P
+ PS=1015000U PD=975000U
* device instance $8 r0 *1 1.82,0.56 nfet_01v8
M$8 6 5 9 10 nfet_01v8 L=150000U W=650000U AS=105625000000P AD=175500000000P
+ PS=975000U PD=1840000U
.ENDS sky130_fd_sc_hd__a31oi_1

* cell sky130_fd_sc_hd__xor2_2
* pin VGND
* pin A
* pin B
* pin X
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__xor2_2 1 3 4 6 8 10 11
* net 1 VGND
* net 3 A
* net 4 B
* net 6 X
* net 8 VPWR
* net 10 VPB
* device instance $1 r0 *1 4.94,1.985 pfet_01v8_hvt
M$1 6 2 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=415000000000P PS=3790000U PD=3830000U
* device instance $3 r0 *1 2.685,1.985 pfet_01v8_hvt
M$3 8 3 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=395000000000P
+ AD=270000000000P PS=3790000U PD=2540000U
* device instance $5 r0 *1 3.525,1.985 pfet_01v8_hvt
M$5 8 4 9 10 pfet_01v8_hvt L=150000U W=2000000U AS=297500000000P
+ AD=422500000000P PS=2595000U PD=3845000U
* device instance $7 r0 *1 0.485,1.985 pfet_01v8_hvt
M$7 8 3 7 10 pfet_01v8_hvt L=150000U W=2000000U AS=410000000000P
+ AD=270000000000P PS=3820000U PD=2540000U
* device instance $9 r0 *1 1.325,1.985 pfet_01v8_hvt
M$9 2 4 7 10 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=395000000000P PS=2540000U PD=3790000U
* device instance $11 r0 *1 4.94,0.56 nfet_01v8
M$11 6 2 1 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=256750000000P
+ PS=2740000U PD=2740000U
* device instance $13 r0 *1 2.685,0.56 nfet_01v8
M$13 1 3 5 11 nfet_01v8 L=150000U W=1300000U AS=256750000000P AD=175500000000P
+ PS=2740000U PD=1840000U
* device instance $15 r0 *1 3.525,0.56 nfet_01v8
M$15 6 4 5 11 nfet_01v8 L=150000U W=1300000U AS=193375000000P AD=274625000000P
+ PS=1895000U PD=2795000U
* device instance $17 r0 *1 0.485,0.56 nfet_01v8
M$17 2 3 1 11 nfet_01v8 L=150000U W=1300000U AS=266500000000P AD=175500000000P
+ PS=2770000U PD=1840000U
* device instance $19 r0 *1 1.325,0.56 nfet_01v8
M$19 2 4 1 11 nfet_01v8 L=150000U W=1300000U AS=175500000000P AD=256750000000P
+ PS=1840000U PD=2740000U
.ENDS sky130_fd_sc_hd__xor2_2

* cell sky130_fd_sc_hd__o31a_1
* pin VGND
* pin X
* pin A1
* pin A2
* pin A3
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o31a_1 1 2 5 6 7 8 9 10 13
* net 1 VGND
* net 2 X
* net 5 A1
* net 6 A2
* net 7 A3
* net 8 B1
* net 9 VPWR
* net 10 VPB
* device instance $1 r0 *1 0.65,1.985 pfet_01v8_hvt
M$1 9 4 2 10 pfet_01v8_hvt L=150000U W=1000000U AS=360000000000P
+ AD=195000000000P PS=2720000U PD=1390000U
* device instance $2 r0 *1 1.19,1.985 pfet_01v8_hvt
M$2 12 5 9 10 pfet_01v8_hvt L=150000U W=1000000U AS=195000000000P
+ AD=135000000000P PS=1390000U PD=1270000U
* device instance $3 r0 *1 1.61,1.985 pfet_01v8_hvt
M$3 11 6 12 10 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=165000000000P PS=1270000U PD=1330000U
* device instance $4 r0 *1 2.09,1.985 pfet_01v8_hvt
M$4 4 7 11 10 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=212500000000P PS=1330000U PD=1425000U
* device instance $5 r0 *1 2.665,1.985 pfet_01v8_hvt
M$5 9 8 4 10 pfet_01v8_hvt L=150000U W=1000000U AS=212500000000P
+ AD=345000000000P PS=1425000U PD=2690000U
* device instance $6 r0 *1 0.65,0.56 nfet_01v8
M$6 1 4 2 13 nfet_01v8 L=150000U W=650000U AS=234000000000P AD=126750000000P
+ PS=2020000U PD=1040000U
* device instance $7 r0 *1 1.19,0.56 nfet_01v8
M$7 3 5 1 13 nfet_01v8 L=150000U W=650000U AS=126750000000P AD=87750000000P
+ PS=1040000U PD=920000U
* device instance $8 r0 *1 1.61,0.56 nfet_01v8
M$8 1 6 3 13 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=107250000000P
+ PS=920000U PD=980000U
* device instance $9 r0 *1 2.09,0.56 nfet_01v8
M$9 3 7 1 13 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=107250000000P
+ PS=980000U PD=980000U
* device instance $10 r0 *1 2.57,0.56 nfet_01v8
M$10 4 8 3 13 nfet_01v8 L=150000U W=650000U AS=107250000000P AD=201500000000P
+ PS=980000U PD=1920000U
.ENDS sky130_fd_sc_hd__o31a_1

* cell sky130_fd_sc_hd__o31ai_4
* pin VGND
* pin B1
* pin Y
* pin A1
* pin A2
* pin A3
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o31ai_4 1 2 4 5 6 7 10 11 12
* net 1 VGND
* net 2 B1
* net 4 Y
* net 5 A1
* net 6 A2
* net 7 A3
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 4.385,1.985 pfet_01v8_hvt
M$1 9 7 4 11 pfet_01v8_hvt L=150000U W=4000000U AS=667800000000P
+ AD=540000000000P PS=6380000U PD=5080000U
* device instance $5 r0 *1 6.065,1.985 pfet_01v8_hvt
M$5 10 2 4 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665000000000P PS=5080000U PD=6330000U
* device instance $9 r0 *1 0.49,1.985 pfet_01v8_hvt
M$9 10 5 8 11 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=540000000000P PS=6370000U PD=5080000U
* device instance $13 r0 *1 2.17,1.985 pfet_01v8_hvt
M$13 9 6 8 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=665500000000P PS=5080000U PD=6370000U
* device instance $17 r0 *1 0.49,0.56 nfet_01v8
M$17 1 5 3 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $21 r0 *1 2.17,0.56 nfet_01v8
M$21 1 6 3 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $25 r0 *1 3.85,0.56 nfet_01v8
M$25 1 7 3 12 nfet_01v8 L=150000U W=2600000U AS=524875000000P AD=524875000000P
+ PS=4215000U PD=4215000U
* device instance $29 r0 *1 6.065,0.56 nfet_01v8
M$29 4 2 3 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__o31ai_4

* cell sky130_fd_sc_hd__o221ai_4
* pin VGND
* pin B2
* pin C1
* pin Y
* pin B1
* pin A1
* pin A2
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__o221ai_4 1 2 4 5 7 8 9 10 11 14
* net 1 VGND
* net 2 B2
* net 4 C1
* net 5 Y
* net 7 B1
* net 8 A1
* net 9 A2
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 5 4 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=685000000000P
+ AD=800000000000P PS=6370000U PD=5600000U
* device instance $5 r0 *1 2.69,1.985 pfet_01v8_hvt
M$5 12 7 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=800000000000P
+ AD=580000000000P PS=5600000U PD=5160000U
* device instance $8 r0 *1 3.95,1.985 pfet_01v8_hvt
M$8 5 2 12 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $13 r0 *1 6.13,1.985 pfet_01v8_hvt
M$13 13 8 10 11 pfet_01v8_hvt L=150000U W=4000000U AS=580000000000P
+ AD=700000000000P PS=5160000U PD=6400000U
* device instance $14 r0 *1 6.55,1.985 pfet_01v8_hvt
M$14 5 9 13 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=540000000000P PS=5080000U PD=5080000U
* device instance $21 r0 *1 2.69,0.56 nfet_01v8
M$21 3 7 6 14 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=377000000000P
+ PS=4580000U PD=3760000U
* device instance $24 r0 *1 3.95,0.56 nfet_01v8
M$24 6 2 3 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $29 r0 *1 6.13,0.56 nfet_01v8
M$29 1 8 6 14 nfet_01v8 L=150000U W=2600000U AS=377000000000P AD=432250000000P
+ PS=3760000U PD=4580000U
* device instance $30 r0 *1 6.55,0.56 nfet_01v8
M$30 6 9 1 14 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=351000000000P
+ PS=3680000U PD=3680000U
* device instance $37 r0 *1 0.49,0.56 nfet_01v8
M$37 5 4 3 14 nfet_01v8 L=150000U W=2600000U AS=445250000000P AD=432250000000P
+ PS=4620000U PD=4580000U
.ENDS sky130_fd_sc_hd__o221ai_4

* cell sky130_fd_sc_hd__a31oi_4
* pin VGND
* pin A3
* pin A2
* pin A1
* pin Y
* pin B1
* pin VPWR
* pin VPB
* pin 
.SUBCKT sky130_fd_sc_hd__a31oi_4 1 2 4 6 7 8 10 11 12
* net 1 VGND
* net 2 A3
* net 4 A2
* net 6 A1
* net 7 Y
* net 8 B1
* net 10 VPWR
* net 11 VPB
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 10 2 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=665000000000P
+ AD=540000000000P PS=6330000U PD=5080000U
* device instance $5 r0 *1 2.15,1.985 pfet_01v8_hvt
M$5 10 4 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=540000000000P
+ AD=550000000000P PS=5080000U PD=5100000U
* device instance $9 r0 *1 3.85,1.985 pfet_01v8_hvt
M$9 10 6 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=550000000000P
+ AD=790000000000P PS=5100000U PD=5580000U
* device instance $13 r0 *1 6.03,1.985 pfet_01v8_hvt
M$13 7 8 9 11 pfet_01v8_hvt L=150000U W=4000000U AS=790000000000P
+ AD=725000000000P PS=5580000U PD=6450000U
* device instance $17 r0 *1 4.35,0.56 nfet_01v8
M$17 5 6 7 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $21 r0 *1 6.03,0.56 nfet_01v8
M$21 1 8 7 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=471250000000P
+ PS=3680000U PD=4700000U
* device instance $25 r0 *1 0.47,0.56 nfet_01v8
M$25 1 2 3 12 nfet_01v8 L=150000U W=2600000U AS=432250000000P AD=351000000000P
+ PS=4580000U PD=3680000U
* device instance $29 r0 *1 2.15,0.56 nfet_01v8
M$29 5 4 3 12 nfet_01v8 L=150000U W=2600000U AS=351000000000P AD=432250000000P
+ PS=3680000U PD=4580000U
.ENDS sky130_fd_sc_hd__a31oi_4

* cell sky130_fd_sc_hd__a21oi_2
* pin VPB
* pin A1
* pin B1
* pin A2
* pin VPWR
* pin Y
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__a21oi_2 1 2 3 4 5 7 8 9
* net 1 VPB
* net 2 A1
* net 3 B1
* net 4 A2
* net 5 VPWR
* net 7 Y
* net 8 VGND
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 5 4 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=415000000000P
+ AD=275000000000P PS=3830000U PD=2550000U
* device instance $2 r0 *1 0.92,1.985 pfet_01v8_hvt
M$2 6 2 5 1 pfet_01v8_hvt L=150000U W=2000000U AS=280000000000P
+ AD=275000000000P PS=2560000U PD=2550000U
* device instance $5 r0 *1 2.19,1.985 pfet_01v8_hvt
M$5 7 3 6 1 pfet_01v8_hvt L=150000U W=2000000U AS=270000000000P
+ AD=495000000000P PS=2540000U PD=3990000U
* device instance $7 r0 *1 0.495,0.56 nfet_01v8
M$7 10 4 8 9 nfet_01v8 L=150000U W=650000U AS=185250000000P AD=89375000000P
+ PS=1870000U PD=925000U
* device instance $8 r0 *1 0.92,0.56 nfet_01v8
M$8 7 2 10 9 nfet_01v8 L=150000U W=650000U AS=89375000000P AD=91000000000P
+ PS=925000U PD=930000U
* device instance $9 r0 *1 1.35,0.56 nfet_01v8
M$9 11 2 7 9 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=68250000000P
+ PS=930000U PD=860000U
* device instance $10 r0 *1 1.71,0.56 nfet_01v8
M$10 8 4 11 9 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=107250000000P
+ PS=860000U PD=980000U
* device instance $11 r0 *1 2.19,0.56 nfet_01v8
M$11 7 3 8 9 nfet_01v8 L=150000U W=1300000U AS=195000000000P AD=347750000000P
+ PS=1900000U PD=3020000U
.ENDS sky130_fd_sc_hd__a21oi_2

* cell sky130_fd_sc_hd__xnor2_1
* pin VPB
* pin B
* pin A
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__xnor2_1 1 2 3 4 5 7 9
* net 1 VPB
* net 2 B
* net 3 A
* net 4 Y
* net 5 VPWR
* net 7 VGND
* device instance $1 r0 *1 0.51,1.985 pfet_01v8_hvt
M$1 8 2 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=300000000000P
+ AD=135000000000P PS=2600000U PD=1270000U
* device instance $2 r0 *1 0.93,1.985 pfet_01v8_hvt
M$2 5 3 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=365000000000P PS=1270000U PD=1730000U
* device instance $3 r0 *1 1.81,1.985 pfet_01v8_hvt
M$3 10 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=365000000000P
+ AD=105000000000P PS=1730000U PD=1210000U
* device instance $4 r0 *1 2.17,1.985 pfet_01v8_hvt
M$4 4 2 10 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=165000000000P PS=1210000U PD=1330000U
* device instance $5 r0 *1 2.65,1.985 pfet_01v8_hvt
M$5 5 8 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=165000000000P
+ AD=360000000000P PS=1330000U PD=2720000U
* device instance $6 r0 *1 2.29,0.56 nfet_01v8
M$6 6 2 7 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $7 r0 *1 2.71,0.56 nfet_01v8
M$7 4 8 6 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=195000000000P
+ PS=920000U PD=1900000U
* device instance $8 r0 *1 0.57,0.56 nfet_01v8
M$8 11 2 8 9 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=68250000000P
+ PS=1820000U PD=860000U
* device instance $9 r0 *1 0.93,0.56 nfet_01v8
M$9 7 3 11 9 nfet_01v8 L=150000U W=650000U AS=68250000000P AD=87750000000P
+ PS=860000U PD=920000U
* device instance $10 r0 *1 1.35,0.56 nfet_01v8
M$10 6 3 7 9 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__xnor2_1

* cell sky130_fd_sc_hd__a21o_1
* pin VPB
* pin A1
* pin A2
* pin B1
* pin VGND
* pin VPWR
* pin X
* pin 
.SUBCKT sky130_fd_sc_hd__a21o_1 1 2 3 4 5 7 9 10
* net 1 VPB
* net 2 A1
* net 3 A2
* net 4 B1
* net 5 VGND
* net 7 VPWR
* net 9 X
* device instance $1 r0 *1 1.42,1.985 pfet_01v8_hvt
M$1 6 4 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=137500000000P PS=2520000U PD=1275000U
* device instance $2 r0 *1 1.845,1.985 pfet_01v8_hvt
M$2 7 2 6 1 pfet_01v8_hvt L=150000U W=1000000U AS=137500000000P
+ AD=140000000000P PS=1275000U PD=1280000U
* device instance $3 r0 *1 2.275,1.985 pfet_01v8_hvt
M$3 6 3 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=140000000000P
+ AD=265000000000P PS=1280000U PD=2530000U
* device instance $4 r0 *1 0.48,1.985 pfet_01v8_hvt
M$4 7 8 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=260000000000P PS=2520000U PD=2520000U
* device instance $5 r0 *1 0.48,0.56 nfet_01v8
M$5 5 8 9 10 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=256750000000P
+ PS=1820000U PD=1440000U
* device instance $6 r0 *1 1.42,0.56 nfet_01v8
M$6 8 4 5 10 nfet_01v8 L=150000U W=650000U AS=256750000000P AD=89375000000P
+ PS=1440000U PD=925000U
* device instance $7 r0 *1 1.845,0.56 nfet_01v8
M$7 11 2 8 10 nfet_01v8 L=150000U W=650000U AS=89375000000P AD=91000000000P
+ PS=925000U PD=930000U
* device instance $8 r0 *1 2.275,0.56 nfet_01v8
M$8 5 3 11 10 nfet_01v8 L=150000U W=650000U AS=91000000000P AD=172250000000P
+ PS=930000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21o_1

* cell sky130_fd_sc_hd__nor2b_1
* pin VPB
* pin A
* pin B_N
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor2b_1 1 2 3 4 6 7 8
* net 1 VPB
* net 2 A
* net 3 B_N
* net 4 Y
* net 6 VGND
* net 7 VPWR
* device instance $1 r0 *1 0.71,1.695 pfet_01v8_hvt
M$1 7 3 5 1 pfet_01v8_hvt L=150000U W=420000U AS=109200000000P AD=157300000000P
+ PS=1360000U PD=1390000U
* device instance $2 r0 *1 1.25,1.985 pfet_01v8_hvt
M$2 9 2 7 1 pfet_01v8_hvt L=150000U W=1000000U AS=157300000000P
+ AD=105000000000P PS=1390000U PD=1210000U
* device instance $3 r0 *1 1.61,1.985 pfet_01v8_hvt
M$3 4 5 9 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $4 r0 *1 0.705,0.445 nfet_01v8
M$4 6 3 5 8 nfet_01v8 L=150000U W=420000U AS=109200000000P AD=100250000000P
+ PS=1360000U PD=985000U
* device instance $5 r0 *1 1.19,0.56 nfet_01v8
M$5 4 2 6 8 nfet_01v8 L=150000U W=650000U AS=100250000000P AD=87750000000P
+ PS=985000U PD=920000U
* device instance $6 r0 *1 1.61,0.56 nfet_01v8
M$6 6 5 4 8 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2b_1

* cell sky130_fd_sc_hd__nand2_1
* pin VPB
* pin A
* pin B
* pin Y
* pin VPWR
* pin VGND
* pin 
.SUBCKT sky130_fd_sc_hd__nand2_1 1 2 3 4 5 6 7
* net 1 VPB
* net 2 A
* net 3 B
* net 4 Y
* net 5 VPWR
* net 6 VGND
* device instance $1 r0 *1 0.49,1.985 pfet_01v8_hvt
M$1 4 3 5 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=135000000000P PS=2520000U PD=1270000U
* device instance $2 r0 *1 0.91,1.985 pfet_01v8_hvt
M$2 5 2 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=135000000000P
+ AD=260000000000P PS=1270000U PD=2520000U
* device instance $3 r0 *1 0.49,0.56 nfet_01v8
M$3 8 3 6 7 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $4 r0 *1 0.91,0.56 nfet_01v8
M$4 4 2 8 7 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2_1

* cell sky130_fd_sc_hd__nor2_1
* pin VPB
* pin A
* pin B
* pin Y
* pin VGND
* pin VPWR
* pin 
.SUBCKT sky130_fd_sc_hd__nor2_1 1 2 3 4 5 6 7
* net 1 VPB
* net 2 A
* net 3 B
* net 4 Y
* net 5 VGND
* net 6 VPWR
* device instance $1 r0 *1 0.47,1.985 pfet_01v8_hvt
M$1 8 3 4 1 pfet_01v8_hvt L=150000U W=1000000U AS=260000000000P
+ AD=105000000000P PS=2520000U PD=1210000U
* device instance $2 r0 *1 0.83,1.985 pfet_01v8_hvt
M$2 6 2 8 1 pfet_01v8_hvt L=150000U W=1000000U AS=105000000000P
+ AD=260000000000P PS=1210000U PD=2520000U
* device instance $3 r0 *1 0.47,0.56 nfet_01v8
M$3 4 3 5 7 nfet_01v8 L=150000U W=650000U AS=169000000000P AD=87750000000P
+ PS=1820000U PD=920000U
* device instance $4 r0 *1 0.89,0.56 nfet_01v8
M$4 5 2 4 7 nfet_01v8 L=150000U W=650000U AS=87750000000P AD=169000000000P
+ PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2_1
