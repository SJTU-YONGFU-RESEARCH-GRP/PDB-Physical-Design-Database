module basic_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire spi_clk_en;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 BUF_X4 _203_ (.A(\bit_count[2] ),
    .Z(_038_));
 INV_X1 _204_ (.A(\bit_count[3] ),
    .ZN(_039_));
 BUF_X4 _205_ (.A(_183_),
    .Z(_040_));
 NAND3_X2 _206_ (.A1(_038_),
    .A2(_039_),
    .A3(_040_),
    .ZN(_189_));
 INV_X1 _207_ (.A(_189_),
    .ZN(_194_));
 BUF_X2 _208_ (.A(rst_n),
    .Z(_041_));
 INV_X1 _209_ (.A(_041_),
    .ZN(_042_));
 CLKBUF_X3 _210_ (.A(_042_),
    .Z(_043_));
 CLKBUF_X2 _211_ (.A(\state[0] ),
    .Z(_044_));
 NAND2_X1 _212_ (.A1(net10),
    .A2(_044_),
    .ZN(_045_));
 CLKBUF_X3 _213_ (.A(\state[2] ),
    .Z(_046_));
 CLKBUF_X3 _214_ (.A(_046_),
    .Z(_047_));
 BUF_X4 _215_ (.A(net20),
    .Z(_048_));
 INV_X1 _216_ (.A(_048_),
    .ZN(_049_));
 NAND2_X1 _217_ (.A1(spi_clk_en),
    .A2(_049_),
    .ZN(_050_));
 OAI21_X1 _218_ (.A(_047_),
    .B1(_189_),
    .B2(_050_),
    .ZN(_051_));
 AOI21_X1 _219_ (.A(_043_),
    .B1(_045_),
    .B2(_051_),
    .ZN(_002_));
 CLKBUF_X3 _220_ (.A(\state[1] ),
    .Z(_052_));
 INV_X1 _221_ (.A(_044_),
    .ZN(_053_));
 OAI21_X1 _222_ (.A(_041_),
    .B1(_053_),
    .B2(net10),
    .ZN(_054_));
 OR2_X1 _223_ (.A1(_052_),
    .A2(_054_),
    .ZN(_001_));
 BUF_X2 _224_ (.A(_041_),
    .Z(_055_));
 NAND2_X2 _225_ (.A1(spi_clk_en),
    .A2(_046_),
    .ZN(_056_));
 NOR2_X2 _226_ (.A1(_048_),
    .A2(_056_),
    .ZN(_057_));
 AND3_X1 _227_ (.A1(_055_),
    .A2(_194_),
    .A3(_057_),
    .ZN(_000_));
 NAND3_X1 _228_ (.A1(_038_),
    .A2(\bit_count[0] ),
    .A3(\bit_count[1] ),
    .ZN(_186_));
 OR2_X1 _229_ (.A1(\bit_count[3] ),
    .A2(_186_),
    .ZN(_197_));
 NAND3_X1 _230_ (.A1(_038_),
    .A2(_039_),
    .A3(_040_),
    .ZN(_200_));
 OAI221_X1 _231_ (.A(\bit_count[0] ),
    .B1(_056_),
    .B2(_048_),
    .C1(_047_),
    .C2(_053_),
    .ZN(_058_));
 INV_X1 _232_ (.A(\bit_count[0] ),
    .ZN(_059_));
 NAND2_X1 _233_ (.A1(_059_),
    .A2(_057_),
    .ZN(_060_));
 AOI21_X1 _234_ (.A(_043_),
    .B1(_058_),
    .B2(_060_),
    .ZN(_005_));
 NAND2_X1 _235_ (.A1(_184_),
    .A2(_057_),
    .ZN(_061_));
 OAI221_X1 _236_ (.A(\bit_count[1] ),
    .B1(_056_),
    .B2(_048_),
    .C1(_047_),
    .C2(_053_),
    .ZN(_062_));
 AOI21_X1 _237_ (.A(_043_),
    .B1(_061_),
    .B2(_062_),
    .ZN(_006_));
 INV_X2 _238_ (.A(_046_),
    .ZN(_063_));
 NAND2_X1 _239_ (.A1(_044_),
    .A2(_063_),
    .ZN(_064_));
 NAND2_X1 _240_ (.A1(_038_),
    .A2(_064_),
    .ZN(_065_));
 NAND2_X1 _241_ (.A1(_040_),
    .A2(_057_),
    .ZN(_066_));
 MUX2_X1 _242_ (.A(_038_),
    .B(_065_),
    .S(_066_),
    .Z(_067_));
 NOR2_X1 _243_ (.A1(_043_),
    .A2(_067_),
    .ZN(_007_));
 NAND2_X1 _244_ (.A1(_188_),
    .A2(_057_),
    .ZN(_068_));
 OAI221_X1 _245_ (.A(\bit_count[3] ),
    .B1(_048_),
    .B2(_056_),
    .C1(_047_),
    .C2(_053_),
    .ZN(_069_));
 AOI21_X1 _246_ (.A(_043_),
    .B1(_068_),
    .B2(_069_),
    .ZN(_008_));
 BUF_X2 _247_ (.A(_055_),
    .Z(_070_));
 MUX2_X1 _248_ (.A(net11),
    .B(\rx_shift_reg[0] ),
    .S(_052_),
    .Z(_071_));
 AND2_X1 _249_ (.A1(_070_),
    .A2(_071_),
    .ZN(_009_));
 MUX2_X1 _250_ (.A(net12),
    .B(\rx_shift_reg[1] ),
    .S(_052_),
    .Z(_072_));
 AND2_X1 _251_ (.A1(_070_),
    .A2(_072_),
    .ZN(_010_));
 MUX2_X1 _252_ (.A(net13),
    .B(\rx_shift_reg[2] ),
    .S(_052_),
    .Z(_073_));
 AND2_X1 _253_ (.A1(_070_),
    .A2(_073_),
    .ZN(_011_));
 MUX2_X1 _254_ (.A(net14),
    .B(\rx_shift_reg[3] ),
    .S(_052_),
    .Z(_074_));
 AND2_X1 _255_ (.A1(_070_),
    .A2(_074_),
    .ZN(_012_));
 MUX2_X1 _256_ (.A(net15),
    .B(\rx_shift_reg[4] ),
    .S(_052_),
    .Z(_075_));
 AND2_X1 _257_ (.A1(_070_),
    .A2(_075_),
    .ZN(_013_));
 MUX2_X1 _258_ (.A(net16),
    .B(\rx_shift_reg[5] ),
    .S(_052_),
    .Z(_076_));
 AND2_X1 _259_ (.A1(_070_),
    .A2(_076_),
    .ZN(_014_));
 MUX2_X1 _260_ (.A(net17),
    .B(\rx_shift_reg[6] ),
    .S(_052_),
    .Z(_077_));
 AND2_X1 _261_ (.A1(_070_),
    .A2(_077_),
    .ZN(_015_));
 MUX2_X1 _262_ (.A(net18),
    .B(\rx_shift_reg[7] ),
    .S(_052_),
    .Z(_078_));
 AND2_X1 _263_ (.A1(_070_),
    .A2(_078_),
    .ZN(_016_));
 AND2_X1 _264_ (.A1(_055_),
    .A2(\rx_shift_reg[0] ),
    .ZN(_079_));
 AND2_X1 _265_ (.A1(_041_),
    .A2(net1),
    .ZN(_080_));
 INV_X1 _266_ (.A(_202_),
    .ZN(_081_));
 NOR2_X1 _267_ (.A1(_191_),
    .A2(_199_),
    .ZN(_082_));
 AND2_X1 _268_ (.A1(_198_),
    .A2(_201_),
    .ZN(_083_));
 AND4_X1 _269_ (.A1(_081_),
    .A2(_187_),
    .A3(_082_),
    .A4(_083_),
    .ZN(_084_));
 NOR4_X1 _270_ (.A1(_081_),
    .A2(_187_),
    .A3(_198_),
    .A4(_201_),
    .ZN(_085_));
 AND2_X1 _271_ (.A1(_191_),
    .A2(_199_),
    .ZN(_086_));
 AOI21_X1 _272_ (.A(_084_),
    .B1(_085_),
    .B2(_086_),
    .ZN(_087_));
 INV_X1 _273_ (.A(_003_),
    .ZN(_088_));
 NAND3_X1 _274_ (.A1(_191_),
    .A2(_088_),
    .A3(_188_),
    .ZN(_089_));
 XNOR2_X2 _275_ (.A(_038_),
    .B(_040_),
    .ZN(_090_));
 NOR2_X2 _276_ (.A1(_195_),
    .A2(_192_),
    .ZN(_091_));
 NAND2_X1 _277_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 INV_X1 _278_ (.A(spi_clk_en),
    .ZN(_093_));
 OR3_X2 _279_ (.A1(_093_),
    .A2(_048_),
    .A3(_004_),
    .ZN(_094_));
 OR4_X1 _280_ (.A1(_184_),
    .A2(_089_),
    .A3(_092_),
    .A4(_094_),
    .ZN(_095_));
 NOR2_X1 _281_ (.A1(_087_),
    .A2(_095_),
    .ZN(_096_));
 MUX2_X1 _282_ (.A(_079_),
    .B(_080_),
    .S(_096_),
    .Z(_017_));
 XOR2_X2 _283_ (.A(_038_),
    .B(_040_),
    .Z(_097_));
 NAND3_X2 _284_ (.A1(_084_),
    .A2(_097_),
    .A3(_091_),
    .ZN(_098_));
 INV_X1 _285_ (.A(_184_),
    .ZN(_099_));
 OR3_X2 _286_ (.A1(_099_),
    .A2(_188_),
    .A3(_094_),
    .ZN(_100_));
 NAND2_X1 _287_ (.A1(_059_),
    .A2(net1),
    .ZN(_101_));
 OR3_X1 _288_ (.A1(_098_),
    .A2(_100_),
    .A3(_101_),
    .ZN(_102_));
 NAND3_X1 _289_ (.A1(_039_),
    .A2(_059_),
    .A3(_097_),
    .ZN(_103_));
 OAI21_X1 _290_ (.A(\rx_shift_reg[1] ),
    .B1(_100_),
    .B2(_103_),
    .ZN(_104_));
 AOI21_X1 _291_ (.A(_043_),
    .B1(_102_),
    .B2(_104_),
    .ZN(_018_));
 AND2_X1 _292_ (.A1(_055_),
    .A2(\rx_shift_reg[2] ),
    .ZN(_105_));
 NOR3_X1 _293_ (.A1(_003_),
    .A2(_098_),
    .A3(_100_),
    .ZN(_106_));
 MUX2_X1 _294_ (.A(_105_),
    .B(_080_),
    .S(_106_),
    .Z(_019_));
 OR3_X2 _295_ (.A1(_184_),
    .A2(_188_),
    .A3(_094_),
    .ZN(_107_));
 OR3_X1 _296_ (.A1(_098_),
    .A2(_101_),
    .A3(_107_),
    .ZN(_108_));
 OAI21_X1 _297_ (.A(\rx_shift_reg[3] ),
    .B1(_103_),
    .B2(_107_),
    .ZN(_109_));
 AOI21_X1 _298_ (.A(_043_),
    .B1(_108_),
    .B2(_109_),
    .ZN(_020_));
 AND2_X1 _299_ (.A1(_041_),
    .A2(\rx_shift_reg[4] ),
    .ZN(_110_));
 NOR3_X1 _300_ (.A1(_003_),
    .A2(_098_),
    .A3(_107_),
    .ZN(_111_));
 MUX2_X1 _301_ (.A(_110_),
    .B(_080_),
    .S(_111_),
    .Z(_021_));
 NAND3_X1 _302_ (.A1(_084_),
    .A2(_090_),
    .A3(_091_),
    .ZN(_112_));
 OR3_X1 _303_ (.A1(_100_),
    .A2(_101_),
    .A3(_112_),
    .ZN(_113_));
 NAND3_X1 _304_ (.A1(_039_),
    .A2(_059_),
    .A3(_090_),
    .ZN(_114_));
 OAI21_X1 _305_ (.A(\rx_shift_reg[5] ),
    .B1(_100_),
    .B2(_114_),
    .ZN(_115_));
 AOI21_X1 _306_ (.A(_043_),
    .B1(_113_),
    .B2(_115_),
    .ZN(_022_));
 AND2_X1 _307_ (.A1(_041_),
    .A2(\rx_shift_reg[6] ),
    .ZN(_116_));
 NOR3_X1 _308_ (.A1(_003_),
    .A2(_100_),
    .A3(_112_),
    .ZN(_117_));
 MUX2_X1 _309_ (.A(_116_),
    .B(_080_),
    .S(_117_),
    .Z(_023_));
 OR3_X1 _310_ (.A1(_101_),
    .A2(_107_),
    .A3(_112_),
    .ZN(_118_));
 OAI21_X1 _311_ (.A(\rx_shift_reg[7] ),
    .B1(_107_),
    .B2(_114_),
    .ZN(_119_));
 AOI21_X1 _312_ (.A(_042_),
    .B1(_118_),
    .B2(_119_),
    .ZN(_024_));
 AND2_X1 _313_ (.A1(_052_),
    .A2(_055_),
    .ZN(_025_));
 MUX2_X1 _314_ (.A(_053_),
    .B(_093_),
    .S(_047_),
    .Z(_120_));
 AOI21_X1 _315_ (.A(_057_),
    .B1(_120_),
    .B2(_048_),
    .ZN(_121_));
 NOR2_X1 _316_ (.A1(_043_),
    .A2(_121_),
    .ZN(_026_));
 NAND2_X1 _317_ (.A1(net10),
    .A2(_063_),
    .ZN(_122_));
 OAI21_X1 _318_ (.A(_047_),
    .B1(_048_),
    .B2(_093_),
    .ZN(_123_));
 OAI221_X1 _319_ (.A(_123_),
    .B1(_094_),
    .B2(_194_),
    .C1(_044_),
    .C2(_047_),
    .ZN(_124_));
 MUX2_X1 _320_ (.A(_122_),
    .B(_093_),
    .S(_124_),
    .Z(_125_));
 NOR2_X1 _321_ (.A1(_043_),
    .A2(_125_),
    .ZN(_027_));
 AND2_X1 _322_ (.A1(_053_),
    .A2(net21),
    .ZN(_126_));
 OR2_X1 _323_ (.A1(_001_),
    .A2(_126_),
    .ZN(_028_));
 MUX2_X1 _324_ (.A(net9),
    .B(\tx_shift_reg[6] ),
    .S(_047_),
    .Z(_127_));
 MUX2_X1 _325_ (.A(_046_),
    .B(net10),
    .S(_044_),
    .Z(_128_));
 AND2_X1 _326_ (.A1(spi_clk_en),
    .A2(_048_),
    .ZN(_129_));
 OAI21_X4 _327_ (.A(_128_),
    .B1(_129_),
    .B2(_063_),
    .ZN(_130_));
 NOR3_X1 _328_ (.A1(_049_),
    .A2(_190_),
    .A3(_056_),
    .ZN(_131_));
 NOR2_X1 _329_ (.A1(_130_),
    .A2(_131_),
    .ZN(_132_));
 MUX2_X1 _330_ (.A(net22),
    .B(_127_),
    .S(_132_),
    .Z(_133_));
 AND2_X1 _331_ (.A1(_070_),
    .A2(_133_),
    .ZN(_029_));
 INV_X1 _332_ (.A(_054_),
    .ZN(_134_));
 INV_X1 _333_ (.A(net23),
    .ZN(_135_));
 OAI21_X1 _334_ (.A(_134_),
    .B1(_135_),
    .B2(_044_),
    .ZN(_030_));
 NAND2_X1 _335_ (.A1(\tx_shift_reg[0] ),
    .A2(_130_),
    .ZN(_136_));
 NAND3_X1 _336_ (.A1(_063_),
    .A2(net2),
    .A3(_128_),
    .ZN(_137_));
 AOI21_X1 _337_ (.A(_042_),
    .B1(_136_),
    .B2(_137_),
    .ZN(_031_));
 MUX2_X1 _338_ (.A(net3),
    .B(\tx_shift_reg[0] ),
    .S(_047_),
    .Z(_138_));
 MUX2_X1 _339_ (.A(_138_),
    .B(\tx_shift_reg[1] ),
    .S(_130_),
    .Z(_139_));
 AND2_X1 _340_ (.A1(_070_),
    .A2(_139_),
    .ZN(_032_));
 MUX2_X1 _341_ (.A(net4),
    .B(\tx_shift_reg[1] ),
    .S(_047_),
    .Z(_140_));
 MUX2_X1 _342_ (.A(_140_),
    .B(\tx_shift_reg[2] ),
    .S(_130_),
    .Z(_141_));
 AND2_X1 _343_ (.A1(_055_),
    .A2(_141_),
    .ZN(_033_));
 MUX2_X1 _344_ (.A(net5),
    .B(\tx_shift_reg[2] ),
    .S(_046_),
    .Z(_142_));
 MUX2_X1 _345_ (.A(_142_),
    .B(\tx_shift_reg[3] ),
    .S(_130_),
    .Z(_143_));
 AND2_X1 _346_ (.A1(_055_),
    .A2(_143_),
    .ZN(_034_));
 MUX2_X1 _347_ (.A(net6),
    .B(\tx_shift_reg[3] ),
    .S(_046_),
    .Z(_144_));
 MUX2_X1 _348_ (.A(_144_),
    .B(\tx_shift_reg[4] ),
    .S(_130_),
    .Z(_145_));
 AND2_X1 _349_ (.A1(_055_),
    .A2(_145_),
    .ZN(_035_));
 MUX2_X1 _350_ (.A(net7),
    .B(\tx_shift_reg[4] ),
    .S(_046_),
    .Z(_146_));
 MUX2_X1 _351_ (.A(_146_),
    .B(\tx_shift_reg[5] ),
    .S(_130_),
    .Z(_147_));
 AND2_X1 _352_ (.A1(_055_),
    .A2(_147_),
    .ZN(_036_));
 MUX2_X1 _353_ (.A(net8),
    .B(\tx_shift_reg[5] ),
    .S(_046_),
    .Z(_148_));
 MUX2_X1 _354_ (.A(_148_),
    .B(\tx_shift_reg[6] ),
    .S(_130_),
    .Z(_149_));
 AND2_X1 _355_ (.A1(_055_),
    .A2(_149_),
    .ZN(_037_));
 HA_X1 _356_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_183_),
    .S(_184_));
 HA_X1 _357_ (.A(_185_),
    .B(_186_),
    .CO(_187_),
    .S(_188_));
 HA_X1 _358_ (.A(_185_),
    .B(_189_),
    .CO(_190_),
    .S(_191_));
 HA_X1 _359_ (.A(\bit_count[3] ),
    .B(_189_),
    .CO(_192_),
    .S(_193_));
 HA_X1 _360_ (.A(\bit_count[3] ),
    .B(_194_),
    .CO(_195_),
    .S(_196_));
 HA_X1 _361_ (.A(_185_),
    .B(_197_),
    .CO(_198_),
    .S(_199_));
 HA_X1 _362_ (.A(_185_),
    .B(_200_),
    .CO(_201_),
    .S(_202_));
 DFF_X2 \bit_count[0]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[0] ),
    .QN(_003_));
 DFF_X1 \bit_count[1]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\bit_count[1] ),
    .QN(_179_));
 DFF_X1 \bit_count[2]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\bit_count[2] ),
    .QN(_178_));
 DFF_X2 \bit_count[3]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\bit_count[3] ),
    .QN(_185_));
 DFF_X1 \rx_data[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net11),
    .QN(_177_));
 DFF_X1 \rx_data[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net12),
    .QN(_176_));
 DFF_X1 \rx_data[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net13),
    .QN(_175_));
 DFF_X1 \rx_data[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net14),
    .QN(_174_));
 DFF_X1 \rx_data[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net15),
    .QN(_173_));
 DFF_X1 \rx_data[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net16),
    .QN(_172_));
 DFF_X1 \rx_data[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net17),
    .QN(_171_));
 DFF_X1 \rx_data[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net18),
    .QN(_170_));
 DFF_X1 \rx_shift_reg[0]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[0] ),
    .QN(_169_));
 DFF_X1 \rx_shift_reg[1]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[1] ),
    .QN(_168_));
 DFF_X1 \rx_shift_reg[2]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[2] ),
    .QN(_167_));
 DFF_X1 \rx_shift_reg[3]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[3] ),
    .QN(_166_));
 DFF_X1 \rx_shift_reg[4]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[4] ),
    .QN(_165_));
 DFF_X1 \rx_shift_reg[5]$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[5] ),
    .QN(_164_));
 DFF_X1 \rx_shift_reg[6]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[6] ),
    .QN(_163_));
 DFF_X1 \rx_shift_reg[7]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[7] ),
    .QN(_162_));
 DFF_X1 \rx_valid$_SDFF_PN0_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net19),
    .QN(_161_));
 DFF_X1 \spi_clk$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net20),
    .QN(_160_));
 DFF_X1 \spi_clk_en$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_2_0__leaf_clk),
    .Q(spi_clk_en),
    .QN(_159_));
 DFF_X1 \spi_cs_n$_SDFFE_PN1P_  (.D(_028_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net21),
    .QN(_158_));
 DFF_X1 \spi_mosi$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net22),
    .QN(_180_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\state[0] ),
    .QN(_181_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[1] ),
    .QN(_182_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\state[2] ),
    .QN(_004_));
 DFF_X1 \tx_ready$_SDFFE_PN1P_  (.D(_030_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net23),
    .QN(_157_));
 DFF_X1 \tx_shift_reg[0]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[0] ),
    .QN(_156_));
 DFF_X1 \tx_shift_reg[1]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[1] ),
    .QN(_155_));
 DFF_X1 \tx_shift_reg[2]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[2] ),
    .QN(_154_));
 DFF_X1 \tx_shift_reg[3]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\tx_shift_reg[3] ),
    .QN(_153_));
 DFF_X1 \tx_shift_reg[4]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[4] ),
    .QN(_152_));
 DFF_X1 \tx_shift_reg[5]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[5] ),
    .QN(_151_));
 DFF_X1 \tx_shift_reg[6]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_shift_reg[6] ),
    .QN(_150_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_85 ();
 BUF_X1 input1 (.A(spi_miso),
    .Z(net1));
 BUF_X1 input2 (.A(tx_data[0]),
    .Z(net2));
 BUF_X1 input3 (.A(tx_data[1]),
    .Z(net3));
 BUF_X1 input4 (.A(tx_data[2]),
    .Z(net4));
 BUF_X1 input5 (.A(tx_data[3]),
    .Z(net5));
 BUF_X1 input6 (.A(tx_data[4]),
    .Z(net6));
 BUF_X1 input7 (.A(tx_data[5]),
    .Z(net7));
 BUF_X1 input8 (.A(tx_data[6]),
    .Z(net8));
 BUF_X1 input9 (.A(tx_data[7]),
    .Z(net9));
 BUF_X1 input10 (.A(tx_valid),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(rx_data[0]));
 BUF_X1 output12 (.A(net12),
    .Z(rx_data[1]));
 BUF_X1 output13 (.A(net13),
    .Z(rx_data[2]));
 BUF_X1 output14 (.A(net14),
    .Z(rx_data[3]));
 BUF_X1 output15 (.A(net15),
    .Z(rx_data[4]));
 BUF_X1 output16 (.A(net16),
    .Z(rx_data[5]));
 BUF_X1 output17 (.A(net17),
    .Z(rx_data[6]));
 BUF_X1 output18 (.A(net18),
    .Z(rx_data[7]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_valid));
 BUF_X1 output20 (.A(net20),
    .Z(spi_clk));
 BUF_X1 output21 (.A(net21),
    .Z(spi_cs_n));
 BUF_X1 output22 (.A(net22),
    .Z(spi_mosi));
 BUF_X1 output23 (.A(net23),
    .Z(tx_ready));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X1 clkload0 (.A(clknet_2_1__leaf_clk));
 INV_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_129 ();
 FILLCELL_X1 FILLER_0_133 ();
 FILLCELL_X4 FILLER_0_137 ();
 FILLCELL_X1 FILLER_0_141 ();
 FILLCELL_X8 FILLER_0_145 ();
 FILLCELL_X1 FILLER_0_153 ();
 FILLCELL_X2 FILLER_0_160 ();
 FILLCELL_X2 FILLER_0_168 ();
 FILLCELL_X1 FILLER_0_170 ();
 FILLCELL_X8 FILLER_0_174 ();
 FILLCELL_X4 FILLER_0_182 ();
 FILLCELL_X2 FILLER_0_186 ();
 FILLCELL_X1 FILLER_0_188 ();
 FILLCELL_X16 FILLER_0_192 ();
 FILLCELL_X2 FILLER_0_208 ();
 FILLCELL_X32 FILLER_0_219 ();
 FILLCELL_X32 FILLER_0_251 ();
 FILLCELL_X32 FILLER_0_283 ();
 FILLCELL_X4 FILLER_0_315 ();
 FILLCELL_X2 FILLER_0_319 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X4 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_165 ();
 FILLCELL_X4 FILLER_1_174 ();
 FILLCELL_X2 FILLER_1_178 ();
 FILLCELL_X4 FILLER_1_187 ();
 FILLCELL_X8 FILLER_1_198 ();
 FILLCELL_X4 FILLER_1_206 ();
 FILLCELL_X1 FILLER_1_210 ();
 FILLCELL_X4 FILLER_1_218 ();
 FILLCELL_X2 FILLER_1_222 ();
 FILLCELL_X32 FILLER_1_231 ();
 FILLCELL_X32 FILLER_1_263 ();
 FILLCELL_X16 FILLER_1_295 ();
 FILLCELL_X8 FILLER_1_311 ();
 FILLCELL_X2 FILLER_1_319 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X8 FILLER_2_161 ();
 FILLCELL_X1 FILLER_2_169 ();
 FILLCELL_X2 FILLER_2_181 ();
 FILLCELL_X8 FILLER_2_187 ();
 FILLCELL_X2 FILLER_2_195 ();
 FILLCELL_X1 FILLER_2_197 ();
 FILLCELL_X16 FILLER_2_205 ();
 FILLCELL_X1 FILLER_2_221 ();
 FILLCELL_X32 FILLER_2_233 ();
 FILLCELL_X32 FILLER_2_265 ();
 FILLCELL_X16 FILLER_2_297 ();
 FILLCELL_X8 FILLER_2_313 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X16 FILLER_3_129 ();
 FILLCELL_X8 FILLER_3_145 ();
 FILLCELL_X2 FILLER_3_153 ();
 FILLCELL_X1 FILLER_3_155 ();
 FILLCELL_X4 FILLER_3_173 ();
 FILLCELL_X2 FILLER_3_177 ();
 FILLCELL_X1 FILLER_3_179 ();
 FILLCELL_X8 FILLER_3_218 ();
 FILLCELL_X4 FILLER_3_226 ();
 FILLCELL_X32 FILLER_3_247 ();
 FILLCELL_X32 FILLER_3_279 ();
 FILLCELL_X8 FILLER_3_311 ();
 FILLCELL_X2 FILLER_3_319 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X4 FILLER_4_161 ();
 FILLCELL_X2 FILLER_4_165 ();
 FILLCELL_X32 FILLER_4_174 ();
 FILLCELL_X8 FILLER_4_206 ();
 FILLCELL_X4 FILLER_4_221 ();
 FILLCELL_X2 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_234 ();
 FILLCELL_X32 FILLER_4_266 ();
 FILLCELL_X16 FILLER_4_298 ();
 FILLCELL_X4 FILLER_4_314 ();
 FILLCELL_X2 FILLER_4_318 ();
 FILLCELL_X1 FILLER_4_320 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X16 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_145 ();
 FILLCELL_X32 FILLER_5_177 ();
 FILLCELL_X32 FILLER_5_235 ();
 FILLCELL_X32 FILLER_5_267 ();
 FILLCELL_X16 FILLER_5_299 ();
 FILLCELL_X4 FILLER_5_315 ();
 FILLCELL_X2 FILLER_5_319 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X4 FILLER_6_161 ();
 FILLCELL_X2 FILLER_6_165 ();
 FILLCELL_X1 FILLER_6_167 ();
 FILLCELL_X32 FILLER_6_175 ();
 FILLCELL_X32 FILLER_6_207 ();
 FILLCELL_X32 FILLER_6_239 ();
 FILLCELL_X32 FILLER_6_271 ();
 FILLCELL_X16 FILLER_6_303 ();
 FILLCELL_X2 FILLER_6_319 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X8 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_176 ();
 FILLCELL_X32 FILLER_7_208 ();
 FILLCELL_X32 FILLER_7_240 ();
 FILLCELL_X32 FILLER_7_272 ();
 FILLCELL_X16 FILLER_7_304 ();
 FILLCELL_X1 FILLER_7_320 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X16 FILLER_8_129 ();
 FILLCELL_X8 FILLER_8_145 ();
 FILLCELL_X4 FILLER_8_153 ();
 FILLCELL_X1 FILLER_8_157 ();
 FILLCELL_X16 FILLER_8_179 ();
 FILLCELL_X1 FILLER_8_195 ();
 FILLCELL_X16 FILLER_8_213 ();
 FILLCELL_X2 FILLER_8_236 ();
 FILLCELL_X8 FILLER_8_242 ();
 FILLCELL_X4 FILLER_8_250 ();
 FILLCELL_X2 FILLER_8_254 ();
 FILLCELL_X32 FILLER_8_260 ();
 FILLCELL_X16 FILLER_8_292 ();
 FILLCELL_X8 FILLER_8_308 ();
 FILLCELL_X4 FILLER_8_316 ();
 FILLCELL_X1 FILLER_8_320 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X1 FILLER_9_129 ();
 FILLCELL_X1 FILLER_9_149 ();
 FILLCELL_X8 FILLER_9_154 ();
 FILLCELL_X1 FILLER_9_162 ();
 FILLCELL_X8 FILLER_9_191 ();
 FILLCELL_X2 FILLER_9_199 ();
 FILLCELL_X16 FILLER_9_226 ();
 FILLCELL_X32 FILLER_9_259 ();
 FILLCELL_X16 FILLER_9_291 ();
 FILLCELL_X8 FILLER_9_307 ();
 FILLCELL_X4 FILLER_9_315 ();
 FILLCELL_X2 FILLER_9_319 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X8 FILLER_10_161 ();
 FILLCELL_X4 FILLER_10_169 ();
 FILLCELL_X8 FILLER_10_176 ();
 FILLCELL_X4 FILLER_10_184 ();
 FILLCELL_X1 FILLER_10_188 ();
 FILLCELL_X4 FILLER_10_196 ();
 FILLCELL_X1 FILLER_10_203 ();
 FILLCELL_X2 FILLER_10_215 ();
 FILLCELL_X1 FILLER_10_217 ();
 FILLCELL_X32 FILLER_10_222 ();
 FILLCELL_X32 FILLER_10_254 ();
 FILLCELL_X32 FILLER_10_286 ();
 FILLCELL_X2 FILLER_10_318 ();
 FILLCELL_X1 FILLER_10_320 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X8 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_137 ();
 FILLCELL_X2 FILLER_11_141 ();
 FILLCELL_X8 FILLER_11_147 ();
 FILLCELL_X2 FILLER_11_155 ();
 FILLCELL_X1 FILLER_11_157 ();
 FILLCELL_X8 FILLER_11_160 ();
 FILLCELL_X4 FILLER_11_168 ();
 FILLCELL_X4 FILLER_11_176 ();
 FILLCELL_X2 FILLER_11_180 ();
 FILLCELL_X1 FILLER_11_182 ();
 FILLCELL_X1 FILLER_11_195 ();
 FILLCELL_X1 FILLER_11_207 ();
 FILLCELL_X32 FILLER_11_212 ();
 FILLCELL_X32 FILLER_11_244 ();
 FILLCELL_X32 FILLER_11_276 ();
 FILLCELL_X8 FILLER_11_308 ();
 FILLCELL_X4 FILLER_11_316 ();
 FILLCELL_X1 FILLER_11_320 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_113 ();
 FILLCELL_X4 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_125 ();
 FILLCELL_X1 FILLER_12_127 ();
 FILLCELL_X2 FILLER_12_149 ();
 FILLCELL_X8 FILLER_12_155 ();
 FILLCELL_X4 FILLER_12_163 ();
 FILLCELL_X4 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_180 ();
 FILLCELL_X1 FILLER_12_182 ();
 FILLCELL_X1 FILLER_12_193 ();
 FILLCELL_X4 FILLER_12_200 ();
 FILLCELL_X2 FILLER_12_204 ();
 FILLCELL_X16 FILLER_12_211 ();
 FILLCELL_X1 FILLER_12_227 ();
 FILLCELL_X32 FILLER_12_235 ();
 FILLCELL_X32 FILLER_12_267 ();
 FILLCELL_X16 FILLER_12_299 ();
 FILLCELL_X4 FILLER_12_315 ();
 FILLCELL_X2 FILLER_12_319 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X4 FILLER_13_129 ();
 FILLCELL_X2 FILLER_13_133 ();
 FILLCELL_X16 FILLER_13_152 ();
 FILLCELL_X8 FILLER_13_168 ();
 FILLCELL_X4 FILLER_13_176 ();
 FILLCELL_X1 FILLER_13_180 ();
 FILLCELL_X16 FILLER_13_190 ();
 FILLCELL_X4 FILLER_13_206 ();
 FILLCELL_X1 FILLER_13_210 ();
 FILLCELL_X16 FILLER_13_218 ();
 FILLCELL_X8 FILLER_13_234 ();
 FILLCELL_X2 FILLER_13_242 ();
 FILLCELL_X1 FILLER_13_244 ();
 FILLCELL_X8 FILLER_13_267 ();
 FILLCELL_X2 FILLER_13_275 ();
 FILLCELL_X1 FILLER_13_277 ();
 FILLCELL_X32 FILLER_13_282 ();
 FILLCELL_X4 FILLER_13_314 ();
 FILLCELL_X2 FILLER_13_318 ();
 FILLCELL_X1 FILLER_13_320 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X16 FILLER_14_193 ();
 FILLCELL_X4 FILLER_14_209 ();
 FILLCELL_X1 FILLER_14_213 ();
 FILLCELL_X32 FILLER_14_224 ();
 FILLCELL_X32 FILLER_14_256 ();
 FILLCELL_X32 FILLER_14_288 ();
 FILLCELL_X1 FILLER_14_320 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X16 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_145 ();
 FILLCELL_X1 FILLER_15_153 ();
 FILLCELL_X8 FILLER_15_171 ();
 FILLCELL_X1 FILLER_15_179 ();
 FILLCELL_X16 FILLER_15_183 ();
 FILLCELL_X2 FILLER_15_199 ();
 FILLCELL_X8 FILLER_15_207 ();
 FILLCELL_X4 FILLER_15_215 ();
 FILLCELL_X2 FILLER_15_219 ();
 FILLCELL_X32 FILLER_15_236 ();
 FILLCELL_X16 FILLER_15_268 ();
 FILLCELL_X4 FILLER_15_284 ();
 FILLCELL_X2 FILLER_15_288 ();
 FILLCELL_X4 FILLER_15_294 ();
 FILLCELL_X2 FILLER_15_315 ();
 FILLCELL_X1 FILLER_15_320 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X1 FILLER_16_161 ();
 FILLCELL_X8 FILLER_16_169 ();
 FILLCELL_X4 FILLER_16_177 ();
 FILLCELL_X8 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_201 ();
 FILLCELL_X1 FILLER_16_203 ();
 FILLCELL_X4 FILLER_16_208 ();
 FILLCELL_X32 FILLER_16_231 ();
 FILLCELL_X16 FILLER_16_263 ();
 FILLCELL_X8 FILLER_16_279 ();
 FILLCELL_X4 FILLER_16_287 ();
 FILLCELL_X16 FILLER_16_294 ();
 FILLCELL_X8 FILLER_16_310 ();
 FILLCELL_X2 FILLER_16_318 ();
 FILLCELL_X1 FILLER_16_320 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_161 ();
 FILLCELL_X4 FILLER_17_169 ();
 FILLCELL_X2 FILLER_17_173 ();
 FILLCELL_X1 FILLER_17_175 ();
 FILLCELL_X4 FILLER_17_197 ();
 FILLCELL_X2 FILLER_17_201 ();
 FILLCELL_X1 FILLER_17_203 ();
 FILLCELL_X8 FILLER_17_207 ();
 FILLCELL_X4 FILLER_17_215 ();
 FILLCELL_X2 FILLER_17_219 ();
 FILLCELL_X1 FILLER_17_221 ();
 FILLCELL_X32 FILLER_17_232 ();
 FILLCELL_X32 FILLER_17_264 ();
 FILLCELL_X8 FILLER_17_313 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X2 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_38 ();
 FILLCELL_X32 FILLER_18_70 ();
 FILLCELL_X32 FILLER_18_102 ();
 FILLCELL_X32 FILLER_18_134 ();
 FILLCELL_X8 FILLER_18_166 ();
 FILLCELL_X1 FILLER_18_174 ();
 FILLCELL_X1 FILLER_18_178 ();
 FILLCELL_X2 FILLER_18_183 ();
 FILLCELL_X2 FILLER_18_195 ();
 FILLCELL_X2 FILLER_18_201 ();
 FILLCELL_X4 FILLER_18_212 ();
 FILLCELL_X2 FILLER_18_216 ();
 FILLCELL_X8 FILLER_18_254 ();
 FILLCELL_X2 FILLER_18_262 ();
 FILLCELL_X2 FILLER_18_285 ();
 FILLCELL_X2 FILLER_18_294 ();
 FILLCELL_X1 FILLER_18_296 ();
 FILLCELL_X8 FILLER_18_301 ();
 FILLCELL_X4 FILLER_18_309 ();
 FILLCELL_X1 FILLER_18_316 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X8 FILLER_19_200 ();
 FILLCELL_X8 FILLER_19_212 ();
 FILLCELL_X4 FILLER_19_220 ();
 FILLCELL_X1 FILLER_19_224 ();
 FILLCELL_X2 FILLER_19_248 ();
 FILLCELL_X8 FILLER_19_256 ();
 FILLCELL_X1 FILLER_19_264 ();
 FILLCELL_X32 FILLER_19_272 ();
 FILLCELL_X16 FILLER_19_304 ();
 FILLCELL_X1 FILLER_19_320 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_169 ();
 FILLCELL_X1 FILLER_20_173 ();
 FILLCELL_X1 FILLER_20_177 ();
 FILLCELL_X32 FILLER_20_181 ();
 FILLCELL_X8 FILLER_20_213 ();
 FILLCELL_X4 FILLER_20_221 ();
 FILLCELL_X2 FILLER_20_225 ();
 FILLCELL_X8 FILLER_20_233 ();
 FILLCELL_X2 FILLER_20_241 ();
 FILLCELL_X8 FILLER_20_254 ();
 FILLCELL_X4 FILLER_20_262 ();
 FILLCELL_X16 FILLER_20_270 ();
 FILLCELL_X4 FILLER_20_286 ();
 FILLCELL_X2 FILLER_20_290 ();
 FILLCELL_X8 FILLER_20_303 ();
 FILLCELL_X4 FILLER_20_311 ();
 FILLCELL_X1 FILLER_20_315 ();
 FILLCELL_X2 FILLER_20_319 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_169 ();
 FILLCELL_X1 FILLER_21_171 ();
 FILLCELL_X8 FILLER_21_179 ();
 FILLCELL_X4 FILLER_21_187 ();
 FILLCELL_X16 FILLER_21_210 ();
 FILLCELL_X2 FILLER_21_226 ();
 FILLCELL_X32 FILLER_21_231 ();
 FILLCELL_X1 FILLER_21_263 ();
 FILLCELL_X8 FILLER_21_288 ();
 FILLCELL_X2 FILLER_21_296 ();
 FILLCELL_X1 FILLER_21_298 ();
 FILLCELL_X4 FILLER_21_316 ();
 FILLCELL_X1 FILLER_21_320 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X16 FILLER_22_129 ();
 FILLCELL_X8 FILLER_22_145 ();
 FILLCELL_X16 FILLER_22_180 ();
 FILLCELL_X2 FILLER_22_196 ();
 FILLCELL_X1 FILLER_22_198 ();
 FILLCELL_X32 FILLER_22_201 ();
 FILLCELL_X32 FILLER_22_233 ();
 FILLCELL_X32 FILLER_22_265 ();
 FILLCELL_X16 FILLER_22_297 ();
 FILLCELL_X8 FILLER_22_313 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_197 ();
 FILLCELL_X8 FILLER_23_212 ();
 FILLCELL_X2 FILLER_23_237 ();
 FILLCELL_X1 FILLER_23_239 ();
 FILLCELL_X8 FILLER_23_244 ();
 FILLCELL_X4 FILLER_23_252 ();
 FILLCELL_X2 FILLER_23_256 ();
 FILLCELL_X32 FILLER_23_263 ();
 FILLCELL_X16 FILLER_23_295 ();
 FILLCELL_X8 FILLER_23_311 ();
 FILLCELL_X2 FILLER_23_319 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X16 FILLER_24_193 ();
 FILLCELL_X4 FILLER_24_209 ();
 FILLCELL_X16 FILLER_24_220 ();
 FILLCELL_X16 FILLER_24_244 ();
 FILLCELL_X8 FILLER_24_260 ();
 FILLCELL_X1 FILLER_24_268 ();
 FILLCELL_X2 FILLER_24_276 ();
 FILLCELL_X8 FILLER_24_282 ();
 FILLCELL_X1 FILLER_24_290 ();
 FILLCELL_X8 FILLER_24_302 ();
 FILLCELL_X4 FILLER_24_310 ();
 FILLCELL_X2 FILLER_24_314 ();
 FILLCELL_X1 FILLER_24_316 ();
 FILLCELL_X1 FILLER_24_320 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X16 FILLER_25_161 ();
 FILLCELL_X4 FILLER_25_177 ();
 FILLCELL_X2 FILLER_25_181 ();
 FILLCELL_X8 FILLER_25_185 ();
 FILLCELL_X4 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_200 ();
 FILLCELL_X16 FILLER_25_232 ();
 FILLCELL_X8 FILLER_25_248 ();
 FILLCELL_X1 FILLER_25_256 ();
 FILLCELL_X8 FILLER_25_261 ();
 FILLCELL_X4 FILLER_25_269 ();
 FILLCELL_X2 FILLER_25_273 ();
 FILLCELL_X4 FILLER_25_292 ();
 FILLCELL_X8 FILLER_25_313 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X16 FILLER_26_161 ();
 FILLCELL_X8 FILLER_26_177 ();
 FILLCELL_X2 FILLER_26_185 ();
 FILLCELL_X1 FILLER_26_187 ();
 FILLCELL_X1 FILLER_26_196 ();
 FILLCELL_X16 FILLER_26_207 ();
 FILLCELL_X2 FILLER_26_223 ();
 FILLCELL_X16 FILLER_26_235 ();
 FILLCELL_X8 FILLER_26_251 ();
 FILLCELL_X4 FILLER_26_259 ();
 FILLCELL_X2 FILLER_26_263 ();
 FILLCELL_X1 FILLER_26_265 ();
 FILLCELL_X4 FILLER_26_273 ();
 FILLCELL_X32 FILLER_26_281 ();
 FILLCELL_X8 FILLER_26_313 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X16 FILLER_27_161 ();
 FILLCELL_X2 FILLER_27_177 ();
 FILLCELL_X8 FILLER_27_204 ();
 FILLCELL_X4 FILLER_27_212 ();
 FILLCELL_X2 FILLER_27_216 ();
 FILLCELL_X4 FILLER_27_226 ();
 FILLCELL_X1 FILLER_27_230 ();
 FILLCELL_X16 FILLER_27_239 ();
 FILLCELL_X8 FILLER_27_255 ();
 FILLCELL_X2 FILLER_27_263 ();
 FILLCELL_X1 FILLER_27_265 ();
 FILLCELL_X2 FILLER_27_283 ();
 FILLCELL_X1 FILLER_27_285 ();
 FILLCELL_X16 FILLER_27_297 ();
 FILLCELL_X8 FILLER_27_313 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X16 FILLER_28_161 ();
 FILLCELL_X4 FILLER_28_177 ();
 FILLCELL_X2 FILLER_28_181 ();
 FILLCELL_X8 FILLER_28_200 ();
 FILLCELL_X4 FILLER_28_208 ();
 FILLCELL_X2 FILLER_28_229 ();
 FILLCELL_X1 FILLER_28_231 ();
 FILLCELL_X32 FILLER_28_249 ();
 FILLCELL_X8 FILLER_28_281 ();
 FILLCELL_X2 FILLER_28_289 ();
 FILLCELL_X1 FILLER_28_291 ();
 FILLCELL_X2 FILLER_28_309 ();
 FILLCELL_X4 FILLER_28_314 ();
 FILLCELL_X2 FILLER_28_318 ();
 FILLCELL_X1 FILLER_28_320 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X4 FILLER_29_161 ();
 FILLCELL_X1 FILLER_29_165 ();
 FILLCELL_X32 FILLER_29_173 ();
 FILLCELL_X32 FILLER_29_205 ();
 FILLCELL_X8 FILLER_29_237 ();
 FILLCELL_X4 FILLER_29_245 ();
 FILLCELL_X2 FILLER_29_249 ();
 FILLCELL_X1 FILLER_29_251 ();
 FILLCELL_X32 FILLER_29_263 ();
 FILLCELL_X16 FILLER_29_295 ();
 FILLCELL_X8 FILLER_29_311 ();
 FILLCELL_X2 FILLER_29_319 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X16 FILLER_30_129 ();
 FILLCELL_X4 FILLER_30_145 ();
 FILLCELL_X1 FILLER_30_149 ();
 FILLCELL_X1 FILLER_30_167 ();
 FILLCELL_X32 FILLER_30_172 ();
 FILLCELL_X32 FILLER_30_204 ();
 FILLCELL_X16 FILLER_30_236 ();
 FILLCELL_X8 FILLER_30_252 ();
 FILLCELL_X1 FILLER_30_260 ();
 FILLCELL_X32 FILLER_30_278 ();
 FILLCELL_X8 FILLER_30_310 ();
 FILLCELL_X2 FILLER_30_318 ();
 FILLCELL_X1 FILLER_30_320 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X16 FILLER_31_161 ();
 FILLCELL_X4 FILLER_31_177 ();
 FILLCELL_X2 FILLER_31_181 ();
 FILLCELL_X1 FILLER_31_183 ();
 FILLCELL_X16 FILLER_31_195 ();
 FILLCELL_X4 FILLER_31_211 ();
 FILLCELL_X32 FILLER_31_226 ();
 FILLCELL_X16 FILLER_31_258 ();
 FILLCELL_X8 FILLER_31_274 ();
 FILLCELL_X4 FILLER_31_282 ();
 FILLCELL_X2 FILLER_31_286 ();
 FILLCELL_X16 FILLER_31_291 ();
 FILLCELL_X8 FILLER_31_307 ();
 FILLCELL_X4 FILLER_31_315 ();
 FILLCELL_X2 FILLER_31_319 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X16 FILLER_32_161 ();
 FILLCELL_X1 FILLER_32_177 ();
 FILLCELL_X16 FILLER_32_195 ();
 FILLCELL_X32 FILLER_32_228 ();
 FILLCELL_X32 FILLER_32_260 ();
 FILLCELL_X16 FILLER_32_292 ();
 FILLCELL_X8 FILLER_32_308 ();
 FILLCELL_X4 FILLER_32_316 ();
 FILLCELL_X1 FILLER_32_320 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X16 FILLER_42_129 ();
 FILLCELL_X8 FILLER_42_145 ();
 FILLCELL_X2 FILLER_42_153 ();
 FILLCELL_X16 FILLER_42_158 ();
 FILLCELL_X8 FILLER_42_174 ();
 FILLCELL_X4 FILLER_42_182 ();
 FILLCELL_X2 FILLER_42_186 ();
 FILLCELL_X1 FILLER_42_188 ();
 FILLCELL_X2 FILLER_42_192 ();
 FILLCELL_X1 FILLER_42_194 ();
 FILLCELL_X16 FILLER_42_198 ();
 FILLCELL_X4 FILLER_42_214 ();
 FILLCELL_X1 FILLER_42_218 ();
 FILLCELL_X32 FILLER_42_222 ();
 FILLCELL_X32 FILLER_42_254 ();
 FILLCELL_X32 FILLER_42_286 ();
 FILLCELL_X2 FILLER_42_318 ();
 FILLCELL_X1 FILLER_42_320 ();
endmodule
